// Verilog netlist created by TD v4.5.12562
// Thu Dec 19 17:42:10 2019

`timescale 1ns / 1ps
module CPLD_SOC_AHB_TOP  // CPLD_SOC_AHB_TOP.v(1)
  (
  clkin,
  limit_l,
  limit_r,
  rst_n,
  dir,
  gpio_out,
  ledout,
  pwm
  );

  input clkin;  // CPLD_SOC_AHB_TOP.v(3)
  input [15:0] limit_l;  // CPLD_SOC_AHB_TOP.v(5)
  input [15:0] limit_r;  // CPLD_SOC_AHB_TOP.v(6)
  input rst_n;  // CPLD_SOC_AHB_TOP.v(4)
  output [15:0] dir;  // CPLD_SOC_AHB_TOP.v(7)
  output [31:0] gpio_out;  // CPLD_SOC_AHB_TOP.v(8)
  output [3:0] ledout;  // CPLD_SOC_AHB_TOP.v(10)
  output [15:0] pwm;  // CPLD_SOC_AHB_TOP.v(7)

  wire [26:0] \PWM0/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWM0/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWM0/n12 ;
  wire [24:0] \PWM0/n26 ;
  wire [31:0] \PWM0/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWM1/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWM1/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWM1/n12 ;
  wire [24:0] \PWM1/n26 ;
  wire [31:0] \PWM1/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWM2/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWM2/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWM2/n12 ;
  wire [24:0] \PWM2/n26 ;
  wire [31:0] \PWM2/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWM3/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWM3/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWM3/n12 ;
  wire [24:0] \PWM3/n26 ;
  wire [31:0] \PWM3/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWM4/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWM4/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWM4/n12 ;
  wire [24:0] \PWM4/n26 ;
  wire [31:0] \PWM4/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWM5/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWM5/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWM5/n12 ;
  wire [24:0] \PWM5/n26 ;
  wire [31:0] \PWM5/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWM6/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWM6/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWM6/n12 ;
  wire [24:0] \PWM6/n26 ;
  wire [31:0] \PWM6/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWM7/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWM7/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWM7/n12 ;
  wire [24:0] \PWM7/n26 ;
  wire [31:0] \PWM7/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWM8/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWM8/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWM8/n12 ;
  wire [24:0] \PWM8/n26 ;
  wire [31:0] \PWM8/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWM9/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWM9/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWM9/n12 ;
  wire [24:0] \PWM9/n26 ;
  wire [31:0] \PWM9/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWMA/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWMA/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWMA/n12 ;
  wire [24:0] \PWMA/n26 ;
  wire [31:0] \PWMA/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWMB/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWMB/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWMB/n12 ;
  wire [24:0] \PWMB/n26 ;
  wire [31:0] \PWMB/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWMC/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWMC/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWMC/n12 ;
  wire [24:0] \PWMC/n26 ;
  wire [31:0] \PWMC/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWMD/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWMD/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWMD/n12 ;
  wire [24:0] \PWMD/n26 ;
  wire [31:0] \PWMD/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWME/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWME/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWME/n12 ;
  wire [24:0] \PWME/n26 ;
  wire [31:0] \PWME/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWMF/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWMF/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWMF/n12 ;
  wire [24:0] \PWMF/n26 ;
  wire [31:0] \PWMF/pnumr ;  // src/OnePWM.v(47)
  wire [31:0] \U_AHB/h2h_haddr ;  // src/AHB.v(23)
  wire [31:0] \U_AHB/h2h_haddrw ;  // src/AHB.v(16)
  wire [31:0] \U_AHB/h2h_hrdata ;  // src/AHB.v(18)
  wire [31:0] \U_AHB/h2h_hwdata ;  // src/AHB.v(17)
  wire [15:0] dir_pad;  // CPLD_SOC_AHB_TOP.v(7)
  wire [31:0] freq0;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freq1;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freq2;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freq3;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freq4;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freq5;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freq6;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freq7;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freq8;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freq9;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freqA;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freqB;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freqC;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freqD;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freqE;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freqF;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] gpio_out_pad;  // CPLD_SOC_AHB_TOP.v(8)
  wire [3:0] ledout_pad;  // CPLD_SOC_AHB_TOP.v(10)
  wire [15:0] limit_l_pad;  // CPLD_SOC_AHB_TOP.v(5)
  wire [15:0] limit_r_pad;  // CPLD_SOC_AHB_TOP.v(6)
  wire [31:0] n2;
  wire [32:0] pnum0;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnum1;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnum2;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnum3;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnum4;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnum5;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnum6;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnum7;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnum8;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnum9;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnumA;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnumB;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnumC;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnumD;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnumE;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnumF;  // CPLD_SOC_AHB_TOP.v(54)
  wire [23:0] pnumcnt0;  // CPLD_SOC_AHB_TOP.v(61)
  wire [23:0] pnumcnt1;  // CPLD_SOC_AHB_TOP.v(62)
  wire [23:0] pnumcnt2;  // CPLD_SOC_AHB_TOP.v(63)
  wire [23:0] pnumcnt3;  // CPLD_SOC_AHB_TOP.v(64)
  wire [23:0] pnumcnt4;  // CPLD_SOC_AHB_TOP.v(65)
  wire [23:0] pnumcnt5;  // CPLD_SOC_AHB_TOP.v(66)
  wire [23:0] pnumcnt6;  // CPLD_SOC_AHB_TOP.v(67)
  wire [23:0] pnumcnt7;  // CPLD_SOC_AHB_TOP.v(68)
  wire [23:0] pnumcnt8;  // CPLD_SOC_AHB_TOP.v(69)
  wire [23:0] pnumcnt9;  // CPLD_SOC_AHB_TOP.v(70)
  wire [23:0] pnumcntA;  // CPLD_SOC_AHB_TOP.v(71)
  wire [23:0] pnumcntB;  // CPLD_SOC_AHB_TOP.v(72)
  wire [23:0] pnumcntC;  // CPLD_SOC_AHB_TOP.v(73)
  wire [23:0] pnumcntD;  // CPLD_SOC_AHB_TOP.v(74)
  wire [23:0] pnumcntE;  // CPLD_SOC_AHB_TOP.v(75)
  wire [23:0] pnumcntF;  // CPLD_SOC_AHB_TOP.v(76)
  wire [15:0] pwm_pad;  // CPLD_SOC_AHB_TOP.v(7)
  wire [31:0] pwm_start_stop;  // CPLD_SOC_AHB_TOP.v(52)
  wire [15:0] pwm_state_read;  // CPLD_SOC_AHB_TOP.v(78)
  wire [31:0] timer;  // CPLD_SOC_AHB_TOP.v(26)
  wire \PWM0/RemaTxNum[0]_keep ;
  wire \PWM0/RemaTxNum[10]_keep ;
  wire \PWM0/RemaTxNum[11]_keep ;
  wire \PWM0/RemaTxNum[12]_keep ;
  wire \PWM0/RemaTxNum[13]_keep ;
  wire \PWM0/RemaTxNum[14]_keep ;
  wire \PWM0/RemaTxNum[15]_keep ;
  wire \PWM0/RemaTxNum[16]_keep ;
  wire \PWM0/RemaTxNum[17]_keep ;
  wire \PWM0/RemaTxNum[18]_keep ;
  wire \PWM0/RemaTxNum[19]_keep ;
  wire \PWM0/RemaTxNum[1]_keep ;
  wire \PWM0/RemaTxNum[20]_keep ;
  wire \PWM0/RemaTxNum[21]_keep ;
  wire \PWM0/RemaTxNum[22]_keep ;
  wire \PWM0/RemaTxNum[23]_keep ;
  wire \PWM0/RemaTxNum[2]_keep ;
  wire \PWM0/RemaTxNum[3]_keep ;
  wire \PWM0/RemaTxNum[4]_keep ;
  wire \PWM0/RemaTxNum[5]_keep ;
  wire \PWM0/RemaTxNum[6]_keep ;
  wire \PWM0/RemaTxNum[7]_keep ;
  wire \PWM0/RemaTxNum[8]_keep ;
  wire \PWM0/RemaTxNum[9]_keep ;
  wire \PWM0/dir_keep ;
  wire \PWM0/mux3_b0_sel_is_3_o ;
  wire \PWM0/n0_lutinv ;
  wire \PWM0/n11 ;
  wire \PWM0/n24 ;
  wire \PWM0/n25_neg_lutinv ;
  wire \PWM0/pnumr[0]_keep ;
  wire \PWM0/pnumr[10]_keep ;
  wire \PWM0/pnumr[11]_keep ;
  wire \PWM0/pnumr[12]_keep ;
  wire \PWM0/pnumr[13]_keep ;
  wire \PWM0/pnumr[14]_keep ;
  wire \PWM0/pnumr[15]_keep ;
  wire \PWM0/pnumr[16]_keep ;
  wire \PWM0/pnumr[17]_keep ;
  wire \PWM0/pnumr[18]_keep ;
  wire \PWM0/pnumr[19]_keep ;
  wire \PWM0/pnumr[1]_keep ;
  wire \PWM0/pnumr[20]_keep ;
  wire \PWM0/pnumr[21]_keep ;
  wire \PWM0/pnumr[22]_keep ;
  wire \PWM0/pnumr[23]_keep ;
  wire \PWM0/pnumr[24]_keep ;
  wire \PWM0/pnumr[25]_keep ;
  wire \PWM0/pnumr[26]_keep ;
  wire \PWM0/pnumr[27]_keep ;
  wire \PWM0/pnumr[28]_keep ;
  wire \PWM0/pnumr[29]_keep ;
  wire \PWM0/pnumr[2]_keep ;
  wire \PWM0/pnumr[30]_keep ;
  wire \PWM0/pnumr[31]_keep ;
  wire \PWM0/pnumr[3]_keep ;
  wire \PWM0/pnumr[4]_keep ;
  wire \PWM0/pnumr[5]_keep ;
  wire \PWM0/pnumr[6]_keep ;
  wire \PWM0/pnumr[7]_keep ;
  wire \PWM0/pnumr[8]_keep ;
  wire \PWM0/pnumr[9]_keep ;
  wire \PWM0/pwm_keep ;
  wire \PWM0/stopreq ;  // src/OnePWM.v(14)
  wire \PWM0/stopreq_keep ;
  wire \PWM0/sub0/c11 ;
  wire \PWM0/sub0/c15 ;
  wire \PWM0/sub0/c19 ;
  wire \PWM0/sub0/c23 ;
  wire \PWM0/sub0/c3 ;
  wire \PWM0/sub0/c7 ;
  wire \PWM0/sub1/c1 ;
  wire \PWM0/sub1/c11 ;
  wire \PWM0/sub1/c13 ;
  wire \PWM0/sub1/c15 ;
  wire \PWM0/sub1/c17 ;
  wire \PWM0/sub1/c19 ;
  wire \PWM0/sub1/c21 ;
  wire \PWM0/sub1/c23 ;
  wire \PWM0/sub1/c3 ;
  wire \PWM0/sub1/c5 ;
  wire \PWM0/sub1/c7 ;
  wire \PWM0/sub1/c9 ;
  wire \PWM0/u14_sel_is_1_o ;
  wire \PWM1/RemaTxNum[0]_keep ;
  wire \PWM1/RemaTxNum[10]_keep ;
  wire \PWM1/RemaTxNum[11]_keep ;
  wire \PWM1/RemaTxNum[12]_keep ;
  wire \PWM1/RemaTxNum[13]_keep ;
  wire \PWM1/RemaTxNum[14]_keep ;
  wire \PWM1/RemaTxNum[15]_keep ;
  wire \PWM1/RemaTxNum[16]_keep ;
  wire \PWM1/RemaTxNum[17]_keep ;
  wire \PWM1/RemaTxNum[18]_keep ;
  wire \PWM1/RemaTxNum[19]_keep ;
  wire \PWM1/RemaTxNum[1]_keep ;
  wire \PWM1/RemaTxNum[20]_keep ;
  wire \PWM1/RemaTxNum[21]_keep ;
  wire \PWM1/RemaTxNum[22]_keep ;
  wire \PWM1/RemaTxNum[23]_keep ;
  wire \PWM1/RemaTxNum[2]_keep ;
  wire \PWM1/RemaTxNum[3]_keep ;
  wire \PWM1/RemaTxNum[4]_keep ;
  wire \PWM1/RemaTxNum[5]_keep ;
  wire \PWM1/RemaTxNum[6]_keep ;
  wire \PWM1/RemaTxNum[7]_keep ;
  wire \PWM1/RemaTxNum[8]_keep ;
  wire \PWM1/RemaTxNum[9]_keep ;
  wire \PWM1/dir_keep ;
  wire \PWM1/mux3_b0_sel_is_3_o ;
  wire \PWM1/n0_lutinv ;
  wire \PWM1/n11 ;
  wire \PWM1/n24 ;
  wire \PWM1/n25_neg_lutinv ;
  wire \PWM1/pnumr[0]_keep ;
  wire \PWM1/pnumr[10]_keep ;
  wire \PWM1/pnumr[11]_keep ;
  wire \PWM1/pnumr[12]_keep ;
  wire \PWM1/pnumr[13]_keep ;
  wire \PWM1/pnumr[14]_keep ;
  wire \PWM1/pnumr[15]_keep ;
  wire \PWM1/pnumr[16]_keep ;
  wire \PWM1/pnumr[17]_keep ;
  wire \PWM1/pnumr[18]_keep ;
  wire \PWM1/pnumr[19]_keep ;
  wire \PWM1/pnumr[1]_keep ;
  wire \PWM1/pnumr[20]_keep ;
  wire \PWM1/pnumr[21]_keep ;
  wire \PWM1/pnumr[22]_keep ;
  wire \PWM1/pnumr[23]_keep ;
  wire \PWM1/pnumr[24]_keep ;
  wire \PWM1/pnumr[25]_keep ;
  wire \PWM1/pnumr[26]_keep ;
  wire \PWM1/pnumr[27]_keep ;
  wire \PWM1/pnumr[28]_keep ;
  wire \PWM1/pnumr[29]_keep ;
  wire \PWM1/pnumr[2]_keep ;
  wire \PWM1/pnumr[30]_keep ;
  wire \PWM1/pnumr[31]_keep ;
  wire \PWM1/pnumr[3]_keep ;
  wire \PWM1/pnumr[4]_keep ;
  wire \PWM1/pnumr[5]_keep ;
  wire \PWM1/pnumr[6]_keep ;
  wire \PWM1/pnumr[7]_keep ;
  wire \PWM1/pnumr[8]_keep ;
  wire \PWM1/pnumr[9]_keep ;
  wire \PWM1/pwm_keep ;
  wire \PWM1/stopreq ;  // src/OnePWM.v(14)
  wire \PWM1/stopreq_keep ;
  wire \PWM1/sub0/c11 ;
  wire \PWM1/sub0/c15 ;
  wire \PWM1/sub0/c19 ;
  wire \PWM1/sub0/c23 ;
  wire \PWM1/sub0/c3 ;
  wire \PWM1/sub0/c7 ;
  wire \PWM1/sub1/c1 ;
  wire \PWM1/sub1/c11 ;
  wire \PWM1/sub1/c13 ;
  wire \PWM1/sub1/c15 ;
  wire \PWM1/sub1/c17 ;
  wire \PWM1/sub1/c19 ;
  wire \PWM1/sub1/c21 ;
  wire \PWM1/sub1/c23 ;
  wire \PWM1/sub1/c3 ;
  wire \PWM1/sub1/c5 ;
  wire \PWM1/sub1/c7 ;
  wire \PWM1/sub1/c9 ;
  wire \PWM1/u14_sel_is_1_o ;
  wire \PWM2/RemaTxNum[0]_keep ;
  wire \PWM2/RemaTxNum[10]_keep ;
  wire \PWM2/RemaTxNum[11]_keep ;
  wire \PWM2/RemaTxNum[12]_keep ;
  wire \PWM2/RemaTxNum[13]_keep ;
  wire \PWM2/RemaTxNum[14]_keep ;
  wire \PWM2/RemaTxNum[15]_keep ;
  wire \PWM2/RemaTxNum[16]_keep ;
  wire \PWM2/RemaTxNum[17]_keep ;
  wire \PWM2/RemaTxNum[18]_keep ;
  wire \PWM2/RemaTxNum[19]_keep ;
  wire \PWM2/RemaTxNum[1]_keep ;
  wire \PWM2/RemaTxNum[20]_keep ;
  wire \PWM2/RemaTxNum[21]_keep ;
  wire \PWM2/RemaTxNum[22]_keep ;
  wire \PWM2/RemaTxNum[23]_keep ;
  wire \PWM2/RemaTxNum[2]_keep ;
  wire \PWM2/RemaTxNum[3]_keep ;
  wire \PWM2/RemaTxNum[4]_keep ;
  wire \PWM2/RemaTxNum[5]_keep ;
  wire \PWM2/RemaTxNum[6]_keep ;
  wire \PWM2/RemaTxNum[7]_keep ;
  wire \PWM2/RemaTxNum[8]_keep ;
  wire \PWM2/RemaTxNum[9]_keep ;
  wire \PWM2/dir_keep ;
  wire \PWM2/mux3_b0_sel_is_3_o ;
  wire \PWM2/n0_lutinv ;
  wire \PWM2/n11 ;
  wire \PWM2/n24 ;
  wire \PWM2/n25_neg_lutinv ;
  wire \PWM2/pnumr[0]_keep ;
  wire \PWM2/pnumr[10]_keep ;
  wire \PWM2/pnumr[11]_keep ;
  wire \PWM2/pnumr[12]_keep ;
  wire \PWM2/pnumr[13]_keep ;
  wire \PWM2/pnumr[14]_keep ;
  wire \PWM2/pnumr[15]_keep ;
  wire \PWM2/pnumr[16]_keep ;
  wire \PWM2/pnumr[17]_keep ;
  wire \PWM2/pnumr[18]_keep ;
  wire \PWM2/pnumr[19]_keep ;
  wire \PWM2/pnumr[1]_keep ;
  wire \PWM2/pnumr[20]_keep ;
  wire \PWM2/pnumr[21]_keep ;
  wire \PWM2/pnumr[22]_keep ;
  wire \PWM2/pnumr[23]_keep ;
  wire \PWM2/pnumr[24]_keep ;
  wire \PWM2/pnumr[25]_keep ;
  wire \PWM2/pnumr[26]_keep ;
  wire \PWM2/pnumr[27]_keep ;
  wire \PWM2/pnumr[28]_keep ;
  wire \PWM2/pnumr[29]_keep ;
  wire \PWM2/pnumr[2]_keep ;
  wire \PWM2/pnumr[30]_keep ;
  wire \PWM2/pnumr[31]_keep ;
  wire \PWM2/pnumr[3]_keep ;
  wire \PWM2/pnumr[4]_keep ;
  wire \PWM2/pnumr[5]_keep ;
  wire \PWM2/pnumr[6]_keep ;
  wire \PWM2/pnumr[7]_keep ;
  wire \PWM2/pnumr[8]_keep ;
  wire \PWM2/pnumr[9]_keep ;
  wire \PWM2/pwm_keep ;
  wire \PWM2/stopreq ;  // src/OnePWM.v(14)
  wire \PWM2/stopreq_keep ;
  wire \PWM2/sub0/c11 ;
  wire \PWM2/sub0/c15 ;
  wire \PWM2/sub0/c19 ;
  wire \PWM2/sub0/c23 ;
  wire \PWM2/sub0/c3 ;
  wire \PWM2/sub0/c7 ;
  wire \PWM2/sub1/c1 ;
  wire \PWM2/sub1/c11 ;
  wire \PWM2/sub1/c13 ;
  wire \PWM2/sub1/c15 ;
  wire \PWM2/sub1/c17 ;
  wire \PWM2/sub1/c19 ;
  wire \PWM2/sub1/c21 ;
  wire \PWM2/sub1/c23 ;
  wire \PWM2/sub1/c3 ;
  wire \PWM2/sub1/c5 ;
  wire \PWM2/sub1/c7 ;
  wire \PWM2/sub1/c9 ;
  wire \PWM2/u14_sel_is_1_o ;
  wire \PWM3/RemaTxNum[0]_keep ;
  wire \PWM3/RemaTxNum[10]_keep ;
  wire \PWM3/RemaTxNum[11]_keep ;
  wire \PWM3/RemaTxNum[12]_keep ;
  wire \PWM3/RemaTxNum[13]_keep ;
  wire \PWM3/RemaTxNum[14]_keep ;
  wire \PWM3/RemaTxNum[15]_keep ;
  wire \PWM3/RemaTxNum[16]_keep ;
  wire \PWM3/RemaTxNum[17]_keep ;
  wire \PWM3/RemaTxNum[18]_keep ;
  wire \PWM3/RemaTxNum[19]_keep ;
  wire \PWM3/RemaTxNum[1]_keep ;
  wire \PWM3/RemaTxNum[20]_keep ;
  wire \PWM3/RemaTxNum[21]_keep ;
  wire \PWM3/RemaTxNum[22]_keep ;
  wire \PWM3/RemaTxNum[23]_keep ;
  wire \PWM3/RemaTxNum[2]_keep ;
  wire \PWM3/RemaTxNum[3]_keep ;
  wire \PWM3/RemaTxNum[4]_keep ;
  wire \PWM3/RemaTxNum[5]_keep ;
  wire \PWM3/RemaTxNum[6]_keep ;
  wire \PWM3/RemaTxNum[7]_keep ;
  wire \PWM3/RemaTxNum[8]_keep ;
  wire \PWM3/RemaTxNum[9]_keep ;
  wire \PWM3/dir_keep ;
  wire \PWM3/mux3_b0_sel_is_3_o ;
  wire \PWM3/n0_lutinv ;
  wire \PWM3/n11 ;
  wire \PWM3/n24 ;
  wire \PWM3/n25_neg_lutinv ;
  wire \PWM3/pnumr[0]_keep ;
  wire \PWM3/pnumr[10]_keep ;
  wire \PWM3/pnumr[11]_keep ;
  wire \PWM3/pnumr[12]_keep ;
  wire \PWM3/pnumr[13]_keep ;
  wire \PWM3/pnumr[14]_keep ;
  wire \PWM3/pnumr[15]_keep ;
  wire \PWM3/pnumr[16]_keep ;
  wire \PWM3/pnumr[17]_keep ;
  wire \PWM3/pnumr[18]_keep ;
  wire \PWM3/pnumr[19]_keep ;
  wire \PWM3/pnumr[1]_keep ;
  wire \PWM3/pnumr[20]_keep ;
  wire \PWM3/pnumr[21]_keep ;
  wire \PWM3/pnumr[22]_keep ;
  wire \PWM3/pnumr[23]_keep ;
  wire \PWM3/pnumr[24]_keep ;
  wire \PWM3/pnumr[25]_keep ;
  wire \PWM3/pnumr[26]_keep ;
  wire \PWM3/pnumr[27]_keep ;
  wire \PWM3/pnumr[28]_keep ;
  wire \PWM3/pnumr[29]_keep ;
  wire \PWM3/pnumr[2]_keep ;
  wire \PWM3/pnumr[30]_keep ;
  wire \PWM3/pnumr[31]_keep ;
  wire \PWM3/pnumr[3]_keep ;
  wire \PWM3/pnumr[4]_keep ;
  wire \PWM3/pnumr[5]_keep ;
  wire \PWM3/pnumr[6]_keep ;
  wire \PWM3/pnumr[7]_keep ;
  wire \PWM3/pnumr[8]_keep ;
  wire \PWM3/pnumr[9]_keep ;
  wire \PWM3/pwm_keep ;
  wire \PWM3/stopreq ;  // src/OnePWM.v(14)
  wire \PWM3/stopreq_keep ;
  wire \PWM3/sub0/c11 ;
  wire \PWM3/sub0/c15 ;
  wire \PWM3/sub0/c19 ;
  wire \PWM3/sub0/c23 ;
  wire \PWM3/sub0/c3 ;
  wire \PWM3/sub0/c7 ;
  wire \PWM3/sub1/c1 ;
  wire \PWM3/sub1/c11 ;
  wire \PWM3/sub1/c13 ;
  wire \PWM3/sub1/c15 ;
  wire \PWM3/sub1/c17 ;
  wire \PWM3/sub1/c19 ;
  wire \PWM3/sub1/c21 ;
  wire \PWM3/sub1/c23 ;
  wire \PWM3/sub1/c3 ;
  wire \PWM3/sub1/c5 ;
  wire \PWM3/sub1/c7 ;
  wire \PWM3/sub1/c9 ;
  wire \PWM3/u14_sel_is_1_o ;
  wire \PWM4/RemaTxNum[0]_keep ;
  wire \PWM4/RemaTxNum[10]_keep ;
  wire \PWM4/RemaTxNum[11]_keep ;
  wire \PWM4/RemaTxNum[12]_keep ;
  wire \PWM4/RemaTxNum[13]_keep ;
  wire \PWM4/RemaTxNum[14]_keep ;
  wire \PWM4/RemaTxNum[15]_keep ;
  wire \PWM4/RemaTxNum[16]_keep ;
  wire \PWM4/RemaTxNum[17]_keep ;
  wire \PWM4/RemaTxNum[18]_keep ;
  wire \PWM4/RemaTxNum[19]_keep ;
  wire \PWM4/RemaTxNum[1]_keep ;
  wire \PWM4/RemaTxNum[20]_keep ;
  wire \PWM4/RemaTxNum[21]_keep ;
  wire \PWM4/RemaTxNum[22]_keep ;
  wire \PWM4/RemaTxNum[23]_keep ;
  wire \PWM4/RemaTxNum[2]_keep ;
  wire \PWM4/RemaTxNum[3]_keep ;
  wire \PWM4/RemaTxNum[4]_keep ;
  wire \PWM4/RemaTxNum[5]_keep ;
  wire \PWM4/RemaTxNum[6]_keep ;
  wire \PWM4/RemaTxNum[7]_keep ;
  wire \PWM4/RemaTxNum[8]_keep ;
  wire \PWM4/RemaTxNum[9]_keep ;
  wire \PWM4/dir_keep ;
  wire \PWM4/mux3_b0_sel_is_3_o ;
  wire \PWM4/n0_lutinv ;
  wire \PWM4/n11 ;
  wire \PWM4/n24 ;
  wire \PWM4/n25_neg_lutinv ;
  wire \PWM4/pnumr[0]_keep ;
  wire \PWM4/pnumr[10]_keep ;
  wire \PWM4/pnumr[11]_keep ;
  wire \PWM4/pnumr[12]_keep ;
  wire \PWM4/pnumr[13]_keep ;
  wire \PWM4/pnumr[14]_keep ;
  wire \PWM4/pnumr[15]_keep ;
  wire \PWM4/pnumr[16]_keep ;
  wire \PWM4/pnumr[17]_keep ;
  wire \PWM4/pnumr[18]_keep ;
  wire \PWM4/pnumr[19]_keep ;
  wire \PWM4/pnumr[1]_keep ;
  wire \PWM4/pnumr[20]_keep ;
  wire \PWM4/pnumr[21]_keep ;
  wire \PWM4/pnumr[22]_keep ;
  wire \PWM4/pnumr[23]_keep ;
  wire \PWM4/pnumr[24]_keep ;
  wire \PWM4/pnumr[25]_keep ;
  wire \PWM4/pnumr[26]_keep ;
  wire \PWM4/pnumr[27]_keep ;
  wire \PWM4/pnumr[28]_keep ;
  wire \PWM4/pnumr[29]_keep ;
  wire \PWM4/pnumr[2]_keep ;
  wire \PWM4/pnumr[30]_keep ;
  wire \PWM4/pnumr[31]_keep ;
  wire \PWM4/pnumr[3]_keep ;
  wire \PWM4/pnumr[4]_keep ;
  wire \PWM4/pnumr[5]_keep ;
  wire \PWM4/pnumr[6]_keep ;
  wire \PWM4/pnumr[7]_keep ;
  wire \PWM4/pnumr[8]_keep ;
  wire \PWM4/pnumr[9]_keep ;
  wire \PWM4/pwm_keep ;
  wire \PWM4/stopreq ;  // src/OnePWM.v(14)
  wire \PWM4/stopreq_keep ;
  wire \PWM4/sub0/c11 ;
  wire \PWM4/sub0/c15 ;
  wire \PWM4/sub0/c19 ;
  wire \PWM4/sub0/c23 ;
  wire \PWM4/sub0/c3 ;
  wire \PWM4/sub0/c7 ;
  wire \PWM4/sub1/c1 ;
  wire \PWM4/sub1/c11 ;
  wire \PWM4/sub1/c13 ;
  wire \PWM4/sub1/c15 ;
  wire \PWM4/sub1/c17 ;
  wire \PWM4/sub1/c19 ;
  wire \PWM4/sub1/c21 ;
  wire \PWM4/sub1/c23 ;
  wire \PWM4/sub1/c3 ;
  wire \PWM4/sub1/c5 ;
  wire \PWM4/sub1/c7 ;
  wire \PWM4/sub1/c9 ;
  wire \PWM4/u14_sel_is_1_o ;
  wire \PWM5/RemaTxNum[0]_keep ;
  wire \PWM5/RemaTxNum[10]_keep ;
  wire \PWM5/RemaTxNum[11]_keep ;
  wire \PWM5/RemaTxNum[12]_keep ;
  wire \PWM5/RemaTxNum[13]_keep ;
  wire \PWM5/RemaTxNum[14]_keep ;
  wire \PWM5/RemaTxNum[15]_keep ;
  wire \PWM5/RemaTxNum[16]_keep ;
  wire \PWM5/RemaTxNum[17]_keep ;
  wire \PWM5/RemaTxNum[18]_keep ;
  wire \PWM5/RemaTxNum[19]_keep ;
  wire \PWM5/RemaTxNum[1]_keep ;
  wire \PWM5/RemaTxNum[20]_keep ;
  wire \PWM5/RemaTxNum[21]_keep ;
  wire \PWM5/RemaTxNum[22]_keep ;
  wire \PWM5/RemaTxNum[23]_keep ;
  wire \PWM5/RemaTxNum[2]_keep ;
  wire \PWM5/RemaTxNum[3]_keep ;
  wire \PWM5/RemaTxNum[4]_keep ;
  wire \PWM5/RemaTxNum[5]_keep ;
  wire \PWM5/RemaTxNum[6]_keep ;
  wire \PWM5/RemaTxNum[7]_keep ;
  wire \PWM5/RemaTxNum[8]_keep ;
  wire \PWM5/RemaTxNum[9]_keep ;
  wire \PWM5/dir_keep ;
  wire \PWM5/mux3_b0_sel_is_3_o ;
  wire \PWM5/n0_lutinv ;
  wire \PWM5/n11 ;
  wire \PWM5/n24 ;
  wire \PWM5/n25_neg_lutinv ;
  wire \PWM5/pnumr[0]_keep ;
  wire \PWM5/pnumr[10]_keep ;
  wire \PWM5/pnumr[11]_keep ;
  wire \PWM5/pnumr[12]_keep ;
  wire \PWM5/pnumr[13]_keep ;
  wire \PWM5/pnumr[14]_keep ;
  wire \PWM5/pnumr[15]_keep ;
  wire \PWM5/pnumr[16]_keep ;
  wire \PWM5/pnumr[17]_keep ;
  wire \PWM5/pnumr[18]_keep ;
  wire \PWM5/pnumr[19]_keep ;
  wire \PWM5/pnumr[1]_keep ;
  wire \PWM5/pnumr[20]_keep ;
  wire \PWM5/pnumr[21]_keep ;
  wire \PWM5/pnumr[22]_keep ;
  wire \PWM5/pnumr[23]_keep ;
  wire \PWM5/pnumr[24]_keep ;
  wire \PWM5/pnumr[25]_keep ;
  wire \PWM5/pnumr[26]_keep ;
  wire \PWM5/pnumr[27]_keep ;
  wire \PWM5/pnumr[28]_keep ;
  wire \PWM5/pnumr[29]_keep ;
  wire \PWM5/pnumr[2]_keep ;
  wire \PWM5/pnumr[30]_keep ;
  wire \PWM5/pnumr[31]_keep ;
  wire \PWM5/pnumr[3]_keep ;
  wire \PWM5/pnumr[4]_keep ;
  wire \PWM5/pnumr[5]_keep ;
  wire \PWM5/pnumr[6]_keep ;
  wire \PWM5/pnumr[7]_keep ;
  wire \PWM5/pnumr[8]_keep ;
  wire \PWM5/pnumr[9]_keep ;
  wire \PWM5/pwm_keep ;
  wire \PWM5/stopreq ;  // src/OnePWM.v(14)
  wire \PWM5/stopreq_keep ;
  wire \PWM5/sub0/c11 ;
  wire \PWM5/sub0/c15 ;
  wire \PWM5/sub0/c19 ;
  wire \PWM5/sub0/c23 ;
  wire \PWM5/sub0/c3 ;
  wire \PWM5/sub0/c7 ;
  wire \PWM5/sub1/c1 ;
  wire \PWM5/sub1/c11 ;
  wire \PWM5/sub1/c13 ;
  wire \PWM5/sub1/c15 ;
  wire \PWM5/sub1/c17 ;
  wire \PWM5/sub1/c19 ;
  wire \PWM5/sub1/c21 ;
  wire \PWM5/sub1/c23 ;
  wire \PWM5/sub1/c3 ;
  wire \PWM5/sub1/c5 ;
  wire \PWM5/sub1/c7 ;
  wire \PWM5/sub1/c9 ;
  wire \PWM5/u14_sel_is_1_o ;
  wire \PWM6/RemaTxNum[0]_keep ;
  wire \PWM6/RemaTxNum[10]_keep ;
  wire \PWM6/RemaTxNum[11]_keep ;
  wire \PWM6/RemaTxNum[12]_keep ;
  wire \PWM6/RemaTxNum[13]_keep ;
  wire \PWM6/RemaTxNum[14]_keep ;
  wire \PWM6/RemaTxNum[15]_keep ;
  wire \PWM6/RemaTxNum[16]_keep ;
  wire \PWM6/RemaTxNum[17]_keep ;
  wire \PWM6/RemaTxNum[18]_keep ;
  wire \PWM6/RemaTxNum[19]_keep ;
  wire \PWM6/RemaTxNum[1]_keep ;
  wire \PWM6/RemaTxNum[20]_keep ;
  wire \PWM6/RemaTxNum[21]_keep ;
  wire \PWM6/RemaTxNum[22]_keep ;
  wire \PWM6/RemaTxNum[23]_keep ;
  wire \PWM6/RemaTxNum[2]_keep ;
  wire \PWM6/RemaTxNum[3]_keep ;
  wire \PWM6/RemaTxNum[4]_keep ;
  wire \PWM6/RemaTxNum[5]_keep ;
  wire \PWM6/RemaTxNum[6]_keep ;
  wire \PWM6/RemaTxNum[7]_keep ;
  wire \PWM6/RemaTxNum[8]_keep ;
  wire \PWM6/RemaTxNum[9]_keep ;
  wire \PWM6/dir_keep ;
  wire \PWM6/mux3_b0_sel_is_3_o ;
  wire \PWM6/n0_lutinv ;
  wire \PWM6/n11 ;
  wire \PWM6/n18_lutinv ;
  wire \PWM6/n24 ;
  wire \PWM6/n25_neg_lutinv ;
  wire \PWM6/pnumr[0]_keep ;
  wire \PWM6/pnumr[10]_keep ;
  wire \PWM6/pnumr[11]_keep ;
  wire \PWM6/pnumr[12]_keep ;
  wire \PWM6/pnumr[13]_keep ;
  wire \PWM6/pnumr[14]_keep ;
  wire \PWM6/pnumr[15]_keep ;
  wire \PWM6/pnumr[16]_keep ;
  wire \PWM6/pnumr[17]_keep ;
  wire \PWM6/pnumr[18]_keep ;
  wire \PWM6/pnumr[19]_keep ;
  wire \PWM6/pnumr[1]_keep ;
  wire \PWM6/pnumr[20]_keep ;
  wire \PWM6/pnumr[21]_keep ;
  wire \PWM6/pnumr[22]_keep ;
  wire \PWM6/pnumr[23]_keep ;
  wire \PWM6/pnumr[24]_keep ;
  wire \PWM6/pnumr[25]_keep ;
  wire \PWM6/pnumr[26]_keep ;
  wire \PWM6/pnumr[27]_keep ;
  wire \PWM6/pnumr[28]_keep ;
  wire \PWM6/pnumr[29]_keep ;
  wire \PWM6/pnumr[2]_keep ;
  wire \PWM6/pnumr[30]_keep ;
  wire \PWM6/pnumr[31]_keep ;
  wire \PWM6/pnumr[3]_keep ;
  wire \PWM6/pnumr[4]_keep ;
  wire \PWM6/pnumr[5]_keep ;
  wire \PWM6/pnumr[6]_keep ;
  wire \PWM6/pnumr[7]_keep ;
  wire \PWM6/pnumr[8]_keep ;
  wire \PWM6/pnumr[9]_keep ;
  wire \PWM6/pwm_keep ;
  wire \PWM6/stopreq ;  // src/OnePWM.v(14)
  wire \PWM6/stopreq_keep ;
  wire \PWM6/sub0/c11 ;
  wire \PWM6/sub0/c15 ;
  wire \PWM6/sub0/c19 ;
  wire \PWM6/sub0/c23 ;
  wire \PWM6/sub0/c3 ;
  wire \PWM6/sub0/c7 ;
  wire \PWM6/sub1/c1 ;
  wire \PWM6/sub1/c11 ;
  wire \PWM6/sub1/c13 ;
  wire \PWM6/sub1/c15 ;
  wire \PWM6/sub1/c17 ;
  wire \PWM6/sub1/c19 ;
  wire \PWM6/sub1/c21 ;
  wire \PWM6/sub1/c23 ;
  wire \PWM6/sub1/c3 ;
  wire \PWM6/sub1/c5 ;
  wire \PWM6/sub1/c7 ;
  wire \PWM6/sub1/c9 ;
  wire \PWM6/u14_sel_is_1_o ;
  wire \PWM7/RemaTxNum[0]_keep ;
  wire \PWM7/RemaTxNum[10]_keep ;
  wire \PWM7/RemaTxNum[11]_keep ;
  wire \PWM7/RemaTxNum[12]_keep ;
  wire \PWM7/RemaTxNum[13]_keep ;
  wire \PWM7/RemaTxNum[14]_keep ;
  wire \PWM7/RemaTxNum[15]_keep ;
  wire \PWM7/RemaTxNum[16]_keep ;
  wire \PWM7/RemaTxNum[17]_keep ;
  wire \PWM7/RemaTxNum[18]_keep ;
  wire \PWM7/RemaTxNum[19]_keep ;
  wire \PWM7/RemaTxNum[1]_keep ;
  wire \PWM7/RemaTxNum[20]_keep ;
  wire \PWM7/RemaTxNum[21]_keep ;
  wire \PWM7/RemaTxNum[22]_keep ;
  wire \PWM7/RemaTxNum[23]_keep ;
  wire \PWM7/RemaTxNum[2]_keep ;
  wire \PWM7/RemaTxNum[3]_keep ;
  wire \PWM7/RemaTxNum[4]_keep ;
  wire \PWM7/RemaTxNum[5]_keep ;
  wire \PWM7/RemaTxNum[6]_keep ;
  wire \PWM7/RemaTxNum[7]_keep ;
  wire \PWM7/RemaTxNum[8]_keep ;
  wire \PWM7/RemaTxNum[9]_keep ;
  wire \PWM7/dir_keep ;
  wire \PWM7/mux3_b0_sel_is_3_o ;
  wire \PWM7/n0_lutinv ;
  wire \PWM7/n11 ;
  wire \PWM7/n24 ;
  wire \PWM7/n25_neg_lutinv ;
  wire \PWM7/pnumr[0]_keep ;
  wire \PWM7/pnumr[10]_keep ;
  wire \PWM7/pnumr[11]_keep ;
  wire \PWM7/pnumr[12]_keep ;
  wire \PWM7/pnumr[13]_keep ;
  wire \PWM7/pnumr[14]_keep ;
  wire \PWM7/pnumr[15]_keep ;
  wire \PWM7/pnumr[16]_keep ;
  wire \PWM7/pnumr[17]_keep ;
  wire \PWM7/pnumr[18]_keep ;
  wire \PWM7/pnumr[19]_keep ;
  wire \PWM7/pnumr[1]_keep ;
  wire \PWM7/pnumr[20]_keep ;
  wire \PWM7/pnumr[21]_keep ;
  wire \PWM7/pnumr[22]_keep ;
  wire \PWM7/pnumr[23]_keep ;
  wire \PWM7/pnumr[24]_keep ;
  wire \PWM7/pnumr[25]_keep ;
  wire \PWM7/pnumr[26]_keep ;
  wire \PWM7/pnumr[27]_keep ;
  wire \PWM7/pnumr[28]_keep ;
  wire \PWM7/pnumr[29]_keep ;
  wire \PWM7/pnumr[2]_keep ;
  wire \PWM7/pnumr[30]_keep ;
  wire \PWM7/pnumr[31]_keep ;
  wire \PWM7/pnumr[3]_keep ;
  wire \PWM7/pnumr[4]_keep ;
  wire \PWM7/pnumr[5]_keep ;
  wire \PWM7/pnumr[6]_keep ;
  wire \PWM7/pnumr[7]_keep ;
  wire \PWM7/pnumr[8]_keep ;
  wire \PWM7/pnumr[9]_keep ;
  wire \PWM7/pwm_keep ;
  wire \PWM7/stopreq ;  // src/OnePWM.v(14)
  wire \PWM7/stopreq_keep ;
  wire \PWM7/sub0/c11 ;
  wire \PWM7/sub0/c15 ;
  wire \PWM7/sub0/c19 ;
  wire \PWM7/sub0/c23 ;
  wire \PWM7/sub0/c3 ;
  wire \PWM7/sub0/c7 ;
  wire \PWM7/sub1/c1 ;
  wire \PWM7/sub1/c11 ;
  wire \PWM7/sub1/c13 ;
  wire \PWM7/sub1/c15 ;
  wire \PWM7/sub1/c17 ;
  wire \PWM7/sub1/c19 ;
  wire \PWM7/sub1/c21 ;
  wire \PWM7/sub1/c23 ;
  wire \PWM7/sub1/c3 ;
  wire \PWM7/sub1/c5 ;
  wire \PWM7/sub1/c7 ;
  wire \PWM7/sub1/c9 ;
  wire \PWM7/u14_sel_is_1_o ;
  wire \PWM8/RemaTxNum[0]_keep ;
  wire \PWM8/RemaTxNum[10]_keep ;
  wire \PWM8/RemaTxNum[11]_keep ;
  wire \PWM8/RemaTxNum[12]_keep ;
  wire \PWM8/RemaTxNum[13]_keep ;
  wire \PWM8/RemaTxNum[14]_keep ;
  wire \PWM8/RemaTxNum[15]_keep ;
  wire \PWM8/RemaTxNum[16]_keep ;
  wire \PWM8/RemaTxNum[17]_keep ;
  wire \PWM8/RemaTxNum[18]_keep ;
  wire \PWM8/RemaTxNum[19]_keep ;
  wire \PWM8/RemaTxNum[1]_keep ;
  wire \PWM8/RemaTxNum[20]_keep ;
  wire \PWM8/RemaTxNum[21]_keep ;
  wire \PWM8/RemaTxNum[22]_keep ;
  wire \PWM8/RemaTxNum[23]_keep ;
  wire \PWM8/RemaTxNum[2]_keep ;
  wire \PWM8/RemaTxNum[3]_keep ;
  wire \PWM8/RemaTxNum[4]_keep ;
  wire \PWM8/RemaTxNum[5]_keep ;
  wire \PWM8/RemaTxNum[6]_keep ;
  wire \PWM8/RemaTxNum[7]_keep ;
  wire \PWM8/RemaTxNum[8]_keep ;
  wire \PWM8/RemaTxNum[9]_keep ;
  wire \PWM8/dir_keep ;
  wire \PWM8/mux3_b0_sel_is_3_o ;
  wire \PWM8/n0_lutinv ;
  wire \PWM8/n11 ;
  wire \PWM8/n24 ;
  wire \PWM8/n25_neg_lutinv ;
  wire \PWM8/pnumr[0]_keep ;
  wire \PWM8/pnumr[10]_keep ;
  wire \PWM8/pnumr[11]_keep ;
  wire \PWM8/pnumr[12]_keep ;
  wire \PWM8/pnumr[13]_keep ;
  wire \PWM8/pnumr[14]_keep ;
  wire \PWM8/pnumr[15]_keep ;
  wire \PWM8/pnumr[16]_keep ;
  wire \PWM8/pnumr[17]_keep ;
  wire \PWM8/pnumr[18]_keep ;
  wire \PWM8/pnumr[19]_keep ;
  wire \PWM8/pnumr[1]_keep ;
  wire \PWM8/pnumr[20]_keep ;
  wire \PWM8/pnumr[21]_keep ;
  wire \PWM8/pnumr[22]_keep ;
  wire \PWM8/pnumr[23]_keep ;
  wire \PWM8/pnumr[24]_keep ;
  wire \PWM8/pnumr[25]_keep ;
  wire \PWM8/pnumr[26]_keep ;
  wire \PWM8/pnumr[27]_keep ;
  wire \PWM8/pnumr[28]_keep ;
  wire \PWM8/pnumr[29]_keep ;
  wire \PWM8/pnumr[2]_keep ;
  wire \PWM8/pnumr[30]_keep ;
  wire \PWM8/pnumr[31]_keep ;
  wire \PWM8/pnumr[3]_keep ;
  wire \PWM8/pnumr[4]_keep ;
  wire \PWM8/pnumr[5]_keep ;
  wire \PWM8/pnumr[6]_keep ;
  wire \PWM8/pnumr[7]_keep ;
  wire \PWM8/pnumr[8]_keep ;
  wire \PWM8/pnumr[9]_keep ;
  wire \PWM8/pwm_keep ;
  wire \PWM8/stopreq ;  // src/OnePWM.v(14)
  wire \PWM8/stopreq_keep ;
  wire \PWM8/sub0/c11 ;
  wire \PWM8/sub0/c15 ;
  wire \PWM8/sub0/c19 ;
  wire \PWM8/sub0/c23 ;
  wire \PWM8/sub0/c3 ;
  wire \PWM8/sub0/c7 ;
  wire \PWM8/sub1/c1 ;
  wire \PWM8/sub1/c11 ;
  wire \PWM8/sub1/c13 ;
  wire \PWM8/sub1/c15 ;
  wire \PWM8/sub1/c17 ;
  wire \PWM8/sub1/c19 ;
  wire \PWM8/sub1/c21 ;
  wire \PWM8/sub1/c23 ;
  wire \PWM8/sub1/c3 ;
  wire \PWM8/sub1/c5 ;
  wire \PWM8/sub1/c7 ;
  wire \PWM8/sub1/c9 ;
  wire \PWM8/u14_sel_is_1_o ;
  wire \PWM9/RemaTxNum[0]_keep ;
  wire \PWM9/RemaTxNum[10]_keep ;
  wire \PWM9/RemaTxNum[11]_keep ;
  wire \PWM9/RemaTxNum[12]_keep ;
  wire \PWM9/RemaTxNum[13]_keep ;
  wire \PWM9/RemaTxNum[14]_keep ;
  wire \PWM9/RemaTxNum[15]_keep ;
  wire \PWM9/RemaTxNum[16]_keep ;
  wire \PWM9/RemaTxNum[17]_keep ;
  wire \PWM9/RemaTxNum[18]_keep ;
  wire \PWM9/RemaTxNum[19]_keep ;
  wire \PWM9/RemaTxNum[1]_keep ;
  wire \PWM9/RemaTxNum[20]_keep ;
  wire \PWM9/RemaTxNum[21]_keep ;
  wire \PWM9/RemaTxNum[22]_keep ;
  wire \PWM9/RemaTxNum[23]_keep ;
  wire \PWM9/RemaTxNum[2]_keep ;
  wire \PWM9/RemaTxNum[3]_keep ;
  wire \PWM9/RemaTxNum[4]_keep ;
  wire \PWM9/RemaTxNum[5]_keep ;
  wire \PWM9/RemaTxNum[6]_keep ;
  wire \PWM9/RemaTxNum[7]_keep ;
  wire \PWM9/RemaTxNum[8]_keep ;
  wire \PWM9/RemaTxNum[9]_keep ;
  wire \PWM9/dir_keep ;
  wire \PWM9/mux3_b0_sel_is_3_o ;
  wire \PWM9/n0_lutinv ;
  wire \PWM9/n11 ;
  wire \PWM9/n24 ;
  wire \PWM9/n25_neg_lutinv ;
  wire \PWM9/pnumr[0]_keep ;
  wire \PWM9/pnumr[10]_keep ;
  wire \PWM9/pnumr[11]_keep ;
  wire \PWM9/pnumr[12]_keep ;
  wire \PWM9/pnumr[13]_keep ;
  wire \PWM9/pnumr[14]_keep ;
  wire \PWM9/pnumr[15]_keep ;
  wire \PWM9/pnumr[16]_keep ;
  wire \PWM9/pnumr[17]_keep ;
  wire \PWM9/pnumr[18]_keep ;
  wire \PWM9/pnumr[19]_keep ;
  wire \PWM9/pnumr[1]_keep ;
  wire \PWM9/pnumr[20]_keep ;
  wire \PWM9/pnumr[21]_keep ;
  wire \PWM9/pnumr[22]_keep ;
  wire \PWM9/pnumr[23]_keep ;
  wire \PWM9/pnumr[24]_keep ;
  wire \PWM9/pnumr[25]_keep ;
  wire \PWM9/pnumr[26]_keep ;
  wire \PWM9/pnumr[27]_keep ;
  wire \PWM9/pnumr[28]_keep ;
  wire \PWM9/pnumr[29]_keep ;
  wire \PWM9/pnumr[2]_keep ;
  wire \PWM9/pnumr[30]_keep ;
  wire \PWM9/pnumr[31]_keep ;
  wire \PWM9/pnumr[3]_keep ;
  wire \PWM9/pnumr[4]_keep ;
  wire \PWM9/pnumr[5]_keep ;
  wire \PWM9/pnumr[6]_keep ;
  wire \PWM9/pnumr[7]_keep ;
  wire \PWM9/pnumr[8]_keep ;
  wire \PWM9/pnumr[9]_keep ;
  wire \PWM9/pwm_keep ;
  wire \PWM9/stopreq ;  // src/OnePWM.v(14)
  wire \PWM9/stopreq_keep ;
  wire \PWM9/sub0/c11 ;
  wire \PWM9/sub0/c15 ;
  wire \PWM9/sub0/c19 ;
  wire \PWM9/sub0/c23 ;
  wire \PWM9/sub0/c3 ;
  wire \PWM9/sub0/c7 ;
  wire \PWM9/sub1/c1 ;
  wire \PWM9/sub1/c11 ;
  wire \PWM9/sub1/c13 ;
  wire \PWM9/sub1/c15 ;
  wire \PWM9/sub1/c17 ;
  wire \PWM9/sub1/c19 ;
  wire \PWM9/sub1/c21 ;
  wire \PWM9/sub1/c23 ;
  wire \PWM9/sub1/c3 ;
  wire \PWM9/sub1/c5 ;
  wire \PWM9/sub1/c7 ;
  wire \PWM9/sub1/c9 ;
  wire \PWM9/u14_sel_is_1_o ;
  wire \PWMA/RemaTxNum[0]_keep ;
  wire \PWMA/RemaTxNum[10]_keep ;
  wire \PWMA/RemaTxNum[11]_keep ;
  wire \PWMA/RemaTxNum[12]_keep ;
  wire \PWMA/RemaTxNum[13]_keep ;
  wire \PWMA/RemaTxNum[14]_keep ;
  wire \PWMA/RemaTxNum[15]_keep ;
  wire \PWMA/RemaTxNum[16]_keep ;
  wire \PWMA/RemaTxNum[17]_keep ;
  wire \PWMA/RemaTxNum[18]_keep ;
  wire \PWMA/RemaTxNum[19]_keep ;
  wire \PWMA/RemaTxNum[1]_keep ;
  wire \PWMA/RemaTxNum[20]_keep ;
  wire \PWMA/RemaTxNum[21]_keep ;
  wire \PWMA/RemaTxNum[22]_keep ;
  wire \PWMA/RemaTxNum[23]_keep ;
  wire \PWMA/RemaTxNum[2]_keep ;
  wire \PWMA/RemaTxNum[3]_keep ;
  wire \PWMA/RemaTxNum[4]_keep ;
  wire \PWMA/RemaTxNum[5]_keep ;
  wire \PWMA/RemaTxNum[6]_keep ;
  wire \PWMA/RemaTxNum[7]_keep ;
  wire \PWMA/RemaTxNum[8]_keep ;
  wire \PWMA/RemaTxNum[9]_keep ;
  wire \PWMA/dir_keep ;
  wire \PWMA/mux3_b0_sel_is_3_o ;
  wire \PWMA/n0_lutinv ;
  wire \PWMA/n11 ;
  wire \PWMA/n24 ;
  wire \PWMA/n25_neg_lutinv ;
  wire \PWMA/pnumr[0]_keep ;
  wire \PWMA/pnumr[10]_keep ;
  wire \PWMA/pnumr[11]_keep ;
  wire \PWMA/pnumr[12]_keep ;
  wire \PWMA/pnumr[13]_keep ;
  wire \PWMA/pnumr[14]_keep ;
  wire \PWMA/pnumr[15]_keep ;
  wire \PWMA/pnumr[16]_keep ;
  wire \PWMA/pnumr[17]_keep ;
  wire \PWMA/pnumr[18]_keep ;
  wire \PWMA/pnumr[19]_keep ;
  wire \PWMA/pnumr[1]_keep ;
  wire \PWMA/pnumr[20]_keep ;
  wire \PWMA/pnumr[21]_keep ;
  wire \PWMA/pnumr[22]_keep ;
  wire \PWMA/pnumr[23]_keep ;
  wire \PWMA/pnumr[24]_keep ;
  wire \PWMA/pnumr[25]_keep ;
  wire \PWMA/pnumr[26]_keep ;
  wire \PWMA/pnumr[27]_keep ;
  wire \PWMA/pnumr[28]_keep ;
  wire \PWMA/pnumr[29]_keep ;
  wire \PWMA/pnumr[2]_keep ;
  wire \PWMA/pnumr[30]_keep ;
  wire \PWMA/pnumr[31]_keep ;
  wire \PWMA/pnumr[3]_keep ;
  wire \PWMA/pnumr[4]_keep ;
  wire \PWMA/pnumr[5]_keep ;
  wire \PWMA/pnumr[6]_keep ;
  wire \PWMA/pnumr[7]_keep ;
  wire \PWMA/pnumr[8]_keep ;
  wire \PWMA/pnumr[9]_keep ;
  wire \PWMA/pwm_keep ;
  wire \PWMA/stopreq ;  // src/OnePWM.v(14)
  wire \PWMA/stopreq_keep ;
  wire \PWMA/sub0/c11 ;
  wire \PWMA/sub0/c15 ;
  wire \PWMA/sub0/c19 ;
  wire \PWMA/sub0/c23 ;
  wire \PWMA/sub0/c3 ;
  wire \PWMA/sub0/c7 ;
  wire \PWMA/sub1/c1 ;
  wire \PWMA/sub1/c11 ;
  wire \PWMA/sub1/c13 ;
  wire \PWMA/sub1/c15 ;
  wire \PWMA/sub1/c17 ;
  wire \PWMA/sub1/c19 ;
  wire \PWMA/sub1/c21 ;
  wire \PWMA/sub1/c23 ;
  wire \PWMA/sub1/c3 ;
  wire \PWMA/sub1/c5 ;
  wire \PWMA/sub1/c7 ;
  wire \PWMA/sub1/c9 ;
  wire \PWMA/u14_sel_is_1_o ;
  wire \PWMB/RemaTxNum[0]_keep ;
  wire \PWMB/RemaTxNum[10]_keep ;
  wire \PWMB/RemaTxNum[11]_keep ;
  wire \PWMB/RemaTxNum[12]_keep ;
  wire \PWMB/RemaTxNum[13]_keep ;
  wire \PWMB/RemaTxNum[14]_keep ;
  wire \PWMB/RemaTxNum[15]_keep ;
  wire \PWMB/RemaTxNum[16]_keep ;
  wire \PWMB/RemaTxNum[17]_keep ;
  wire \PWMB/RemaTxNum[18]_keep ;
  wire \PWMB/RemaTxNum[19]_keep ;
  wire \PWMB/RemaTxNum[1]_keep ;
  wire \PWMB/RemaTxNum[20]_keep ;
  wire \PWMB/RemaTxNum[21]_keep ;
  wire \PWMB/RemaTxNum[22]_keep ;
  wire \PWMB/RemaTxNum[23]_keep ;
  wire \PWMB/RemaTxNum[2]_keep ;
  wire \PWMB/RemaTxNum[3]_keep ;
  wire \PWMB/RemaTxNum[4]_keep ;
  wire \PWMB/RemaTxNum[5]_keep ;
  wire \PWMB/RemaTxNum[6]_keep ;
  wire \PWMB/RemaTxNum[7]_keep ;
  wire \PWMB/RemaTxNum[8]_keep ;
  wire \PWMB/RemaTxNum[9]_keep ;
  wire \PWMB/dir_keep ;
  wire \PWMB/mux3_b0_sel_is_3_o ;
  wire \PWMB/n0_lutinv ;
  wire \PWMB/n11 ;
  wire \PWMB/n24 ;
  wire \PWMB/n25_neg_lutinv ;
  wire \PWMB/pnumr[0]_keep ;
  wire \PWMB/pnumr[10]_keep ;
  wire \PWMB/pnumr[11]_keep ;
  wire \PWMB/pnumr[12]_keep ;
  wire \PWMB/pnumr[13]_keep ;
  wire \PWMB/pnumr[14]_keep ;
  wire \PWMB/pnumr[15]_keep ;
  wire \PWMB/pnumr[16]_keep ;
  wire \PWMB/pnumr[17]_keep ;
  wire \PWMB/pnumr[18]_keep ;
  wire \PWMB/pnumr[19]_keep ;
  wire \PWMB/pnumr[1]_keep ;
  wire \PWMB/pnumr[20]_keep ;
  wire \PWMB/pnumr[21]_keep ;
  wire \PWMB/pnumr[22]_keep ;
  wire \PWMB/pnumr[23]_keep ;
  wire \PWMB/pnumr[24]_keep ;
  wire \PWMB/pnumr[25]_keep ;
  wire \PWMB/pnumr[26]_keep ;
  wire \PWMB/pnumr[27]_keep ;
  wire \PWMB/pnumr[28]_keep ;
  wire \PWMB/pnumr[29]_keep ;
  wire \PWMB/pnumr[2]_keep ;
  wire \PWMB/pnumr[30]_keep ;
  wire \PWMB/pnumr[31]_keep ;
  wire \PWMB/pnumr[3]_keep ;
  wire \PWMB/pnumr[4]_keep ;
  wire \PWMB/pnumr[5]_keep ;
  wire \PWMB/pnumr[6]_keep ;
  wire \PWMB/pnumr[7]_keep ;
  wire \PWMB/pnumr[8]_keep ;
  wire \PWMB/pnumr[9]_keep ;
  wire \PWMB/pwm_keep ;
  wire \PWMB/stopreq ;  // src/OnePWM.v(14)
  wire \PWMB/stopreq_keep ;
  wire \PWMB/sub0/c11 ;
  wire \PWMB/sub0/c15 ;
  wire \PWMB/sub0/c19 ;
  wire \PWMB/sub0/c23 ;
  wire \PWMB/sub0/c3 ;
  wire \PWMB/sub0/c7 ;
  wire \PWMB/sub1/c1 ;
  wire \PWMB/sub1/c11 ;
  wire \PWMB/sub1/c13 ;
  wire \PWMB/sub1/c15 ;
  wire \PWMB/sub1/c17 ;
  wire \PWMB/sub1/c19 ;
  wire \PWMB/sub1/c21 ;
  wire \PWMB/sub1/c23 ;
  wire \PWMB/sub1/c3 ;
  wire \PWMB/sub1/c5 ;
  wire \PWMB/sub1/c7 ;
  wire \PWMB/sub1/c9 ;
  wire \PWMB/u14_sel_is_1_o ;
  wire \PWMC/RemaTxNum[0]_keep ;
  wire \PWMC/RemaTxNum[10]_keep ;
  wire \PWMC/RemaTxNum[11]_keep ;
  wire \PWMC/RemaTxNum[12]_keep ;
  wire \PWMC/RemaTxNum[13]_keep ;
  wire \PWMC/RemaTxNum[14]_keep ;
  wire \PWMC/RemaTxNum[15]_keep ;
  wire \PWMC/RemaTxNum[16]_keep ;
  wire \PWMC/RemaTxNum[17]_keep ;
  wire \PWMC/RemaTxNum[18]_keep ;
  wire \PWMC/RemaTxNum[19]_keep ;
  wire \PWMC/RemaTxNum[1]_keep ;
  wire \PWMC/RemaTxNum[20]_keep ;
  wire \PWMC/RemaTxNum[21]_keep ;
  wire \PWMC/RemaTxNum[22]_keep ;
  wire \PWMC/RemaTxNum[23]_keep ;
  wire \PWMC/RemaTxNum[2]_keep ;
  wire \PWMC/RemaTxNum[3]_keep ;
  wire \PWMC/RemaTxNum[4]_keep ;
  wire \PWMC/RemaTxNum[5]_keep ;
  wire \PWMC/RemaTxNum[6]_keep ;
  wire \PWMC/RemaTxNum[7]_keep ;
  wire \PWMC/RemaTxNum[8]_keep ;
  wire \PWMC/RemaTxNum[9]_keep ;
  wire \PWMC/dir_keep ;
  wire \PWMC/mux3_b0_sel_is_3_o ;
  wire \PWMC/n0_lutinv ;
  wire \PWMC/n11 ;
  wire \PWMC/n24 ;
  wire \PWMC/n25_neg_lutinv ;
  wire \PWMC/pnumr[0]_keep ;
  wire \PWMC/pnumr[10]_keep ;
  wire \PWMC/pnumr[11]_keep ;
  wire \PWMC/pnumr[12]_keep ;
  wire \PWMC/pnumr[13]_keep ;
  wire \PWMC/pnumr[14]_keep ;
  wire \PWMC/pnumr[15]_keep ;
  wire \PWMC/pnumr[16]_keep ;
  wire \PWMC/pnumr[17]_keep ;
  wire \PWMC/pnumr[18]_keep ;
  wire \PWMC/pnumr[19]_keep ;
  wire \PWMC/pnumr[1]_keep ;
  wire \PWMC/pnumr[20]_keep ;
  wire \PWMC/pnumr[21]_keep ;
  wire \PWMC/pnumr[22]_keep ;
  wire \PWMC/pnumr[23]_keep ;
  wire \PWMC/pnumr[24]_keep ;
  wire \PWMC/pnumr[25]_keep ;
  wire \PWMC/pnumr[26]_keep ;
  wire \PWMC/pnumr[27]_keep ;
  wire \PWMC/pnumr[28]_keep ;
  wire \PWMC/pnumr[29]_keep ;
  wire \PWMC/pnumr[2]_keep ;
  wire \PWMC/pnumr[30]_keep ;
  wire \PWMC/pnumr[31]_keep ;
  wire \PWMC/pnumr[3]_keep ;
  wire \PWMC/pnumr[4]_keep ;
  wire \PWMC/pnumr[5]_keep ;
  wire \PWMC/pnumr[6]_keep ;
  wire \PWMC/pnumr[7]_keep ;
  wire \PWMC/pnumr[8]_keep ;
  wire \PWMC/pnumr[9]_keep ;
  wire \PWMC/pwm_keep ;
  wire \PWMC/stopreq ;  // src/OnePWM.v(14)
  wire \PWMC/stopreq_keep ;
  wire \PWMC/sub0/c11 ;
  wire \PWMC/sub0/c15 ;
  wire \PWMC/sub0/c19 ;
  wire \PWMC/sub0/c23 ;
  wire \PWMC/sub0/c3 ;
  wire \PWMC/sub0/c7 ;
  wire \PWMC/sub1/c1 ;
  wire \PWMC/sub1/c11 ;
  wire \PWMC/sub1/c13 ;
  wire \PWMC/sub1/c15 ;
  wire \PWMC/sub1/c17 ;
  wire \PWMC/sub1/c19 ;
  wire \PWMC/sub1/c21 ;
  wire \PWMC/sub1/c23 ;
  wire \PWMC/sub1/c3 ;
  wire \PWMC/sub1/c5 ;
  wire \PWMC/sub1/c7 ;
  wire \PWMC/sub1/c9 ;
  wire \PWMC/u14_sel_is_1_o ;
  wire \PWMD/RemaTxNum[0]_keep ;
  wire \PWMD/RemaTxNum[10]_keep ;
  wire \PWMD/RemaTxNum[11]_keep ;
  wire \PWMD/RemaTxNum[12]_keep ;
  wire \PWMD/RemaTxNum[13]_keep ;
  wire \PWMD/RemaTxNum[14]_keep ;
  wire \PWMD/RemaTxNum[15]_keep ;
  wire \PWMD/RemaTxNum[16]_keep ;
  wire \PWMD/RemaTxNum[17]_keep ;
  wire \PWMD/RemaTxNum[18]_keep ;
  wire \PWMD/RemaTxNum[19]_keep ;
  wire \PWMD/RemaTxNum[1]_keep ;
  wire \PWMD/RemaTxNum[20]_keep ;
  wire \PWMD/RemaTxNum[21]_keep ;
  wire \PWMD/RemaTxNum[22]_keep ;
  wire \PWMD/RemaTxNum[23]_keep ;
  wire \PWMD/RemaTxNum[2]_keep ;
  wire \PWMD/RemaTxNum[3]_keep ;
  wire \PWMD/RemaTxNum[4]_keep ;
  wire \PWMD/RemaTxNum[5]_keep ;
  wire \PWMD/RemaTxNum[6]_keep ;
  wire \PWMD/RemaTxNum[7]_keep ;
  wire \PWMD/RemaTxNum[8]_keep ;
  wire \PWMD/RemaTxNum[9]_keep ;
  wire \PWMD/dir_keep ;
  wire \PWMD/mux3_b0_sel_is_3_o ;
  wire \PWMD/n0_lutinv ;
  wire \PWMD/n11 ;
  wire \PWMD/n24 ;
  wire \PWMD/n25_neg_lutinv ;
  wire \PWMD/pnumr[0]_keep ;
  wire \PWMD/pnumr[10]_keep ;
  wire \PWMD/pnumr[11]_keep ;
  wire \PWMD/pnumr[12]_keep ;
  wire \PWMD/pnumr[13]_keep ;
  wire \PWMD/pnumr[14]_keep ;
  wire \PWMD/pnumr[15]_keep ;
  wire \PWMD/pnumr[16]_keep ;
  wire \PWMD/pnumr[17]_keep ;
  wire \PWMD/pnumr[18]_keep ;
  wire \PWMD/pnumr[19]_keep ;
  wire \PWMD/pnumr[1]_keep ;
  wire \PWMD/pnumr[20]_keep ;
  wire \PWMD/pnumr[21]_keep ;
  wire \PWMD/pnumr[22]_keep ;
  wire \PWMD/pnumr[23]_keep ;
  wire \PWMD/pnumr[24]_keep ;
  wire \PWMD/pnumr[25]_keep ;
  wire \PWMD/pnumr[26]_keep ;
  wire \PWMD/pnumr[27]_keep ;
  wire \PWMD/pnumr[28]_keep ;
  wire \PWMD/pnumr[29]_keep ;
  wire \PWMD/pnumr[2]_keep ;
  wire \PWMD/pnumr[30]_keep ;
  wire \PWMD/pnumr[31]_keep ;
  wire \PWMD/pnumr[3]_keep ;
  wire \PWMD/pnumr[4]_keep ;
  wire \PWMD/pnumr[5]_keep ;
  wire \PWMD/pnumr[6]_keep ;
  wire \PWMD/pnumr[7]_keep ;
  wire \PWMD/pnumr[8]_keep ;
  wire \PWMD/pnumr[9]_keep ;
  wire \PWMD/pwm_keep ;
  wire \PWMD/stopreq ;  // src/OnePWM.v(14)
  wire \PWMD/stopreq_keep ;
  wire \PWMD/sub0/c11 ;
  wire \PWMD/sub0/c15 ;
  wire \PWMD/sub0/c19 ;
  wire \PWMD/sub0/c23 ;
  wire \PWMD/sub0/c3 ;
  wire \PWMD/sub0/c7 ;
  wire \PWMD/sub1/c1 ;
  wire \PWMD/sub1/c11 ;
  wire \PWMD/sub1/c13 ;
  wire \PWMD/sub1/c15 ;
  wire \PWMD/sub1/c17 ;
  wire \PWMD/sub1/c19 ;
  wire \PWMD/sub1/c21 ;
  wire \PWMD/sub1/c23 ;
  wire \PWMD/sub1/c3 ;
  wire \PWMD/sub1/c5 ;
  wire \PWMD/sub1/c7 ;
  wire \PWMD/sub1/c9 ;
  wire \PWMD/u14_sel_is_1_o ;
  wire \PWME/RemaTxNum[0]_keep ;
  wire \PWME/RemaTxNum[10]_keep ;
  wire \PWME/RemaTxNum[11]_keep ;
  wire \PWME/RemaTxNum[12]_keep ;
  wire \PWME/RemaTxNum[13]_keep ;
  wire \PWME/RemaTxNum[14]_keep ;
  wire \PWME/RemaTxNum[15]_keep ;
  wire \PWME/RemaTxNum[16]_keep ;
  wire \PWME/RemaTxNum[17]_keep ;
  wire \PWME/RemaTxNum[18]_keep ;
  wire \PWME/RemaTxNum[19]_keep ;
  wire \PWME/RemaTxNum[1]_keep ;
  wire \PWME/RemaTxNum[20]_keep ;
  wire \PWME/RemaTxNum[21]_keep ;
  wire \PWME/RemaTxNum[22]_keep ;
  wire \PWME/RemaTxNum[23]_keep ;
  wire \PWME/RemaTxNum[2]_keep ;
  wire \PWME/RemaTxNum[3]_keep ;
  wire \PWME/RemaTxNum[4]_keep ;
  wire \PWME/RemaTxNum[5]_keep ;
  wire \PWME/RemaTxNum[6]_keep ;
  wire \PWME/RemaTxNum[7]_keep ;
  wire \PWME/RemaTxNum[8]_keep ;
  wire \PWME/RemaTxNum[9]_keep ;
  wire \PWME/dir_keep ;
  wire \PWME/mux3_b0_sel_is_3_o ;
  wire \PWME/n0_lutinv ;
  wire \PWME/n11 ;
  wire \PWME/n24 ;
  wire \PWME/n25_neg_lutinv ;
  wire \PWME/pnumr[0]_keep ;
  wire \PWME/pnumr[10]_keep ;
  wire \PWME/pnumr[11]_keep ;
  wire \PWME/pnumr[12]_keep ;
  wire \PWME/pnumr[13]_keep ;
  wire \PWME/pnumr[14]_keep ;
  wire \PWME/pnumr[15]_keep ;
  wire \PWME/pnumr[16]_keep ;
  wire \PWME/pnumr[17]_keep ;
  wire \PWME/pnumr[18]_keep ;
  wire \PWME/pnumr[19]_keep ;
  wire \PWME/pnumr[1]_keep ;
  wire \PWME/pnumr[20]_keep ;
  wire \PWME/pnumr[21]_keep ;
  wire \PWME/pnumr[22]_keep ;
  wire \PWME/pnumr[23]_keep ;
  wire \PWME/pnumr[24]_keep ;
  wire \PWME/pnumr[25]_keep ;
  wire \PWME/pnumr[26]_keep ;
  wire \PWME/pnumr[27]_keep ;
  wire \PWME/pnumr[28]_keep ;
  wire \PWME/pnumr[29]_keep ;
  wire \PWME/pnumr[2]_keep ;
  wire \PWME/pnumr[30]_keep ;
  wire \PWME/pnumr[31]_keep ;
  wire \PWME/pnumr[3]_keep ;
  wire \PWME/pnumr[4]_keep ;
  wire \PWME/pnumr[5]_keep ;
  wire \PWME/pnumr[6]_keep ;
  wire \PWME/pnumr[7]_keep ;
  wire \PWME/pnumr[8]_keep ;
  wire \PWME/pnumr[9]_keep ;
  wire \PWME/pwm_keep ;
  wire \PWME/stopreq ;  // src/OnePWM.v(14)
  wire \PWME/stopreq_keep ;
  wire \PWME/sub0/c11 ;
  wire \PWME/sub0/c15 ;
  wire \PWME/sub0/c19 ;
  wire \PWME/sub0/c23 ;
  wire \PWME/sub0/c3 ;
  wire \PWME/sub0/c7 ;
  wire \PWME/sub1/c1 ;
  wire \PWME/sub1/c11 ;
  wire \PWME/sub1/c13 ;
  wire \PWME/sub1/c15 ;
  wire \PWME/sub1/c17 ;
  wire \PWME/sub1/c19 ;
  wire \PWME/sub1/c21 ;
  wire \PWME/sub1/c23 ;
  wire \PWME/sub1/c3 ;
  wire \PWME/sub1/c5 ;
  wire \PWME/sub1/c7 ;
  wire \PWME/sub1/c9 ;
  wire \PWME/u14_sel_is_1_o ;
  wire \PWMF/RemaTxNum[0]_keep ;
  wire \PWMF/RemaTxNum[10]_keep ;
  wire \PWMF/RemaTxNum[11]_keep ;
  wire \PWMF/RemaTxNum[12]_keep ;
  wire \PWMF/RemaTxNum[13]_keep ;
  wire \PWMF/RemaTxNum[14]_keep ;
  wire \PWMF/RemaTxNum[15]_keep ;
  wire \PWMF/RemaTxNum[16]_keep ;
  wire \PWMF/RemaTxNum[17]_keep ;
  wire \PWMF/RemaTxNum[18]_keep ;
  wire \PWMF/RemaTxNum[19]_keep ;
  wire \PWMF/RemaTxNum[1]_keep ;
  wire \PWMF/RemaTxNum[20]_keep ;
  wire \PWMF/RemaTxNum[21]_keep ;
  wire \PWMF/RemaTxNum[22]_keep ;
  wire \PWMF/RemaTxNum[23]_keep ;
  wire \PWMF/RemaTxNum[2]_keep ;
  wire \PWMF/RemaTxNum[3]_keep ;
  wire \PWMF/RemaTxNum[4]_keep ;
  wire \PWMF/RemaTxNum[5]_keep ;
  wire \PWMF/RemaTxNum[6]_keep ;
  wire \PWMF/RemaTxNum[7]_keep ;
  wire \PWMF/RemaTxNum[8]_keep ;
  wire \PWMF/RemaTxNum[9]_keep ;
  wire \PWMF/dir_keep ;
  wire \PWMF/mux3_b0_sel_is_3_o ;
  wire \PWMF/n0_lutinv ;
  wire \PWMF/n11 ;
  wire \PWMF/n24 ;
  wire \PWMF/n25_neg_lutinv ;
  wire \PWMF/pnumr[0]_keep ;
  wire \PWMF/pnumr[10]_keep ;
  wire \PWMF/pnumr[11]_keep ;
  wire \PWMF/pnumr[12]_keep ;
  wire \PWMF/pnumr[13]_keep ;
  wire \PWMF/pnumr[14]_keep ;
  wire \PWMF/pnumr[15]_keep ;
  wire \PWMF/pnumr[16]_keep ;
  wire \PWMF/pnumr[17]_keep ;
  wire \PWMF/pnumr[18]_keep ;
  wire \PWMF/pnumr[19]_keep ;
  wire \PWMF/pnumr[1]_keep ;
  wire \PWMF/pnumr[20]_keep ;
  wire \PWMF/pnumr[21]_keep ;
  wire \PWMF/pnumr[22]_keep ;
  wire \PWMF/pnumr[23]_keep ;
  wire \PWMF/pnumr[24]_keep ;
  wire \PWMF/pnumr[25]_keep ;
  wire \PWMF/pnumr[26]_keep ;
  wire \PWMF/pnumr[27]_keep ;
  wire \PWMF/pnumr[28]_keep ;
  wire \PWMF/pnumr[29]_keep ;
  wire \PWMF/pnumr[2]_keep ;
  wire \PWMF/pnumr[30]_keep ;
  wire \PWMF/pnumr[31]_keep ;
  wire \PWMF/pnumr[3]_keep ;
  wire \PWMF/pnumr[4]_keep ;
  wire \PWMF/pnumr[5]_keep ;
  wire \PWMF/pnumr[6]_keep ;
  wire \PWMF/pnumr[7]_keep ;
  wire \PWMF/pnumr[8]_keep ;
  wire \PWMF/pnumr[9]_keep ;
  wire \PWMF/pwm_keep ;
  wire \PWMF/stopreq ;  // src/OnePWM.v(14)
  wire \PWMF/stopreq_keep ;
  wire \PWMF/sub0/c1 ;
  wire \PWMF/sub0/c11 ;
  wire \PWMF/sub0/c13 ;
  wire \PWMF/sub0/c15 ;
  wire \PWMF/sub0/c17 ;
  wire \PWMF/sub0/c19 ;
  wire \PWMF/sub0/c21 ;
  wire \PWMF/sub0/c23 ;
  wire \PWMF/sub0/c25 ;
  wire \PWMF/sub0/c3 ;
  wire \PWMF/sub0/c5 ;
  wire \PWMF/sub0/c7 ;
  wire \PWMF/sub0/c9 ;
  wire \PWMF/sub1/c1 ;
  wire \PWMF/sub1/c11 ;
  wire \PWMF/sub1/c13 ;
  wire \PWMF/sub1/c15 ;
  wire \PWMF/sub1/c17 ;
  wire \PWMF/sub1/c19 ;
  wire \PWMF/sub1/c21 ;
  wire \PWMF/sub1/c23 ;
  wire \PWMF/sub1/c3 ;
  wire \PWMF/sub1/c5 ;
  wire \PWMF/sub1/c7 ;
  wire \PWMF/sub1/c9 ;
  wire \PWMF/u14_sel_is_1_o ;
  wire \U_AHB/h2h_hwrite ;  // src/AHB.v(22)
  wire \U_AHB/h2h_hwritew ;  // src/AHB.v(19)
  wire \U_AHB/n10 ;
  wire \U_AHB/n102 ;
  wire \U_AHB/n104_lutinv ;
  wire \U_AHB/n105 ;
  wire \U_AHB/n108 ;
  wire \U_AHB/n111 ;
  wire \U_AHB/n113_lutinv ;
  wire \U_AHB/n12 ;
  wire \U_AHB/n14 ;
  wire \U_AHB/n16 ;
  wire \U_AHB/n18 ;
  wire \U_AHB/n2 ;
  wire \U_AHB/n20 ;
  wire \U_AHB/n22 ;
  wire \U_AHB/n24 ;
  wire \U_AHB/n26 ;
  wire \U_AHB/n28 ;
  wire \U_AHB/n30 ;
  wire \U_AHB/n32 ;
  wire \U_AHB/n34 ;
  wire \U_AHB/n36 ;
  wire \U_AHB/n38 ;
  wire \U_AHB/n4 ;
  wire \U_AHB/n45 ;
  wire \U_AHB/n47 ;
  wire \U_AHB/n51 ;
  wire \U_AHB/n53 ;
  wire \U_AHB/n55 ;
  wire \U_AHB/n57 ;
  wire \U_AHB/n59 ;
  wire \U_AHB/n61 ;
  wire \U_AHB/n63 ;
  wire \U_AHB/n65 ;
  wire \U_AHB/n67 ;
  wire \U_AHB/n69 ;
  wire \U_AHB/n71 ;
  wire \U_AHB/n73 ;
  wire \U_AHB/n75 ;
  wire \U_AHB/n77 ;
  wire \U_AHB/n79 ;
  wire \U_AHB/n8 ;
  wire \U_AHB/n82 ;
  wire \U_AHB/n87 ;
  wire \U_AHB/n90 ;
  wire \U_AHB/n93 ;
  wire \U_AHB/n95_lutinv ;
  wire \U_AHB/n96 ;
  wire \U_AHB/n99 ;
  wire _al_n1_en;
  wire _al_u1030_o;
  wire _al_u1031_o;
  wire _al_u1032_o;
  wire _al_u1033_o;
  wire _al_u1034_o;
  wire _al_u1035_o;
  wire _al_u1036_o;
  wire _al_u1067_o;
  wire _al_u1068_o;
  wire _al_u1069_o;
  wire _al_u1070_o;
  wire _al_u1071_o;
  wire _al_u1072_o;
  wire _al_u1073_o;
  wire _al_u1104_o;
  wire _al_u1105_o;
  wire _al_u1106_o;
  wire _al_u1107_o;
  wire _al_u1108_o;
  wire _al_u1109_o;
  wire _al_u1110_o;
  wire _al_u1141_o;
  wire _al_u1142_o;
  wire _al_u1143_o;
  wire _al_u1144_o;
  wire _al_u1145_o;
  wire _al_u1146_o;
  wire _al_u1147_o;
  wire _al_u1178_o;
  wire _al_u1179_o;
  wire _al_u1180_o;
  wire _al_u1181_o;
  wire _al_u1182_o;
  wire _al_u1183_o;
  wire _al_u1184_o;
  wire _al_u1215_o;
  wire _al_u1216_o;
  wire _al_u1217_o;
  wire _al_u1218_o;
  wire _al_u1219_o;
  wire _al_u1220_o;
  wire _al_u1221_o;
  wire _al_u1252_o;
  wire _al_u1253_o;
  wire _al_u1254_o;
  wire _al_u1255_o;
  wire _al_u1256_o;
  wire _al_u1257_o;
  wire _al_u1258_o;
  wire _al_u1289_o;
  wire _al_u1290_o;
  wire _al_u1291_o;
  wire _al_u1292_o;
  wire _al_u1293_o;
  wire _al_u1294_o;
  wire _al_u1295_o;
  wire _al_u1360_o;
  wire _al_u1361_o;
  wire _al_u1362_o;
  wire _al_u1363_o;
  wire _al_u1364_o;
  wire _al_u1365_o;
  wire _al_u1366_o;
  wire _al_u1367_o;
  wire _al_u1368_o;
  wire _al_u1369_o;
  wire _al_u1370_o;
  wire _al_u1371_o;
  wire _al_u1372_o;
  wire _al_u1373_o;
  wire _al_u1374_o;
  wire _al_u1375_o;
  wire _al_u1376_o;
  wire _al_u1378_o;
  wire _al_u1379_o;
  wire _al_u1380_o;
  wire _al_u1381_o;
  wire _al_u1382_o;
  wire _al_u1383_o;
  wire _al_u1384_o;
  wire _al_u1385_o;
  wire _al_u1386_o;
  wire _al_u1387_o;
  wire _al_u1388_o;
  wire _al_u1389_o;
  wire _al_u1390_o;
  wire _al_u1391_o;
  wire _al_u1392_o;
  wire _al_u1393_o;
  wire _al_u1395_o;
  wire _al_u1396_o;
  wire _al_u1397_o;
  wire _al_u1398_o;
  wire _al_u1399_o;
  wire _al_u1400_o;
  wire _al_u1401_o;
  wire _al_u1402_o;
  wire _al_u1403_o;
  wire _al_u1404_o;
  wire _al_u1405_o;
  wire _al_u1406_o;
  wire _al_u1407_o;
  wire _al_u1408_o;
  wire _al_u1409_o;
  wire _al_u1410_o;
  wire _al_u1411_o;
  wire _al_u1413_o;
  wire _al_u1414_o;
  wire _al_u1415_o;
  wire _al_u1416_o;
  wire _al_u1417_o;
  wire _al_u1418_o;
  wire _al_u1419_o;
  wire _al_u1420_o;
  wire _al_u1421_o;
  wire _al_u1422_o;
  wire _al_u1423_o;
  wire _al_u1424_o;
  wire _al_u1425_o;
  wire _al_u1426_o;
  wire _al_u1427_o;
  wire _al_u1428_o;
  wire _al_u1430_o;
  wire _al_u1431_o;
  wire _al_u1432_o;
  wire _al_u1433_o;
  wire _al_u1434_o;
  wire _al_u1435_o;
  wire _al_u1436_o;
  wire _al_u1437_o;
  wire _al_u1438_o;
  wire _al_u1439_o;
  wire _al_u1440_o;
  wire _al_u1441_o;
  wire _al_u1442_o;
  wire _al_u1443_o;
  wire _al_u1444_o;
  wire _al_u1445_o;
  wire _al_u1447_o;
  wire _al_u1448_o;
  wire _al_u1449_o;
  wire _al_u1450_o;
  wire _al_u1451_o;
  wire _al_u1452_o;
  wire _al_u1453_o;
  wire _al_u1454_o;
  wire _al_u1455_o;
  wire _al_u1456_o;
  wire _al_u1457_o;
  wire _al_u1458_o;
  wire _al_u1459_o;
  wire _al_u1460_o;
  wire _al_u1461_o;
  wire _al_u1462_o;
  wire _al_u1464_o;
  wire _al_u1465_o;
  wire _al_u1466_o;
  wire _al_u1467_o;
  wire _al_u1468_o;
  wire _al_u1469_o;
  wire _al_u1470_o;
  wire _al_u1471_o;
  wire _al_u1472_o;
  wire _al_u1473_o;
  wire _al_u1474_o;
  wire _al_u1475_o;
  wire _al_u1476_o;
  wire _al_u1477_o;
  wire _al_u1480_o;
  wire _al_u1481_o;
  wire _al_u1482_o;
  wire _al_u1483_o;
  wire _al_u1484_o;
  wire _al_u1485_o;
  wire _al_u1486_o;
  wire _al_u1487_o;
  wire _al_u1488_o;
  wire _al_u1489_o;
  wire _al_u1490_o;
  wire _al_u1491_o;
  wire _al_u1492_o;
  wire _al_u1493_o;
  wire _al_u1494_o;
  wire _al_u1495_o;
  wire _al_u1496_o;
  wire _al_u1498_o;
  wire _al_u1499_o;
  wire _al_u1500_o;
  wire _al_u1501_o;
  wire _al_u1502_o;
  wire _al_u1503_o;
  wire _al_u1504_o;
  wire _al_u1505_o;
  wire _al_u1506_o;
  wire _al_u1507_o;
  wire _al_u1508_o;
  wire _al_u1509_o;
  wire _al_u1510_o;
  wire _al_u1511_o;
  wire _al_u1512_o;
  wire _al_u1513_o;
  wire _al_u1514_o;
  wire _al_u1516_o;
  wire _al_u1517_o;
  wire _al_u1518_o;
  wire _al_u1519_o;
  wire _al_u1520_o;
  wire _al_u1521_o;
  wire _al_u1522_o;
  wire _al_u1523_o;
  wire _al_u1524_o;
  wire _al_u1525_o;
  wire _al_u1526_o;
  wire _al_u1527_o;
  wire _al_u1528_o;
  wire _al_u1529_o;
  wire _al_u1530_o;
  wire _al_u1531_o;
  wire _al_u1533_o;
  wire _al_u1534_o;
  wire _al_u1535_o;
  wire _al_u1536_o;
  wire _al_u1537_o;
  wire _al_u1538_o;
  wire _al_u1539_o;
  wire _al_u1540_o;
  wire _al_u1541_o;
  wire _al_u1542_o;
  wire _al_u1543_o;
  wire _al_u1544_o;
  wire _al_u1545_o;
  wire _al_u1546_o;
  wire _al_u1547_o;
  wire _al_u1548_o;
  wire _al_u1549_o;
  wire _al_u1551_o;
  wire _al_u1552_o;
  wire _al_u1553_o;
  wire _al_u1554_o;
  wire _al_u1555_o;
  wire _al_u1556_o;
  wire _al_u1557_o;
  wire _al_u1558_o;
  wire _al_u1559_o;
  wire _al_u1560_o;
  wire _al_u1561_o;
  wire _al_u1562_o;
  wire _al_u1563_o;
  wire _al_u1564_o;
  wire _al_u1565_o;
  wire _al_u1566_o;
  wire _al_u1568_o;
  wire _al_u1569_o;
  wire _al_u1570_o;
  wire _al_u1571_o;
  wire _al_u1572_o;
  wire _al_u1573_o;
  wire _al_u1574_o;
  wire _al_u1575_o;
  wire _al_u1576_o;
  wire _al_u1577_o;
  wire _al_u1578_o;
  wire _al_u1579_o;
  wire _al_u1580_o;
  wire _al_u1581_o;
  wire _al_u1582_o;
  wire _al_u1583_o;
  wire _al_u1585_o;
  wire _al_u1586_o;
  wire _al_u1587_o;
  wire _al_u1588_o;
  wire _al_u1589_o;
  wire _al_u1590_o;
  wire _al_u1591_o;
  wire _al_u1592_o;
  wire _al_u1593_o;
  wire _al_u1594_o;
  wire _al_u1595_o;
  wire _al_u1596_o;
  wire _al_u1597_o;
  wire _al_u1598_o;
  wire _al_u1599_o;
  wire _al_u1600_o;
  wire _al_u1602_o;
  wire _al_u1603_o;
  wire _al_u1604_o;
  wire _al_u1605_o;
  wire _al_u1606_o;
  wire _al_u1607_o;
  wire _al_u1608_o;
  wire _al_u1609_o;
  wire _al_u1610_o;
  wire _al_u1611_o;
  wire _al_u1612_o;
  wire _al_u1613_o;
  wire _al_u1614_o;
  wire _al_u1615_o;
  wire _al_u1616_o;
  wire _al_u1617_o;
  wire _al_u1618_o;
  wire _al_u1620_o;
  wire _al_u1621_o;
  wire _al_u1622_o;
  wire _al_u1623_o;
  wire _al_u1624_o;
  wire _al_u1625_o;
  wire _al_u1626_o;
  wire _al_u1627_o;
  wire _al_u1628_o;
  wire _al_u1629_o;
  wire _al_u1630_o;
  wire _al_u1631_o;
  wire _al_u1632_o;
  wire _al_u1633_o;
  wire _al_u1634_o;
  wire _al_u1635_o;
  wire _al_u1636_o;
  wire _al_u1638_o;
  wire _al_u1639_o;
  wire _al_u1640_o;
  wire _al_u1641_o;
  wire _al_u1642_o;
  wire _al_u1643_o;
  wire _al_u1644_o;
  wire _al_u1645_o;
  wire _al_u1647_o;
  wire _al_u1648_o;
  wire _al_u1649_o;
  wire _al_u1650_o;
  wire _al_u1651_o;
  wire _al_u1652_o;
  wire _al_u1686_o;
  wire _al_u1687_o;
  wire _al_u1688_o;
  wire _al_u1689_o;
  wire _al_u1690_o;
  wire _al_u1691_o;
  wire _al_u1693_o;
  wire _al_u1695_o;
  wire _al_u1697_o;
  wire _al_u1699_o;
  wire _al_u1701_o;
  wire _al_u1703_o;
  wire _al_u1705_o;
  wire _al_u1707_o;
  wire _al_u1709_o;
  wire _al_u1711_o;
  wire _al_u1713_o;
  wire _al_u1715_o;
  wire _al_u1717_o;
  wire _al_u1719_o;
  wire _al_u1721_o;
  wire _al_u1723_o;
  wire _al_u1725_o;
  wire _al_u1727_o;
  wire _al_u1729_o;
  wire _al_u1731_o;
  wire _al_u1733_o;
  wire _al_u1735_o;
  wire _al_u1737_o;
  wire _al_u1739_o;
  wire _al_u1741_o;
  wire _al_u1742_o;
  wire _al_u1743_o;
  wire _al_u1744_o;
  wire _al_u1745_o;
  wire _al_u1746_o;
  wire _al_u1747_o;
  wire _al_u1748_o;
  wire _al_u1749_o;
  wire _al_u1750_o;
  wire _al_u1751_o;
  wire _al_u1752_o;
  wire _al_u1753_o;
  wire _al_u1754_o;
  wire _al_u1755_o;
  wire _al_u1756_o;
  wire _al_u1757_o;
  wire _al_u1758_o;
  wire _al_u1759_o;
  wire _al_u1760_o;
  wire _al_u1761_o;
  wire _al_u1762_o;
  wire _al_u1763_o;
  wire _al_u1764_o;
  wire _al_u1765_o;
  wire _al_u1768_o;
  wire _al_u1769_o;
  wire _al_u1770_o;
  wire _al_u1771_o;
  wire _al_u1772_o;
  wire _al_u1773_o;
  wire _al_u1775_o;
  wire _al_u1777_o;
  wire _al_u1779_o;
  wire _al_u1781_o;
  wire _al_u1783_o;
  wire _al_u1785_o;
  wire _al_u1787_o;
  wire _al_u1789_o;
  wire _al_u1791_o;
  wire _al_u1793_o;
  wire _al_u1795_o;
  wire _al_u1797_o;
  wire _al_u1799_o;
  wire _al_u1801_o;
  wire _al_u1803_o;
  wire _al_u1805_o;
  wire _al_u1807_o;
  wire _al_u1809_o;
  wire _al_u1811_o;
  wire _al_u1813_o;
  wire _al_u1815_o;
  wire _al_u1817_o;
  wire _al_u1819_o;
  wire _al_u1821_o;
  wire _al_u1823_o;
  wire _al_u1824_o;
  wire _al_u1825_o;
  wire _al_u1826_o;
  wire _al_u1827_o;
  wire _al_u1828_o;
  wire _al_u1829_o;
  wire _al_u1830_o;
  wire _al_u1831_o;
  wire _al_u1832_o;
  wire _al_u1833_o;
  wire _al_u1834_o;
  wire _al_u1835_o;
  wire _al_u1836_o;
  wire _al_u1837_o;
  wire _al_u1838_o;
  wire _al_u1839_o;
  wire _al_u1840_o;
  wire _al_u1841_o;
  wire _al_u1842_o;
  wire _al_u1843_o;
  wire _al_u1844_o;
  wire _al_u1845_o;
  wire _al_u1846_o;
  wire _al_u1847_o;
  wire _al_u1850_o;
  wire _al_u1851_o;
  wire _al_u1852_o;
  wire _al_u1853_o;
  wire _al_u1854_o;
  wire _al_u1855_o;
  wire _al_u1857_o;
  wire _al_u1859_o;
  wire _al_u1861_o;
  wire _al_u1863_o;
  wire _al_u1865_o;
  wire _al_u1867_o;
  wire _al_u1869_o;
  wire _al_u1871_o;
  wire _al_u1873_o;
  wire _al_u1875_o;
  wire _al_u1877_o;
  wire _al_u1879_o;
  wire _al_u1881_o;
  wire _al_u1883_o;
  wire _al_u1885_o;
  wire _al_u1887_o;
  wire _al_u1889_o;
  wire _al_u1891_o;
  wire _al_u1893_o;
  wire _al_u1895_o;
  wire _al_u1897_o;
  wire _al_u1899_o;
  wire _al_u1901_o;
  wire _al_u1903_o;
  wire _al_u1905_o;
  wire _al_u1906_o;
  wire _al_u1907_o;
  wire _al_u1908_o;
  wire _al_u1909_o;
  wire _al_u1910_o;
  wire _al_u1911_o;
  wire _al_u1912_o;
  wire _al_u1913_o;
  wire _al_u1914_o;
  wire _al_u1915_o;
  wire _al_u1916_o;
  wire _al_u1917_o;
  wire _al_u1918_o;
  wire _al_u1919_o;
  wire _al_u1920_o;
  wire _al_u1921_o;
  wire _al_u1922_o;
  wire _al_u1923_o;
  wire _al_u1924_o;
  wire _al_u1925_o;
  wire _al_u1926_o;
  wire _al_u1927_o;
  wire _al_u1930_o;
  wire _al_u1931_o;
  wire _al_u1932_o;
  wire _al_u1933_o;
  wire _al_u1934_o;
  wire _al_u1935_o;
  wire _al_u1937_o;
  wire _al_u1939_o;
  wire _al_u1941_o;
  wire _al_u1943_o;
  wire _al_u1945_o;
  wire _al_u1947_o;
  wire _al_u1949_o;
  wire _al_u1951_o;
  wire _al_u1953_o;
  wire _al_u1955_o;
  wire _al_u1957_o;
  wire _al_u1959_o;
  wire _al_u1961_o;
  wire _al_u1963_o;
  wire _al_u1965_o;
  wire _al_u1967_o;
  wire _al_u1969_o;
  wire _al_u1971_o;
  wire _al_u1973_o;
  wire _al_u1975_o;
  wire _al_u1977_o;
  wire _al_u1979_o;
  wire _al_u1981_o;
  wire _al_u1983_o;
  wire _al_u1985_o;
  wire _al_u1986_o;
  wire _al_u1987_o;
  wire _al_u1988_o;
  wire _al_u1989_o;
  wire _al_u1990_o;
  wire _al_u1991_o;
  wire _al_u1992_o;
  wire _al_u1993_o;
  wire _al_u1994_o;
  wire _al_u1995_o;
  wire _al_u1996_o;
  wire _al_u1997_o;
  wire _al_u1998_o;
  wire _al_u1999_o;
  wire _al_u2000_o;
  wire _al_u2001_o;
  wire _al_u2002_o;
  wire _al_u2003_o;
  wire _al_u2004_o;
  wire _al_u2005_o;
  wire _al_u2006_o;
  wire _al_u2007_o;
  wire _al_u2008_o;
  wire _al_u2009_o;
  wire _al_u2012_o;
  wire _al_u2013_o;
  wire _al_u2014_o;
  wire _al_u2015_o;
  wire _al_u2016_o;
  wire _al_u2017_o;
  wire _al_u2019_o;
  wire _al_u2021_o;
  wire _al_u2023_o;
  wire _al_u2025_o;
  wire _al_u2027_o;
  wire _al_u2029_o;
  wire _al_u2031_o;
  wire _al_u2033_o;
  wire _al_u2035_o;
  wire _al_u2037_o;
  wire _al_u2039_o;
  wire _al_u2041_o;
  wire _al_u2043_o;
  wire _al_u2045_o;
  wire _al_u2047_o;
  wire _al_u2049_o;
  wire _al_u2051_o;
  wire _al_u2053_o;
  wire _al_u2055_o;
  wire _al_u2057_o;
  wire _al_u2059_o;
  wire _al_u2061_o;
  wire _al_u2063_o;
  wire _al_u2065_o;
  wire _al_u2067_o;
  wire _al_u2068_o;
  wire _al_u2069_o;
  wire _al_u2070_o;
  wire _al_u2071_o;
  wire _al_u2072_o;
  wire _al_u2073_o;
  wire _al_u2074_o;
  wire _al_u2075_o;
  wire _al_u2076_o;
  wire _al_u2077_o;
  wire _al_u2078_o;
  wire _al_u2079_o;
  wire _al_u2080_o;
  wire _al_u2081_o;
  wire _al_u2082_o;
  wire _al_u2083_o;
  wire _al_u2084_o;
  wire _al_u2085_o;
  wire _al_u2086_o;
  wire _al_u2087_o;
  wire _al_u2088_o;
  wire _al_u2089_o;
  wire _al_u2090_o;
  wire _al_u2091_o;
  wire _al_u2094_o;
  wire _al_u2095_o;
  wire _al_u2096_o;
  wire _al_u2097_o;
  wire _al_u2098_o;
  wire _al_u2099_o;
  wire _al_u2101_o;
  wire _al_u2103_o;
  wire _al_u2105_o;
  wire _al_u2107_o;
  wire _al_u2109_o;
  wire _al_u2111_o;
  wire _al_u2113_o;
  wire _al_u2115_o;
  wire _al_u2117_o;
  wire _al_u2119_o;
  wire _al_u2121_o;
  wire _al_u2123_o;
  wire _al_u2125_o;
  wire _al_u2127_o;
  wire _al_u2129_o;
  wire _al_u2131_o;
  wire _al_u2133_o;
  wire _al_u2135_o;
  wire _al_u2137_o;
  wire _al_u2139_o;
  wire _al_u2141_o;
  wire _al_u2143_o;
  wire _al_u2145_o;
  wire _al_u2147_o;
  wire _al_u2149_o;
  wire _al_u2150_o;
  wire _al_u2151_o;
  wire _al_u2152_o;
  wire _al_u2153_o;
  wire _al_u2154_o;
  wire _al_u2155_o;
  wire _al_u2156_o;
  wire _al_u2157_o;
  wire _al_u2158_o;
  wire _al_u2159_o;
  wire _al_u2160_o;
  wire _al_u2161_o;
  wire _al_u2162_o;
  wire _al_u2163_o;
  wire _al_u2164_o;
  wire _al_u2165_o;
  wire _al_u2166_o;
  wire _al_u2167_o;
  wire _al_u2168_o;
  wire _al_u2169_o;
  wire _al_u2170_o;
  wire _al_u2171_o;
  wire _al_u2172_o;
  wire _al_u2173_o;
  wire _al_u2176_o;
  wire _al_u2177_o;
  wire _al_u2178_o;
  wire _al_u2179_o;
  wire _al_u2180_o;
  wire _al_u2181_o;
  wire _al_u2183_o;
  wire _al_u2185_o;
  wire _al_u2187_o;
  wire _al_u2189_o;
  wire _al_u2191_o;
  wire _al_u2193_o;
  wire _al_u2195_o;
  wire _al_u2197_o;
  wire _al_u2199_o;
  wire _al_u2201_o;
  wire _al_u2203_o;
  wire _al_u2205_o;
  wire _al_u2207_o;
  wire _al_u2209_o;
  wire _al_u2211_o;
  wire _al_u2213_o;
  wire _al_u2215_o;
  wire _al_u2217_o;
  wire _al_u2219_o;
  wire _al_u2221_o;
  wire _al_u2223_o;
  wire _al_u2225_o;
  wire _al_u2227_o;
  wire _al_u2229_o;
  wire _al_u2231_o;
  wire _al_u2232_o;
  wire _al_u2233_o;
  wire _al_u2234_o;
  wire _al_u2235_o;
  wire _al_u2236_o;
  wire _al_u2237_o;
  wire _al_u2238_o;
  wire _al_u2239_o;
  wire _al_u2240_o;
  wire _al_u2241_o;
  wire _al_u2242_o;
  wire _al_u2243_o;
  wire _al_u2244_o;
  wire _al_u2245_o;
  wire _al_u2246_o;
  wire _al_u2247_o;
  wire _al_u2248_o;
  wire _al_u2249_o;
  wire _al_u2250_o;
  wire _al_u2251_o;
  wire _al_u2252_o;
  wire _al_u2253_o;
  wire _al_u2256_o;
  wire _al_u2257_o;
  wire _al_u2258_o;
  wire _al_u2259_o;
  wire _al_u2260_o;
  wire _al_u2261_o;
  wire _al_u2263_o;
  wire _al_u2265_o;
  wire _al_u2267_o;
  wire _al_u2269_o;
  wire _al_u2271_o;
  wire _al_u2273_o;
  wire _al_u2275_o;
  wire _al_u2277_o;
  wire _al_u2279_o;
  wire _al_u2281_o;
  wire _al_u2283_o;
  wire _al_u2285_o;
  wire _al_u2287_o;
  wire _al_u2289_o;
  wire _al_u2291_o;
  wire _al_u2293_o;
  wire _al_u2295_o;
  wire _al_u2297_o;
  wire _al_u2299_o;
  wire _al_u2301_o;
  wire _al_u2303_o;
  wire _al_u2305_o;
  wire _al_u2307_o;
  wire _al_u2309_o;
  wire _al_u2311_o;
  wire _al_u2312_o;
  wire _al_u2313_o;
  wire _al_u2314_o;
  wire _al_u2315_o;
  wire _al_u2316_o;
  wire _al_u2317_o;
  wire _al_u2318_o;
  wire _al_u2319_o;
  wire _al_u2320_o;
  wire _al_u2321_o;
  wire _al_u2322_o;
  wire _al_u2323_o;
  wire _al_u2324_o;
  wire _al_u2325_o;
  wire _al_u2326_o;
  wire _al_u2327_o;
  wire _al_u2328_o;
  wire _al_u2329_o;
  wire _al_u2330_o;
  wire _al_u2331_o;
  wire _al_u2332_o;
  wire _al_u2333_o;
  wire _al_u2334_o;
  wire _al_u2335_o;
  wire _al_u2338_o;
  wire _al_u2339_o;
  wire _al_u2340_o;
  wire _al_u2341_o;
  wire _al_u2342_o;
  wire _al_u2343_o;
  wire _al_u2345_o;
  wire _al_u2347_o;
  wire _al_u2349_o;
  wire _al_u2351_o;
  wire _al_u2353_o;
  wire _al_u2355_o;
  wire _al_u2357_o;
  wire _al_u2359_o;
  wire _al_u2361_o;
  wire _al_u2363_o;
  wire _al_u2365_o;
  wire _al_u2367_o;
  wire _al_u2369_o;
  wire _al_u2371_o;
  wire _al_u2373_o;
  wire _al_u2375_o;
  wire _al_u2377_o;
  wire _al_u2379_o;
  wire _al_u2381_o;
  wire _al_u2383_o;
  wire _al_u2385_o;
  wire _al_u2387_o;
  wire _al_u2389_o;
  wire _al_u2391_o;
  wire _al_u2393_o;
  wire _al_u2394_o;
  wire _al_u2395_o;
  wire _al_u2396_o;
  wire _al_u2397_o;
  wire _al_u2398_o;
  wire _al_u2399_o;
  wire _al_u2400_o;
  wire _al_u2401_o;
  wire _al_u2402_o;
  wire _al_u2403_o;
  wire _al_u2404_o;
  wire _al_u2405_o;
  wire _al_u2406_o;
  wire _al_u2407_o;
  wire _al_u2408_o;
  wire _al_u2409_o;
  wire _al_u2410_o;
  wire _al_u2411_o;
  wire _al_u2412_o;
  wire _al_u2413_o;
  wire _al_u2414_o;
  wire _al_u2415_o;
  wire _al_u2418_o;
  wire _al_u2419_o;
  wire _al_u2420_o;
  wire _al_u2421_o;
  wire _al_u2422_o;
  wire _al_u2423_o;
  wire _al_u2425_o;
  wire _al_u2427_o;
  wire _al_u2429_o;
  wire _al_u2431_o;
  wire _al_u2433_o;
  wire _al_u2435_o;
  wire _al_u2437_o;
  wire _al_u2439_o;
  wire _al_u2441_o;
  wire _al_u2443_o;
  wire _al_u2445_o;
  wire _al_u2447_o;
  wire _al_u2449_o;
  wire _al_u2451_o;
  wire _al_u2453_o;
  wire _al_u2455_o;
  wire _al_u2457_o;
  wire _al_u2459_o;
  wire _al_u2461_o;
  wire _al_u2463_o;
  wire _al_u2465_o;
  wire _al_u2467_o;
  wire _al_u2469_o;
  wire _al_u2471_o;
  wire _al_u2473_o;
  wire _al_u2474_o;
  wire _al_u2475_o;
  wire _al_u2476_o;
  wire _al_u2477_o;
  wire _al_u2478_o;
  wire _al_u2479_o;
  wire _al_u2480_o;
  wire _al_u2481_o;
  wire _al_u2482_o;
  wire _al_u2483_o;
  wire _al_u2484_o;
  wire _al_u2485_o;
  wire _al_u2486_o;
  wire _al_u2487_o;
  wire _al_u2488_o;
  wire _al_u2489_o;
  wire _al_u2490_o;
  wire _al_u2491_o;
  wire _al_u2492_o;
  wire _al_u2493_o;
  wire _al_u2494_o;
  wire _al_u2495_o;
  wire _al_u2496_o;
  wire _al_u2497_o;
  wire _al_u2500_o;
  wire _al_u2501_o;
  wire _al_u2502_o;
  wire _al_u2503_o;
  wire _al_u2504_o;
  wire _al_u2505_o;
  wire _al_u2507_o;
  wire _al_u2509_o;
  wire _al_u2511_o;
  wire _al_u2513_o;
  wire _al_u2515_o;
  wire _al_u2517_o;
  wire _al_u2519_o;
  wire _al_u2521_o;
  wire _al_u2523_o;
  wire _al_u2525_o;
  wire _al_u2527_o;
  wire _al_u2529_o;
  wire _al_u2531_o;
  wire _al_u2533_o;
  wire _al_u2535_o;
  wire _al_u2537_o;
  wire _al_u2539_o;
  wire _al_u2541_o;
  wire _al_u2543_o;
  wire _al_u2545_o;
  wire _al_u2547_o;
  wire _al_u2549_o;
  wire _al_u2551_o;
  wire _al_u2553_o;
  wire _al_u2555_o;
  wire _al_u2556_o;
  wire _al_u2557_o;
  wire _al_u2558_o;
  wire _al_u2559_o;
  wire _al_u2560_o;
  wire _al_u2561_o;
  wire _al_u2562_o;
  wire _al_u2563_o;
  wire _al_u2564_o;
  wire _al_u2565_o;
  wire _al_u2566_o;
  wire _al_u2567_o;
  wire _al_u2568_o;
  wire _al_u2569_o;
  wire _al_u2570_o;
  wire _al_u2571_o;
  wire _al_u2572_o;
  wire _al_u2573_o;
  wire _al_u2574_o;
  wire _al_u2575_o;
  wire _al_u2576_o;
  wire _al_u2579_o;
  wire _al_u2580_o;
  wire _al_u2581_o;
  wire _al_u2582_o;
  wire _al_u2583_o;
  wire _al_u2584_o;
  wire _al_u2586_o;
  wire _al_u2588_o;
  wire _al_u2590_o;
  wire _al_u2592_o;
  wire _al_u2594_o;
  wire _al_u2596_o;
  wire _al_u2598_o;
  wire _al_u2600_o;
  wire _al_u2602_o;
  wire _al_u2604_o;
  wire _al_u2606_o;
  wire _al_u2608_o;
  wire _al_u2610_o;
  wire _al_u2612_o;
  wire _al_u2614_o;
  wire _al_u2616_o;
  wire _al_u2618_o;
  wire _al_u2620_o;
  wire _al_u2622_o;
  wire _al_u2624_o;
  wire _al_u2626_o;
  wire _al_u2628_o;
  wire _al_u2630_o;
  wire _al_u2632_o;
  wire _al_u2634_o;
  wire _al_u2635_o;
  wire _al_u2636_o;
  wire _al_u2637_o;
  wire _al_u2638_o;
  wire _al_u2639_o;
  wire _al_u2640_o;
  wire _al_u2641_o;
  wire _al_u2642_o;
  wire _al_u2643_o;
  wire _al_u2644_o;
  wire _al_u2645_o;
  wire _al_u2646_o;
  wire _al_u2647_o;
  wire _al_u2648_o;
  wire _al_u2649_o;
  wire _al_u2650_o;
  wire _al_u2651_o;
  wire _al_u2652_o;
  wire _al_u2653_o;
  wire _al_u2654_o;
  wire _al_u2655_o;
  wire _al_u2656_o;
  wire _al_u2657_o;
  wire _al_u2658_o;
  wire _al_u2661_o;
  wire _al_u2662_o;
  wire _al_u2663_o;
  wire _al_u2664_o;
  wire _al_u2665_o;
  wire _al_u2666_o;
  wire _al_u2668_o;
  wire _al_u2670_o;
  wire _al_u2672_o;
  wire _al_u2674_o;
  wire _al_u2676_o;
  wire _al_u2678_o;
  wire _al_u2680_o;
  wire _al_u2682_o;
  wire _al_u2684_o;
  wire _al_u2686_o;
  wire _al_u2688_o;
  wire _al_u2690_o;
  wire _al_u2692_o;
  wire _al_u2694_o;
  wire _al_u2696_o;
  wire _al_u2698_o;
  wire _al_u2700_o;
  wire _al_u2702_o;
  wire _al_u2704_o;
  wire _al_u2706_o;
  wire _al_u2708_o;
  wire _al_u2710_o;
  wire _al_u2712_o;
  wire _al_u2714_o;
  wire _al_u2716_o;
  wire _al_u2717_o;
  wire _al_u2718_o;
  wire _al_u2719_o;
  wire _al_u2720_o;
  wire _al_u2721_o;
  wire _al_u2722_o;
  wire _al_u2723_o;
  wire _al_u2724_o;
  wire _al_u2725_o;
  wire _al_u2726_o;
  wire _al_u2727_o;
  wire _al_u2728_o;
  wire _al_u2729_o;
  wire _al_u2730_o;
  wire _al_u2731_o;
  wire _al_u2732_o;
  wire _al_u2733_o;
  wire _al_u2734_o;
  wire _al_u2735_o;
  wire _al_u2736_o;
  wire _al_u2737_o;
  wire _al_u2740_o;
  wire _al_u2741_o;
  wire _al_u2742_o;
  wire _al_u2743_o;
  wire _al_u2744_o;
  wire _al_u2745_o;
  wire _al_u2747_o;
  wire _al_u2749_o;
  wire _al_u2751_o;
  wire _al_u2753_o;
  wire _al_u2755_o;
  wire _al_u2757_o;
  wire _al_u2759_o;
  wire _al_u2761_o;
  wire _al_u2763_o;
  wire _al_u2765_o;
  wire _al_u2767_o;
  wire _al_u2769_o;
  wire _al_u2771_o;
  wire _al_u2773_o;
  wire _al_u2775_o;
  wire _al_u2777_o;
  wire _al_u2779_o;
  wire _al_u2781_o;
  wire _al_u2783_o;
  wire _al_u2785_o;
  wire _al_u2787_o;
  wire _al_u2789_o;
  wire _al_u2791_o;
  wire _al_u2793_o;
  wire _al_u2795_o;
  wire _al_u2796_o;
  wire _al_u2797_o;
  wire _al_u2798_o;
  wire _al_u2799_o;
  wire _al_u2800_o;
  wire _al_u2801_o;
  wire _al_u2802_o;
  wire _al_u2803_o;
  wire _al_u2804_o;
  wire _al_u2805_o;
  wire _al_u2806_o;
  wire _al_u2807_o;
  wire _al_u2808_o;
  wire _al_u2809_o;
  wire _al_u2810_o;
  wire _al_u2811_o;
  wire _al_u2812_o;
  wire _al_u2813_o;
  wire _al_u2814_o;
  wire _al_u2815_o;
  wire _al_u2816_o;
  wire _al_u2817_o;
  wire _al_u2820_o;
  wire _al_u2821_o;
  wire _al_u2822_o;
  wire _al_u2823_o;
  wire _al_u2824_o;
  wire _al_u2825_o;
  wire _al_u2827_o;
  wire _al_u2829_o;
  wire _al_u2831_o;
  wire _al_u2833_o;
  wire _al_u2835_o;
  wire _al_u2837_o;
  wire _al_u2839_o;
  wire _al_u2841_o;
  wire _al_u2843_o;
  wire _al_u2845_o;
  wire _al_u2847_o;
  wire _al_u2849_o;
  wire _al_u2851_o;
  wire _al_u2853_o;
  wire _al_u2855_o;
  wire _al_u2857_o;
  wire _al_u2859_o;
  wire _al_u2861_o;
  wire _al_u2863_o;
  wire _al_u2865_o;
  wire _al_u2867_o;
  wire _al_u2869_o;
  wire _al_u2871_o;
  wire _al_u2873_o;
  wire _al_u2875_o;
  wire _al_u2876_o;
  wire _al_u2877_o;
  wire _al_u2878_o;
  wire _al_u2879_o;
  wire _al_u2880_o;
  wire _al_u2881_o;
  wire _al_u2882_o;
  wire _al_u2883_o;
  wire _al_u2884_o;
  wire _al_u2885_o;
  wire _al_u2886_o;
  wire _al_u2887_o;
  wire _al_u2888_o;
  wire _al_u2889_o;
  wire _al_u2890_o;
  wire _al_u2891_o;
  wire _al_u2892_o;
  wire _al_u2893_o;
  wire _al_u2894_o;
  wire _al_u2895_o;
  wire _al_u2896_o;
  wire _al_u2899_o;
  wire _al_u2900_o;
  wire _al_u2901_o;
  wire _al_u2902_o;
  wire _al_u2903_o;
  wire _al_u2904_o;
  wire _al_u2906_o;
  wire _al_u2908_o;
  wire _al_u2910_o;
  wire _al_u2912_o;
  wire _al_u2914_o;
  wire _al_u2916_o;
  wire _al_u2918_o;
  wire _al_u2920_o;
  wire _al_u2922_o;
  wire _al_u2924_o;
  wire _al_u2926_o;
  wire _al_u2928_o;
  wire _al_u2930_o;
  wire _al_u2932_o;
  wire _al_u2934_o;
  wire _al_u2936_o;
  wire _al_u2938_o;
  wire _al_u2940_o;
  wire _al_u2942_o;
  wire _al_u2944_o;
  wire _al_u2946_o;
  wire _al_u2948_o;
  wire _al_u2950_o;
  wire _al_u2952_o;
  wire _al_u2954_o;
  wire _al_u2955_o;
  wire _al_u2956_o;
  wire _al_u2957_o;
  wire _al_u2958_o;
  wire _al_u2959_o;
  wire _al_u2960_o;
  wire _al_u2961_o;
  wire _al_u2962_o;
  wire _al_u2963_o;
  wire _al_u2964_o;
  wire _al_u2965_o;
  wire _al_u2966_o;
  wire _al_u2967_o;
  wire _al_u2968_o;
  wire _al_u2969_o;
  wire _al_u2970_o;
  wire _al_u2971_o;
  wire _al_u2972_o;
  wire _al_u2973_o;
  wire _al_u2974_o;
  wire _al_u2975_o;
  wire _al_u2976_o;
  wire _al_u2977_o;
  wire _al_u2978_o;
  wire _al_u2980_o;
  wire _al_u2981_o;
  wire _al_u2982_o;
  wire _al_u2983_o;
  wire _al_u2984_o;
  wire _al_u2985_o;
  wire _al_u2986_o;
  wire _al_u2987_o;
  wire _al_u2988_o;
  wire _al_u3007_o;
  wire _al_u3008_o;
  wire _al_u3010_o;
  wire _al_u3011_o;
  wire _al_u3013_o;
  wire _al_u3014_o;
  wire _al_u3016_o;
  wire _al_u3017_o;
  wire _al_u3019_o;
  wire _al_u3020_o;
  wire _al_u3022_o;
  wire _al_u3023_o;
  wire _al_u3025_o;
  wire _al_u3026_o;
  wire _al_u3028_o;
  wire _al_u3029_o;
  wire _al_u3031_o;
  wire _al_u3032_o;
  wire _al_u3034_o;
  wire _al_u3035_o;
  wire _al_u3037_o;
  wire _al_u3038_o;
  wire _al_u3040_o;
  wire _al_u3041_o;
  wire _al_u3043_o;
  wire _al_u3044_o;
  wire _al_u3046_o;
  wire _al_u3047_o;
  wire _al_u3049_o;
  wire _al_u3050_o;
  wire _al_u3052_o;
  wire _al_u3053_o;
  wire _al_u3055_o;
  wire _al_u3061_o;
  wire _al_u3062_o;
  wire _al_u3065_o;
  wire _al_u3068_o;
  wire _al_u3070_o;
  wire _al_u3072_o;
  wire _al_u3074_o;
  wire _al_u3076_o;
  wire _al_u3078_o;
  wire _al_u3080_o;
  wire _al_u3082_o;
  wire _al_u3085_o;
  wire _al_u3087_o;
  wire _al_u3089_o;
  wire _al_u3092_o;
  wire _al_u3094_o;
  wire _al_u3095_o;
  wire _al_u3096_o;
  wire _al_u3097_o;
  wire _al_u3098_o;
  wire _al_u3100_o;
  wire _al_u3101_o;
  wire _al_u3102_o;
  wire _al_u3103_o;
  wire _al_u3104_o;
  wire _al_u3105_o;
  wire _al_u3106_o;
  wire _al_u3107_o;
  wire _al_u3108_o;
  wire _al_u3109_o;
  wire _al_u3111_o;
  wire _al_u3112_o;
  wire _al_u3113_o;
  wire _al_u3114_o;
  wire _al_u3115_o;
  wire _al_u3116_o;
  wire _al_u3117_o;
  wire _al_u3118_o;
  wire _al_u3119_o;
  wire _al_u3120_o;
  wire _al_u3122_o;
  wire _al_u3123_o;
  wire _al_u3124_o;
  wire _al_u3125_o;
  wire _al_u3126_o;
  wire _al_u3127_o;
  wire _al_u3128_o;
  wire _al_u3129_o;
  wire _al_u3130_o;
  wire _al_u3131_o;
  wire _al_u3133_o;
  wire _al_u3134_o;
  wire _al_u3135_o;
  wire _al_u3136_o;
  wire _al_u3137_o;
  wire _al_u3138_o;
  wire _al_u3139_o;
  wire _al_u3140_o;
  wire _al_u3141_o;
  wire _al_u3142_o;
  wire _al_u3143_o;
  wire _al_u3145_o;
  wire _al_u3146_o;
  wire _al_u3147_o;
  wire _al_u3148_o;
  wire _al_u3149_o;
  wire _al_u3150_o;
  wire _al_u3151_o;
  wire _al_u3152_o;
  wire _al_u3153_o;
  wire _al_u3154_o;
  wire _al_u3156_o;
  wire _al_u3157_o;
  wire _al_u3158_o;
  wire _al_u3159_o;
  wire _al_u3160_o;
  wire _al_u3161_o;
  wire _al_u3162_o;
  wire _al_u3163_o;
  wire _al_u3164_o;
  wire _al_u3165_o;
  wire _al_u3167_o;
  wire _al_u3168_o;
  wire _al_u3169_o;
  wire _al_u3170_o;
  wire _al_u3171_o;
  wire _al_u3172_o;
  wire _al_u3173_o;
  wire _al_u3174_o;
  wire _al_u3175_o;
  wire _al_u3176_o;
  wire _al_u3178_o;
  wire _al_u3179_o;
  wire _al_u3180_o;
  wire _al_u3181_o;
  wire _al_u3182_o;
  wire _al_u3183_o;
  wire _al_u3184_o;
  wire _al_u3185_o;
  wire _al_u3186_o;
  wire _al_u3187_o;
  wire _al_u3189_o;
  wire _al_u3190_o;
  wire _al_u3191_o;
  wire _al_u3192_o;
  wire _al_u3193_o;
  wire _al_u3194_o;
  wire _al_u3195_o;
  wire _al_u3196_o;
  wire _al_u3197_o;
  wire _al_u3198_o;
  wire _al_u3200_o;
  wire _al_u3201_o;
  wire _al_u3202_o;
  wire _al_u3203_o;
  wire _al_u3204_o;
  wire _al_u3205_o;
  wire _al_u3206_o;
  wire _al_u3207_o;
  wire _al_u3208_o;
  wire _al_u3209_o;
  wire _al_u3211_o;
  wire _al_u3212_o;
  wire _al_u3213_o;
  wire _al_u3214_o;
  wire _al_u3215_o;
  wire _al_u3216_o;
  wire _al_u3217_o;
  wire _al_u3218_o;
  wire _al_u3219_o;
  wire _al_u3220_o;
  wire _al_u3222_o;
  wire _al_u3223_o;
  wire _al_u3224_o;
  wire _al_u3225_o;
  wire _al_u3226_o;
  wire _al_u3227_o;
  wire _al_u3228_o;
  wire _al_u3229_o;
  wire _al_u3230_o;
  wire _al_u3231_o;
  wire _al_u3233_o;
  wire _al_u3234_o;
  wire _al_u3235_o;
  wire _al_u3236_o;
  wire _al_u3237_o;
  wire _al_u3238_o;
  wire _al_u3239_o;
  wire _al_u3240_o;
  wire _al_u3241_o;
  wire _al_u3242_o;
  wire _al_u3244_o;
  wire _al_u3245_o;
  wire _al_u3246_o;
  wire _al_u3247_o;
  wire _al_u3248_o;
  wire _al_u3249_o;
  wire _al_u3250_o;
  wire _al_u3251_o;
  wire _al_u3252_o;
  wire _al_u3253_o;
  wire _al_u3255_o;
  wire _al_u3256_o;
  wire _al_u3257_o;
  wire _al_u3258_o;
  wire _al_u3259_o;
  wire _al_u3260_o;
  wire _al_u3261_o;
  wire _al_u3262_o;
  wire _al_u3263_o;
  wire _al_u3264_o;
  wire _al_u3266_o;
  wire _al_u3267_o;
  wire _al_u3268_o;
  wire _al_u3269_o;
  wire _al_u3270_o;
  wire _al_u3271_o;
  wire _al_u3272_o;
  wire _al_u3273_o;
  wire _al_u3274_o;
  wire _al_u3275_o;
  wire _al_u3277_o;
  wire _al_u3278_o;
  wire _al_u3279_o;
  wire _al_u3280_o;
  wire _al_u3281_o;
  wire _al_u3282_o;
  wire _al_u3283_o;
  wire _al_u3284_o;
  wire _al_u3285_o;
  wire _al_u3286_o;
  wire _al_u3288_o;
  wire _al_u3289_o;
  wire _al_u3290_o;
  wire _al_u3291_o;
  wire _al_u3292_o;
  wire _al_u3293_o;
  wire _al_u3294_o;
  wire _al_u3295_o;
  wire _al_u3296_o;
  wire _al_u3297_o;
  wire _al_u3299_o;
  wire _al_u3300_o;
  wire _al_u3301_o;
  wire _al_u3302_o;
  wire _al_u3303_o;
  wire _al_u3304_o;
  wire _al_u3305_o;
  wire _al_u3306_o;
  wire _al_u3307_o;
  wire _al_u3308_o;
  wire _al_u3310_o;
  wire _al_u3311_o;
  wire _al_u3312_o;
  wire _al_u3313_o;
  wire _al_u3314_o;
  wire _al_u3315_o;
  wire _al_u3316_o;
  wire _al_u3317_o;
  wire _al_u3318_o;
  wire _al_u3319_o;
  wire _al_u3321_o;
  wire _al_u3322_o;
  wire _al_u3323_o;
  wire _al_u3324_o;
  wire _al_u3325_o;
  wire _al_u3326_o;
  wire _al_u3327_o;
  wire _al_u3328_o;
  wire _al_u3329_o;
  wire _al_u3330_o;
  wire _al_u3332_o;
  wire _al_u3333_o;
  wire _al_u3334_o;
  wire _al_u3335_o;
  wire _al_u3336_o;
  wire _al_u3337_o;
  wire _al_u3338_o;
  wire _al_u3339_o;
  wire _al_u3340_o;
  wire _al_u3341_o;
  wire _al_u3343_o;
  wire _al_u3344_o;
  wire _al_u3345_o;
  wire _al_u3346_o;
  wire _al_u3347_o;
  wire _al_u3348_o;
  wire _al_u3349_o;
  wire _al_u3350_o;
  wire _al_u3351_o;
  wire _al_u3352_o;
  wire _al_u734_o;
  wire _al_u735_o;
  wire _al_u736_o;
  wire _al_u737_o;
  wire _al_u738_o;
  wire _al_u739_o;
  wire _al_u740_o;
  wire _al_u771_o;
  wire _al_u772_o;
  wire _al_u773_o;
  wire _al_u774_o;
  wire _al_u775_o;
  wire _al_u776_o;
  wire _al_u777_o;
  wire _al_u808_o;
  wire _al_u809_o;
  wire _al_u810_o;
  wire _al_u811_o;
  wire _al_u812_o;
  wire _al_u813_o;
  wire _al_u814_o;
  wire _al_u845_o;
  wire _al_u846_o;
  wire _al_u847_o;
  wire _al_u848_o;
  wire _al_u849_o;
  wire _al_u850_o;
  wire _al_u851_o;
  wire _al_u882_o;
  wire _al_u883_o;
  wire _al_u884_o;
  wire _al_u885_o;
  wire _al_u886_o;
  wire _al_u887_o;
  wire _al_u888_o;
  wire _al_u919_o;
  wire _al_u920_o;
  wire _al_u921_o;
  wire _al_u922_o;
  wire _al_u923_o;
  wire _al_u924_o;
  wire _al_u925_o;
  wire _al_u956_o;
  wire _al_u957_o;
  wire _al_u958_o;
  wire _al_u959_o;
  wire _al_u960_o;
  wire _al_u961_o;
  wire _al_u962_o;
  wire _al_u993_o;
  wire _al_u994_o;
  wire _al_u995_o;
  wire _al_u996_o;
  wire _al_u997_o;
  wire _al_u998_o;
  wire _al_u999_o;
  wire \add0/c11 ;
  wire \add0/c15 ;
  wire \add0/c19 ;
  wire \add0/c23 ;
  wire \add0/c27 ;
  wire \add0/c3 ;
  wire \add0/c31 ;
  wire \add0/c7 ;
  wire clk100m;  // CPLD_SOC_AHB_TOP.v(13)
  wire clk100m_keep;
  wire clk25m;  // CPLD_SOC_AHB_TOP.v(13)
  wire clkin_pad;  // CPLD_SOC_AHB_TOP.v(3)
  wire n4_neg;
  wire rst_n_pad;  // CPLD_SOC_AHB_TOP.v(4)
  wire rstn;  // CPLD_SOC_AHB_TOP.v(13)

  // src/OnePWM.v(26)
  // src/OnePWM.v(26)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*~(~D*B*~A))"),
    //.LUTF1("(C*~(~D*B*~A))"),
    //.LUTG0("(C*~(~D*B*~A))"),
    //.LUTG1("(C*~(~D*B*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000010110000),
    .INIT_LUTF1(16'b1111000010110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \PWM0/State_reg|PWMF/State_reg  (
    .a({_al_u3007_o,_al_u3052_o}),
    .b({\PWM0/n0_lutinv ,\PWMF/n0_lutinv }),
    .c({_al_u3008_o,_al_u3053_o}),
    .clk(clk100m),
    .d({pwm_start_stop[16],pwm_start_stop[31]}),
    .sr(rstn),
    .q({pwm_state_read[0],pwm_state_read[15]}));  // src/OnePWM.v(26)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[0]  (
    .i(\PWM0/RemaTxNum[0]_keep ),
    .o(pnumcnt0[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[10]  (
    .i(\PWM0/RemaTxNum[10]_keep ),
    .o(pnumcnt0[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[11]  (
    .i(\PWM0/RemaTxNum[11]_keep ),
    .o(pnumcnt0[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[12]  (
    .i(\PWM0/RemaTxNum[12]_keep ),
    .o(pnumcnt0[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[13]  (
    .i(\PWM0/RemaTxNum[13]_keep ),
    .o(pnumcnt0[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[14]  (
    .i(\PWM0/RemaTxNum[14]_keep ),
    .o(pnumcnt0[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[15]  (
    .i(\PWM0/RemaTxNum[15]_keep ),
    .o(pnumcnt0[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[16]  (
    .i(\PWM0/RemaTxNum[16]_keep ),
    .o(pnumcnt0[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[17]  (
    .i(\PWM0/RemaTxNum[17]_keep ),
    .o(pnumcnt0[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[18]  (
    .i(\PWM0/RemaTxNum[18]_keep ),
    .o(pnumcnt0[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[19]  (
    .i(\PWM0/RemaTxNum[19]_keep ),
    .o(pnumcnt0[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[1]  (
    .i(\PWM0/RemaTxNum[1]_keep ),
    .o(pnumcnt0[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[20]  (
    .i(\PWM0/RemaTxNum[20]_keep ),
    .o(pnumcnt0[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[21]  (
    .i(\PWM0/RemaTxNum[21]_keep ),
    .o(pnumcnt0[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[22]  (
    .i(\PWM0/RemaTxNum[22]_keep ),
    .o(pnumcnt0[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[23]  (
    .i(\PWM0/RemaTxNum[23]_keep ),
    .o(pnumcnt0[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[2]  (
    .i(\PWM0/RemaTxNum[2]_keep ),
    .o(pnumcnt0[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[3]  (
    .i(\PWM0/RemaTxNum[3]_keep ),
    .o(pnumcnt0[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[4]  (
    .i(\PWM0/RemaTxNum[4]_keep ),
    .o(pnumcnt0[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[5]  (
    .i(\PWM0/RemaTxNum[5]_keep ),
    .o(pnumcnt0[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[6]  (
    .i(\PWM0/RemaTxNum[6]_keep ),
    .o(pnumcnt0[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[7]  (
    .i(\PWM0/RemaTxNum[7]_keep ),
    .o(pnumcnt0[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[8]  (
    .i(\PWM0/RemaTxNum[8]_keep ),
    .o(pnumcnt0[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[9]  (
    .i(\PWM0/RemaTxNum[9]_keep ),
    .o(pnumcnt0[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_dir  (
    .i(\PWM0/dir_keep ),
    .o(dir_pad[0]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[0]  (
    .i(\PWM0/pnumr[0]_keep ),
    .o(\PWM0/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[10]  (
    .i(\PWM0/pnumr[10]_keep ),
    .o(\PWM0/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[11]  (
    .i(\PWM0/pnumr[11]_keep ),
    .o(\PWM0/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[12]  (
    .i(\PWM0/pnumr[12]_keep ),
    .o(\PWM0/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[13]  (
    .i(\PWM0/pnumr[13]_keep ),
    .o(\PWM0/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[14]  (
    .i(\PWM0/pnumr[14]_keep ),
    .o(\PWM0/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[15]  (
    .i(\PWM0/pnumr[15]_keep ),
    .o(\PWM0/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[16]  (
    .i(\PWM0/pnumr[16]_keep ),
    .o(\PWM0/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[17]  (
    .i(\PWM0/pnumr[17]_keep ),
    .o(\PWM0/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[18]  (
    .i(\PWM0/pnumr[18]_keep ),
    .o(\PWM0/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[19]  (
    .i(\PWM0/pnumr[19]_keep ),
    .o(\PWM0/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[1]  (
    .i(\PWM0/pnumr[1]_keep ),
    .o(\PWM0/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[20]  (
    .i(\PWM0/pnumr[20]_keep ),
    .o(\PWM0/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[21]  (
    .i(\PWM0/pnumr[21]_keep ),
    .o(\PWM0/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[22]  (
    .i(\PWM0/pnumr[22]_keep ),
    .o(\PWM0/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[23]  (
    .i(\PWM0/pnumr[23]_keep ),
    .o(\PWM0/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[24]  (
    .i(\PWM0/pnumr[24]_keep ),
    .o(\PWM0/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[25]  (
    .i(\PWM0/pnumr[25]_keep ),
    .o(\PWM0/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[26]  (
    .i(\PWM0/pnumr[26]_keep ),
    .o(\PWM0/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[27]  (
    .i(\PWM0/pnumr[27]_keep ),
    .o(\PWM0/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[28]  (
    .i(\PWM0/pnumr[28]_keep ),
    .o(\PWM0/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[29]  (
    .i(\PWM0/pnumr[29]_keep ),
    .o(\PWM0/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[2]  (
    .i(\PWM0/pnumr[2]_keep ),
    .o(\PWM0/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[30]  (
    .i(\PWM0/pnumr[30]_keep ),
    .o(\PWM0/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[31]  (
    .i(\PWM0/pnumr[31]_keep ),
    .o(\PWM0/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[3]  (
    .i(\PWM0/pnumr[3]_keep ),
    .o(\PWM0/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[4]  (
    .i(\PWM0/pnumr[4]_keep ),
    .o(\PWM0/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[5]  (
    .i(\PWM0/pnumr[5]_keep ),
    .o(\PWM0/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[6]  (
    .i(\PWM0/pnumr[6]_keep ),
    .o(\PWM0/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[7]  (
    .i(\PWM0/pnumr[7]_keep ),
    .o(\PWM0/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[8]  (
    .i(\PWM0/pnumr[8]_keep ),
    .o(\PWM0/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[9]  (
    .i(\PWM0/pnumr[9]_keep ),
    .o(\PWM0/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pwm  (
    .i(\PWM0/pwm_keep ),
    .o(pwm_pad[0]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_stopreq  (
    .i(\PWM0/stopreq_keep ),
    .o(\PWM0/stopreq ));  // src/OnePWM.v(14)
  EF2_PHY_MSLICE #(
    //.LUT0("(D*~(C)*~((~0*~(B*A)))+D*C*~((~0*~(B*A)))+~(D)*C*(~0*~(B*A))+D*C*(~0*~(B*A)))"),
    //.LUT1("(D*~(C)*~((~1*~(B*A)))+D*C*~((~1*~(B*A)))+~(D)*C*(~1*~(B*A))+D*C*(~1*~(B*A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111100001110000),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/dir_reg  (
    .a({\PWM0/n24 ,\PWM0/n24 }),
    .b({\PWM0/n25_neg_lutinv ,\PWM0/n25_neg_lutinv }),
    .c({dir_pad[0],dir_pad[0]}),
    .clk(clk100m),
    .d({\PWM0/pnumr [31],\PWM0/pnumr [31]}),
    .mi({open_n33,pwm_start_stop[16]}),
    .q({open_n40,\PWM0/dir_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("~(~0*~(D*C*B*A))"),
    //.LUT1("~(~1*~(D*C*B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b1111111111111111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM0/pwm_reg  (
    .a({_al_u1365_o,_al_u1365_o}),
    .b({_al_u1372_o,_al_u1372_o}),
    .c({_al_u1374_o,_al_u1374_o}),
    .clk(clk100m),
    .d({_al_u1376_o,_al_u1376_o}),
    .mi({open_n52,pwm_pad[0]}),
    .sr(\PWM0/u14_sel_is_1_o ),
    .q({open_n58,\PWM0/pwm_keep }));  // src/OnePWM.v(45)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM0/reg0_b0|PWM0/reg0_b15  (
    .b({\PWM0/n12 [0],\PWM0/n12 [15]}),
    .c({freq0[0],freq0[15]}),
    .clk(clk100m),
    .d({\PWM0/n0_lutinv ,\PWM0/n0_lutinv }),
    .sr(\PWM0/n11 ),
    .q({\PWM0/FreCnt [0],\PWM0/FreCnt [15]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM0/reg0_b10|PWM0/reg0_b12  (
    .b({\PWM0/n12 [10],\PWM0/n12 [12]}),
    .c({freq0[10],freq0[12]}),
    .clk(clk100m),
    .d({\PWM0/n0_lutinv ,\PWM0/n0_lutinv }),
    .sr(\PWM0/n11 ),
    .q({\PWM0/FreCnt [10],\PWM0/FreCnt [12]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM0/reg0_b11|PWM0/reg0_b8  (
    .b({\PWM0/n12 [11],\PWM0/n12 [8]}),
    .c({freq0[11],freq0[8]}),
    .clk(clk100m),
    .d({\PWM0/n0_lutinv ,\PWM0/n0_lutinv }),
    .sr(\PWM0/n11 ),
    .q({\PWM0/FreCnt [11],\PWM0/FreCnt [8]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM0/reg0_b13|PWM0/reg0_b7  (
    .b({\PWM0/n12 [13],\PWM0/n12 [7]}),
    .c({freq0[13],freq0[7]}),
    .clk(clk100m),
    .d({\PWM0/n0_lutinv ,\PWM0/n0_lutinv }),
    .sr(\PWM0/n11 ),
    .q({\PWM0/FreCnt [13],\PWM0/FreCnt [7]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM0/reg0_b14|PWM0/reg0_b5  (
    .b({\PWM0/n12 [14],\PWM0/n12 [5]}),
    .c({freq0[14],freq0[5]}),
    .clk(clk100m),
    .d({\PWM0/n0_lutinv ,\PWM0/n0_lutinv }),
    .sr(\PWM0/n11 ),
    .q({\PWM0/FreCnt [14],\PWM0/FreCnt [5]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM0/reg0_b16|PWM0/reg0_b3  (
    .b({\PWM0/n12 [16],\PWM0/n12 [3]}),
    .c({freq0[16],freq0[3]}),
    .clk(clk100m),
    .d({\PWM0/n0_lutinv ,\PWM0/n0_lutinv }),
    .sr(\PWM0/n11 ),
    .q({\PWM0/FreCnt [16],\PWM0/FreCnt [3]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM0/reg0_b17|PWM0/reg0_b25  (
    .b({\PWM0/n12 [17],\PWM0/n12 [25]}),
    .c({freq0[17],freq0[25]}),
    .clk(clk100m),
    .d({\PWM0/n0_lutinv ,\PWM0/n0_lutinv }),
    .sr(\PWM0/n11 ),
    .q({\PWM0/FreCnt [17],\PWM0/FreCnt [25]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM0/reg0_b18|PWM0/reg0_b23  (
    .b({\PWM0/n12 [18],\PWM0/n12 [23]}),
    .c({freq0[18],freq0[23]}),
    .clk(clk100m),
    .d({\PWM0/n0_lutinv ,\PWM0/n0_lutinv }),
    .sr(\PWM0/n11 ),
    .q({\PWM0/FreCnt [18],\PWM0/FreCnt [23]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM0/reg0_b20|PWM0/reg0_b9  (
    .b({\PWM0/n12 [20],\PWM0/n12 [9]}),
    .c({freq0[20],freq0[9]}),
    .clk(clk100m),
    .d({\PWM0/n0_lutinv ,\PWM0/n0_lutinv }),
    .sr(\PWM0/n11 ),
    .q({\PWM0/FreCnt [20],\PWM0/FreCnt [9]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM0/reg0_b21|PWM0/reg0_b6  (
    .b({\PWM0/n12 [21],\PWM0/n12 [6]}),
    .c({freq0[21],freq0[6]}),
    .clk(clk100m),
    .d({\PWM0/n0_lutinv ,\PWM0/n0_lutinv }),
    .sr(\PWM0/n11 ),
    .q({\PWM0/FreCnt [21],\PWM0/FreCnt [6]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM0/reg0_b22|PWM0/reg0_b4  (
    .b({\PWM0/n12 [22],\PWM0/n12 [4]}),
    .c({freq0[22],freq0[4]}),
    .clk(clk100m),
    .d({\PWM0/n0_lutinv ,\PWM0/n0_lutinv }),
    .sr(\PWM0/n11 ),
    .q({\PWM0/FreCnt [22],\PWM0/FreCnt [4]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM0/reg0_b24|PWM0/reg0_b26  (
    .b({\PWM0/n12 [24],\PWM0/n12 [26]}),
    .c({freq0[24],freq0[26]}),
    .clk(clk100m),
    .d({\PWM0/n0_lutinv ,\PWM0/n0_lutinv }),
    .sr(\PWM0/n11 ),
    .q({\PWM0/FreCnt [24],\PWM0/FreCnt [26]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*B*A*~(0@D))"),
    //.LUTF1("(B*A*~(D@C))"),
    //.LUTG0("(C*B*A*~(1@D))"),
    //.LUTG1("(B*A*~(D@C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b1000000000001000),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b1000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg1_b10|PWM0/reg1_b7  (
    .a({_al_u1742_o,_al_u1744_o}),
    .b({_al_u1743_o,_al_u1746_o}),
    .c({\PWM0/FreCnt [9],_al_u1747_o}),
    .ce(\PWM0/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM0/FreCntr [10],\PWM0/FreCnt [6]}),
    .e({open_n319,\PWM0/FreCntr [7]}),
    .mi({freq0[10],freq0[7]}),
    .f({_al_u1744_o,_al_u1748_o}),
    .q({\PWM0/FreCntr [10],\PWM0/FreCntr [7]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~(D*~B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1100010011110101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg1_b13|PWM0/reg1_b0  (
    .a({\PWM0/FreCnt [12],open_n336}),
    .b({\PWM0/FreCnt [8],open_n337}),
    .c({\PWM0/FreCntr [13],\PWM0/n11 }),
    .ce(\PWM0/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM0/FreCntr [9],\PWM0/n0_lutinv }),
    .mi({freq0[13],freq0[0]}),
    .f({_al_u1743_o,\PWM0/mux3_b0_sel_is_3_o }),
    .q({\PWM0/FreCntr [13],\PWM0/FreCntr [0]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~A*~(0*~C)*~(D@B))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~A*~(1*~C)*~(D@B))"),
    //.LUTG1("(~C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100010000010001),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0100000000010000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg1_b14|PWM0/reg1_b11  (
    .a({open_n352,_al_u1753_o}),
    .b({open_n353,\PWM0/FreCnt [10]}),
    .c({\PWM0/FreCntr [14],\PWM0/FreCnt [16]}),
    .ce(\PWM0/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM0/FreCnt [13],\PWM0/FreCntr [11]}),
    .e({open_n354,\PWM0/FreCntr [17]}),
    .mi({freq0[14],freq0[11]}),
    .f({_al_u1753_o,_al_u1754_o}),
    .q({\PWM0/FreCntr [14],\PWM0/FreCntr [11]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~D*B)*~(~C*A))"),
    //.LUT1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111010100110001),
    .INIT_LUT1(16'b1000010000100001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg1_b15|PWM0/reg1_b9  (
    .a({\PWM0/FreCnt [14],\PWM0/FreCnt [0]}),
    .b({\PWM0/FreCnt [4],\PWM0/FreCnt [8]}),
    .c({\PWM0/FreCntr [15],\PWM0/FreCntr [1]}),
    .ce(\PWM0/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM0/FreCntr [5],\PWM0/FreCntr [9]}),
    .mi({freq0[15],freq0[9]}),
    .f({_al_u1749_o,_al_u1741_o}),
    .q({\PWM0/FreCntr [15],\PWM0/FreCntr [9]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~C*~(~0*B)*~(D@A))"),
    //.LUTF1("(A*~(0@C)*~(D@B))"),
    //.LUTG0("(~C*~(~1*B)*~(D@A))"),
    //.LUTG1("(A*~(1@C)*~(D@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000000001),
    .INIT_LUTF1(16'b0000100000000010),
    .INIT_LUTG0(16'b0000101000000101),
    .INIT_LUTG1(16'b1000000000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg1_b17|PWM0/reg1_b12  (
    .a({_al_u1360_o,\PWM0/FreCnt [11]}),
    .b(\PWM0/FreCnt [17:16]),
    .c({\PWM0/FreCnt [8],\PWM0/FreCnt [26]}),
    .ce(\PWM0/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM0/FreCntr [17],\PWM0/FreCntr [12]}),
    .e({\PWM0/FreCntr [8],\PWM0/FreCntr [17]}),
    .mi({freq0[17],freq0[12]}),
    .f({_al_u1361_o,_al_u1755_o}),
    .q({\PWM0/FreCntr [17],\PWM0/FreCntr [12]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(~0*C)*~(~D*B))"),
    //.LUTF1("(A*~(0*~C)*~(D*~B))"),
    //.LUTG0("(A*~(~1*C)*~(~D*B))"),
    //.LUTG1("(A*~(1*~C)*~(D*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101000000010),
    .INIT_LUTF1(16'b1000100010101010),
    .INIT_LUTG0(16'b1010101000100010),
    .INIT_LUTG1(16'b1000000010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg1_b18|PWM0/reg1_b16  (
    .a({_al_u1757_o,_al_u1761_o}),
    .b({\PWM0/FreCnt [17],\PWM0/FreCnt [15]}),
    .c({\PWM0/FreCnt [19],\PWM0/FreCnt [17]}),
    .ce(\PWM0/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM0/FreCntr [18],\PWM0/FreCntr [16]}),
    .e({\PWM0/FreCntr [20],\PWM0/FreCntr [18]}),
    .mi({freq0[18],freq0[16]}),
    .f({_al_u1758_o,_al_u1762_o}),
    .q({\PWM0/FreCntr [18],\PWM0/FreCntr [16]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*B*A*~(0@D))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(C*B*A*~(1@D))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg1_b19|PWM0/reg1_b3  (
    .a({\PWM0/FreCnt [18],_al_u1361_o}),
    .b({\PWM0/FreCnt [2],_al_u1363_o}),
    .c({\PWM0/FreCntr [19],_al_u1364_o}),
    .ce(\PWM0/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM0/FreCntr [3],\PWM0/FreCnt [3]}),
    .e({open_n417,\PWM0/FreCntr [3]}),
    .mi({freq0[19],freq0[3]}),
    .f({_al_u1751_o,_al_u1365_o}),
    .q({\PWM0/FreCntr [19],\PWM0/FreCntr [3]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(D@B)*~(C@A))"),
    //.LUT1("(D*~(C@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000010000100001),
    .INIT_LUT1(16'b1100001100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg1_b22|PWM0/reg1_b5  (
    .a({open_n434,\PWM0/FreCnt [18]}),
    .b({\PWM0/FreCnt [21],\PWM0/FreCnt [5]}),
    .c({\PWM0/FreCntr [22],\PWM0/FreCntr [18]}),
    .ce(\PWM0/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({_al_u1749_o,\PWM0/FreCntr [5]}),
    .mi({freq0[22],freq0[5]}),
    .f({_al_u1750_o,_al_u1364_o}),
    .q({\PWM0/FreCntr [22],\PWM0/FreCntr [5]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg1_b23|PWM0/reg1_b21  (
    .a({\PWM0/FreCnt [22],_al_u1751_o}),
    .b({\PWM0/FreCnt [23],\PWM0/FreCnt [20]}),
    .c({\PWM0/FreCntr [22],\PWM0/FreCnt [22]}),
    .ce(\PWM0/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM0/FreCntr [23],\PWM0/FreCntr [21]}),
    .e({open_n449,\PWM0/FreCntr [23]}),
    .mi({freq0[23],freq0[21]}),
    .f({_al_u1360_o,_al_u1752_o}),
    .q({\PWM0/FreCntr [23],\PWM0/FreCntr [21]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~A*~(0@C)*~(D*~B))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(~A*~(1@C)*~(D*~B))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010000000101),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b0100000001010000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg1_b25|PWM0/reg1_b1  (
    .a({\PWM0/FreCnt [11],_al_u1763_o}),
    .b({\PWM0/FreCnt [25],\PWM0/FreCnt [0]}),
    .c({\PWM0/FreCntr [11],\PWM0/FreCnt [24]}),
    .ce(\PWM0/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM0/FreCntr [25],\PWM0/FreCntr [1]}),
    .e({open_n466,\PWM0/FreCntr [25]}),
    .mi({freq0[25],freq0[1]}),
    .f({_al_u1373_o,_al_u1764_o}),
    .q({\PWM0/FreCntr [25],\PWM0/FreCntr [1]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~D*B)*~(~C*A))"),
    //.LUTF1("(~(~D*B)*~(C*~A))"),
    //.LUTG0("(~(~D*B)*~(~C*A))"),
    //.LUTG1("(~(~D*B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111010100110001),
    .INIT_LUTF1(16'b1010111100100011),
    .INIT_LUTG0(16'b1111010100110001),
    .INIT_LUTG1(16'b1010111100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg1_b2|PWM0/reg1_b26  (
    .a({\PWM0/FreCnt [1],\PWM0/FreCnt [1]}),
    .b({\PWM0/FreCnt [23],\PWM0/FreCnt [25]}),
    .c({\PWM0/FreCntr [2],\PWM0/FreCntr [2]}),
    .ce(\PWM0/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM0/FreCntr [24],\PWM0/FreCntr [26]}),
    .mi({freq0[2],freq0[26]}),
    .f({_al_u1761_o,_al_u1757_o}),
    .q({\PWM0/FreCntr [2],\PWM0/FreCntr [26]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(D*~B)*~(~C*A))"),
    //.LUT1("(~C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100010011110101),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg1_b4|PWM0/reg1_b20  (
    .a({open_n501,\PWM0/FreCnt [19]}),
    .b({open_n502,\PWM0/FreCnt [3]}),
    .c({\PWM0/FreCntr [4],\PWM0/FreCntr [20]}),
    .ce(\PWM0/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM0/FreCnt [3],\PWM0/FreCntr [4]}),
    .mi({freq0[4],freq0[20]}),
    .f({_al_u1763_o,_al_u1745_o}),
    .q({\PWM0/FreCntr [4],\PWM0/FreCntr [20]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(D*~B)*~(C*~A))"),
    //.LUT1("(~(~D*B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000110010101111),
    .INIT_LUT1(16'b1111010100110001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg1_b6|PWM0/reg1_b8  (
    .a({\PWM0/FreCnt [5],\PWM0/FreCnt [15]}),
    .b({\PWM0/FreCnt [7],\PWM0/FreCnt [7]}),
    .c({\PWM0/FreCntr [6],\PWM0/FreCntr [16]}),
    .ce(\PWM0/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM0/FreCntr [8],\PWM0/FreCntr [8]}),
    .mi({freq0[6],freq0[8]}),
    .f({_al_u1759_o,_al_u1747_o}),
    .q({\PWM0/FreCntr [6],\PWM0/FreCntr [8]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg2_b0|PWM0/reg3_b0  (
    .a({\PWM0/pnumr [0],_al_u1739_o}),
    .b({pnum0[0],\PWM0/n24 }),
    .c({pnum0[32],pnumcnt0[0]}),
    .clk(clk100m),
    .d({pwm_start_stop[16],\PWM0/pnumr [0]}),
    .e({open_n532,pwm_start_stop[16]}),
    .q({\PWM0/pnumr[0]_keep ,\PWM0/RemaTxNum[0]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011100010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011100010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg2_b10|PWM0/reg2_b9  (
    .a(\PWM0/pnumr [10:9]),
    .b({pnum0[10],pnum0[32]}),
    .c({pnum0[32],pnum0[9]}),
    .clk(clk100m),
    .d({pwm_start_stop[16],pwm_start_stop[16]}),
    .q({\PWM0/pnumr[10]_keep ,\PWM0/pnumr[9]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011100010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011100010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg2_b11|PWM0/reg2_b8  (
    .a({\PWM0/pnumr [11],\PWM0/pnumr [8]}),
    .b({pnum0[11],pnum0[32]}),
    .c({pnum0[32],pnum0[8]}),
    .clk(clk100m),
    .d({pwm_start_stop[16],pwm_start_stop[16]}),
    .q({\PWM0/pnumr[11]_keep ,\PWM0/pnumr[8]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg2_b12|PWM0/reg3_b12  (
    .a({\PWM0/pnumr [12],_al_u1731_o}),
    .b({pnum0[12],\PWM0/n24 }),
    .c({pnum0[32],pnumcnt0[12]}),
    .clk(clk100m),
    .d({pwm_start_stop[16],\PWM0/pnumr [12]}),
    .e({open_n600,pwm_start_stop[16]}),
    .q({\PWM0/pnumr[12]_keep ,\PWM0/RemaTxNum[12]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg2_b13|PWM0/reg3_b13  (
    .a({\PWM0/pnumr [13],_al_u1729_o}),
    .b({pnum0[13],\PWM0/n24 }),
    .c({pnum0[32],pnumcnt0[13]}),
    .clk(clk100m),
    .d({pwm_start_stop[16],\PWM0/pnumr [13]}),
    .e({open_n622,pwm_start_stop[16]}),
    .q({\PWM0/pnumr[13]_keep ,\PWM0/RemaTxNum[13]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011100010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg2_b14|PWM0/reg2_b5  (
    .a({\PWM0/pnumr [14],\PWM0/pnumr [5]}),
    .b({pnum0[14],pnum0[32]}),
    .c({pnum0[32],pnum0[5]}),
    .clk(clk100m),
    .d({pwm_start_stop[16],pwm_start_stop[16]}),
    .q({\PWM0/pnumr[14]_keep ,\PWM0/pnumr[5]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011100010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg2_b15|PWM0/reg2_b4  (
    .a({\PWM0/pnumr [15],\PWM0/pnumr [4]}),
    .b({pnum0[15],pnum0[32]}),
    .c({pnum0[32],pnum0[4]}),
    .clk(clk100m),
    .d({pwm_start_stop[16],pwm_start_stop[16]}),
    .q({\PWM0/pnumr[15]_keep ,\PWM0/pnumr[4]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg2_b16|PWM0/reg3_b16  (
    .a({\PWM0/pnumr [16],_al_u1723_o}),
    .b({pnum0[16],\PWM0/n24 }),
    .c({pnum0[32],pnumcnt0[16]}),
    .clk(clk100m),
    .d({pwm_start_stop[16],\PWM0/pnumr [16]}),
    .e({open_n682,pwm_start_stop[16]}),
    .q({\PWM0/pnumr[16]_keep ,\PWM0/RemaTxNum[16]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg2_b17|PWM0/reg3_b17  (
    .a({\PWM0/pnumr [17],_al_u1721_o}),
    .b({pnum0[17],\PWM0/n24 }),
    .c({pnum0[32],pnumcnt0[17]}),
    .clk(clk100m),
    .d({pwm_start_stop[16],\PWM0/pnumr [17]}),
    .e({open_n704,pwm_start_stop[16]}),
    .q({\PWM0/pnumr[17]_keep ,\PWM0/RemaTxNum[17]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg2_b18|PWM0/reg2_b22  (
    .a({\PWM0/pnumr [18],\PWM0/pnumr [22]}),
    .b({pnum0[18],pnum0[22]}),
    .c({pnum0[32],pnum0[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[16],pwm_start_stop[16]}),
    .q({\PWM0/pnumr[18]_keep ,\PWM0/pnumr[22]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg2_b19|PWM0/reg2_b21  (
    .a({\PWM0/pnumr [19],\PWM0/pnumr [21]}),
    .b({pnum0[19],pnum0[21]}),
    .c({pnum0[32],pnum0[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[16],pwm_start_stop[16]}),
    .q({\PWM0/pnumr[19]_keep ,\PWM0/pnumr[21]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg2_b1|PWM0/reg3_b1  (
    .a({\PWM0/pnumr [1],_al_u1737_o}),
    .b({pnum0[1],\PWM0/n24 }),
    .c({pnum0[32],pnumcnt0[1]}),
    .clk(clk100m),
    .d({pwm_start_stop[16],\PWM0/pnumr [1]}),
    .e({open_n772,pwm_start_stop[16]}),
    .q({\PWM0/pnumr[1]_keep ,\PWM0/RemaTxNum[1]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg2_b20|PWM0/reg3_b20  (
    .a({\PWM0/pnumr [20],_al_u1713_o}),
    .b({pnum0[20],\PWM0/n24 }),
    .c({pnum0[32],pnumcnt0[20]}),
    .clk(clk100m),
    .d({pwm_start_stop[16],\PWM0/pnumr [20]}),
    .e({open_n794,pwm_start_stop[16]}),
    .q({\PWM0/pnumr[20]_keep ,\PWM0/RemaTxNum[20]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg2_b23|PWM0/reg3_b23  (
    .a({\PWM0/pnumr [23],_al_u1707_o}),
    .b({pnum0[23],\PWM0/n24 }),
    .c({pnum0[32],pnumcnt0[23]}),
    .clk(clk100m),
    .d({pwm_start_stop[16],\PWM0/pnumr [23]}),
    .e({open_n816,pwm_start_stop[16]}),
    .q({\PWM0/pnumr[23]_keep ,\PWM0/RemaTxNum[23]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg2_b24|PWM0/reg2_b31  (
    .a({\PWM0/pnumr [24],\PWM0/pnumr [31]}),
    .b({pnum0[24],pnum0[31]}),
    .c({pnum0[32],pnum0[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[16],pwm_start_stop[16]}),
    .q({\PWM0/pnumr[24]_keep ,\PWM0/pnumr[31]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg2_b25|PWM0/reg2_b30  (
    .a({\PWM0/pnumr [25],\PWM0/pnumr [30]}),
    .b({pnum0[25],pnum0[30]}),
    .c({pnum0[32],pnum0[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[16],pwm_start_stop[16]}),
    .q({\PWM0/pnumr[25]_keep ,\PWM0/pnumr[30]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg2_b26|PWM0/reg2_b29  (
    .a({\PWM0/pnumr [26],\PWM0/pnumr [29]}),
    .b({pnum0[26],pnum0[29]}),
    .c({pnum0[32],pnum0[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[16],pwm_start_stop[16]}),
    .q({\PWM0/pnumr[26]_keep ,\PWM0/pnumr[29]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg2_b27|PWM0/reg2_b28  (
    .a({\PWM0/pnumr [27],\PWM0/pnumr [28]}),
    .b({pnum0[27],pnum0[28]}),
    .c({pnum0[32],pnum0[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[16],pwm_start_stop[16]}),
    .q({\PWM0/pnumr[27]_keep ,\PWM0/pnumr[28]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg2_b2|PWM0/reg3_b2  (
    .a({\PWM0/pnumr [2],_al_u1715_o}),
    .b({pnum0[2],\PWM0/n24 }),
    .c({pnum0[32],pnumcnt0[2]}),
    .clk(clk100m),
    .d({pwm_start_stop[16],\PWM0/pnumr [2]}),
    .e({open_n922,pwm_start_stop[16]}),
    .q({\PWM0/pnumr[2]_keep ,\PWM0/RemaTxNum[2]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg2_b3|PWM0/reg3_b3  (
    .a({\PWM0/pnumr [3],_al_u1705_o}),
    .b({pnum0[3],\PWM0/n24 }),
    .c({pnum0[32],pnumcnt0[3]}),
    .clk(clk100m),
    .d({pwm_start_stop[16],\PWM0/pnumr [3]}),
    .e({open_n944,pwm_start_stop[16]}),
    .q({\PWM0/pnumr[3]_keep ,\PWM0/RemaTxNum[3]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg2_b6|PWM0/reg3_b6  (
    .a({\PWM0/pnumr [6],_al_u1699_o}),
    .b({pnum0[32],\PWM0/n24 }),
    .c({pnum0[6],pnumcnt0[6]}),
    .clk(clk100m),
    .d({pwm_start_stop[16],\PWM0/pnumr [6]}),
    .e({open_n966,pwm_start_stop[16]}),
    .q({\PWM0/pnumr[6]_keep ,\PWM0/RemaTxNum[6]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg2_b7|PWM0/reg3_b7  (
    .a({\PWM0/pnumr [7],_al_u1697_o}),
    .b({pnum0[32],\PWM0/n24 }),
    .c({pnum0[7],pnumcnt0[7]}),
    .clk(clk100m),
    .d({pwm_start_stop[16],\PWM0/pnumr [7]}),
    .e({open_n988,pwm_start_stop[16]}),
    .q({\PWM0/pnumr[7]_keep ,\PWM0/RemaTxNum[7]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg3_b10  (
    .a({_al_u1735_o,_al_u1735_o}),
    .b({\PWM0/n24 ,\PWM0/n24 }),
    .c({pnumcnt0[10],pnumcnt0[10]}),
    .clk(clk100m),
    .d({\PWM0/pnumr [10],\PWM0/pnumr [10]}),
    .mi({open_n1020,pwm_start_stop[16]}),
    .q({open_n1027,\PWM0/RemaTxNum[10]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg3_b11  (
    .a({_al_u1733_o,_al_u1733_o}),
    .b({\PWM0/n24 ,\PWM0/n24 }),
    .c({pnumcnt0[11],pnumcnt0[11]}),
    .clk(clk100m),
    .d({\PWM0/pnumr [11],\PWM0/pnumr [11]}),
    .mi({open_n1039,pwm_start_stop[16]}),
    .q({open_n1046,\PWM0/RemaTxNum[11]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg3_b14  (
    .a({_al_u1727_o,_al_u1727_o}),
    .b({\PWM0/n24 ,\PWM0/n24 }),
    .c({pnumcnt0[14],pnumcnt0[14]}),
    .clk(clk100m),
    .d({\PWM0/pnumr [14],\PWM0/pnumr [14]}),
    .mi({open_n1058,pwm_start_stop[16]}),
    .q({open_n1065,\PWM0/RemaTxNum[14]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg3_b15  (
    .a({_al_u1725_o,_al_u1725_o}),
    .b({\PWM0/n24 ,\PWM0/n24 }),
    .c({pnumcnt0[15],pnumcnt0[15]}),
    .clk(clk100m),
    .d({\PWM0/pnumr [15],\PWM0/pnumr [15]}),
    .mi({open_n1077,pwm_start_stop[16]}),
    .q({open_n1084,\PWM0/RemaTxNum[15]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg3_b18  (
    .a({_al_u1719_o,_al_u1719_o}),
    .b({\PWM0/n24 ,\PWM0/n24 }),
    .c({pnumcnt0[18],pnumcnt0[18]}),
    .clk(clk100m),
    .d({\PWM0/pnumr [18],\PWM0/pnumr [18]}),
    .mi({open_n1096,pwm_start_stop[16]}),
    .q({open_n1103,\PWM0/RemaTxNum[18]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg3_b19  (
    .a({_al_u1717_o,_al_u1717_o}),
    .b({\PWM0/n24 ,\PWM0/n24 }),
    .c({pnumcnt0[19],pnumcnt0[19]}),
    .clk(clk100m),
    .d({\PWM0/pnumr [19],\PWM0/pnumr [19]}),
    .mi({open_n1115,pwm_start_stop[16]}),
    .q({open_n1122,\PWM0/RemaTxNum[19]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg3_b21  (
    .a({_al_u1711_o,_al_u1711_o}),
    .b({\PWM0/n24 ,\PWM0/n24 }),
    .c({pnumcnt0[21],pnumcnt0[21]}),
    .clk(clk100m),
    .d({\PWM0/pnumr [21],\PWM0/pnumr [21]}),
    .mi({open_n1134,pwm_start_stop[16]}),
    .q({open_n1141,\PWM0/RemaTxNum[21]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg3_b22  (
    .a({_al_u1709_o,_al_u1709_o}),
    .b({\PWM0/n24 ,\PWM0/n24 }),
    .c({pnumcnt0[22],pnumcnt0[22]}),
    .clk(clk100m),
    .d({\PWM0/pnumr [22],\PWM0/pnumr [22]}),
    .mi({open_n1153,pwm_start_stop[16]}),
    .q({open_n1160,\PWM0/RemaTxNum[22]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg3_b4  (
    .a({_al_u1703_o,_al_u1703_o}),
    .b({\PWM0/n24 ,\PWM0/n24 }),
    .c({pnumcnt0[4],pnumcnt0[4]}),
    .clk(clk100m),
    .d({\PWM0/pnumr [4],\PWM0/pnumr [4]}),
    .mi({open_n1172,pwm_start_stop[16]}),
    .q({open_n1179,\PWM0/RemaTxNum[4]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg3_b5  (
    .a({_al_u1701_o,_al_u1701_o}),
    .b({\PWM0/n24 ,\PWM0/n24 }),
    .c({pnumcnt0[5],pnumcnt0[5]}),
    .clk(clk100m),
    .d({\PWM0/pnumr [5],\PWM0/pnumr [5]}),
    .mi({open_n1191,pwm_start_stop[16]}),
    .q({open_n1198,\PWM0/RemaTxNum[5]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg3_b8  (
    .a({_al_u1695_o,_al_u1695_o}),
    .b({\PWM0/n24 ,\PWM0/n24 }),
    .c({pnumcnt0[8],pnumcnt0[8]}),
    .clk(clk100m),
    .d({\PWM0/pnumr [8],\PWM0/pnumr [8]}),
    .mi({open_n1210,pwm_start_stop[16]}),
    .q({open_n1217,\PWM0/RemaTxNum[8]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/reg3_b9  (
    .a({_al_u1693_o,_al_u1693_o}),
    .b({\PWM0/n24 ,\PWM0/n24 }),
    .c({pnumcnt0[9],pnumcnt0[9]}),
    .clk(clk100m),
    .d({\PWM0/pnumr [9],\PWM0/pnumr [9]}),
    .mi({open_n1229,pwm_start_stop[16]}),
    .q({open_n1236,\PWM0/RemaTxNum[9]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_LSLICE #(
    //.MACRO("PWM0/sub0/ucin_al_u3363"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM0/sub0/u11_al_u3366  (
    .a({\PWM0/FreCnt [13],\PWM0/FreCnt [11]}),
    .b({\PWM0/FreCnt [14],\PWM0/FreCnt [12]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM0/sub0/c11 ),
    .f({\PWM0/n12 [13],\PWM0/n12 [11]}),
    .fco(\PWM0/sub0/c15 ),
    .fx({\PWM0/n12 [14],\PWM0/n12 [12]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM0/sub0/ucin_al_u3363"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM0/sub0/u15_al_u3367  (
    .a({\PWM0/FreCnt [17],\PWM0/FreCnt [15]}),
    .b({\PWM0/FreCnt [18],\PWM0/FreCnt [16]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM0/sub0/c15 ),
    .f({\PWM0/n12 [17],\PWM0/n12 [15]}),
    .fco(\PWM0/sub0/c19 ),
    .fx({\PWM0/n12 [18],\PWM0/n12 [16]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM0/sub0/ucin_al_u3363"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM0/sub0/u19_al_u3368  (
    .a({\PWM0/FreCnt [21],\PWM0/FreCnt [19]}),
    .b({\PWM0/FreCnt [22],\PWM0/FreCnt [20]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM0/sub0/c19 ),
    .f({\PWM0/n12 [21],\PWM0/n12 [19]}),
    .fco(\PWM0/sub0/c23 ),
    .fx({\PWM0/n12 [22],\PWM0/n12 [20]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM0/sub0/ucin_al_u3363"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM0/sub0/u23_al_u3369  (
    .a({\PWM0/FreCnt [25],\PWM0/FreCnt [23]}),
    .b({\PWM0/FreCnt [26],\PWM0/FreCnt [24]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM0/sub0/c23 ),
    .f({\PWM0/n12 [25],\PWM0/n12 [23]}),
    .fx({\PWM0/n12 [26],\PWM0/n12 [24]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM0/sub0/ucin_al_u3363"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM0/sub0/u3_al_u3364  (
    .a({\PWM0/FreCnt [5],\PWM0/FreCnt [3]}),
    .b({\PWM0/FreCnt [6],\PWM0/FreCnt [4]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM0/sub0/c3 ),
    .f({\PWM0/n12 [5],\PWM0/n12 [3]}),
    .fco(\PWM0/sub0/c7 ),
    .fx({\PWM0/n12 [6],\PWM0/n12 [4]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM0/sub0/ucin_al_u3363"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM0/sub0/u7_al_u3365  (
    .a({\PWM0/FreCnt [9],\PWM0/FreCnt [7]}),
    .b({\PWM0/FreCnt [10],\PWM0/FreCnt [8]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM0/sub0/c7 ),
    .f({\PWM0/n12 [9],\PWM0/n12 [7]}),
    .fco(\PWM0/sub0/c11 ),
    .fx({\PWM0/n12 [10],\PWM0/n12 [8]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM0/sub0/ucin_al_u3363"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'h0005),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/sub0/ucin_al_u3363  (
    .a({\PWM0/FreCnt [1],1'b0}),
    .b({\PWM0/FreCnt [2],\PWM0/FreCnt [0]}),
    .c(2'b11),
    .ce(\U_AHB/n2 ),
    .clk(clk100m),
    .d(2'b01),
    .e(2'b01),
    .mi({open_n1347,\U_AHB/h2h_hwdata [2]}),
    .f({\PWM0/n12 [1],open_n1360}),
    .fco(\PWM0/sub0/c3 ),
    .fx({\PWM0/n12 [2],\PWM0/n12 [0]}),
    .q({open_n1361,freq0[2]}));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM0/sub1/u0|PWM0/sub1/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("SUB_CARRY"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000101),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM0/sub1/u0|PWM0/sub1/ucin  (
    .a({pnumcnt0[0],1'b0}),
    .b({1'b1,open_n1362}),
    .ce(\U_AHB/n10 ),
    .clk(clk100m),
    .mi({\U_AHB/h2h_hwdata [4],\U_AHB/h2h_hwdata [26]}),
    .f({\PWM0/n26 [0],open_n1378}),
    .fco(\PWM0/sub1/c1 ),
    .q({freq3[4],freq3[26]}));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM0/sub1/u0|PWM0/sub1/ucin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM0/sub1/u10|PWM0/sub1/u9  (
    .a(pnumcnt0[10:9]),
    .b(2'b00),
    .fci(\PWM0/sub1/c9 ),
    .f(\PWM0/n26 [10:9]),
    .fco(\PWM0/sub1/c11 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM0/sub1/u0|PWM0/sub1/ucin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM0/sub1/u12|PWM0/sub1/u11  (
    .a(pnumcnt0[12:11]),
    .b(2'b00),
    .fci(\PWM0/sub1/c11 ),
    .f(\PWM0/n26 [12:11]),
    .fco(\PWM0/sub1/c13 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM0/sub1/u0|PWM0/sub1/ucin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM0/sub1/u14|PWM0/sub1/u13  (
    .a(pnumcnt0[14:13]),
    .b(2'b00),
    .fci(\PWM0/sub1/c13 ),
    .f(\PWM0/n26 [14:13]),
    .fco(\PWM0/sub1/c15 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM0/sub1/u0|PWM0/sub1/ucin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM0/sub1/u16|PWM0/sub1/u15  (
    .a(pnumcnt0[16:15]),
    .b(2'b00),
    .fci(\PWM0/sub1/c15 ),
    .f(\PWM0/n26 [16:15]),
    .fco(\PWM0/sub1/c17 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM0/sub1/u0|PWM0/sub1/ucin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM0/sub1/u18|PWM0/sub1/u17  (
    .a(pnumcnt0[18:17]),
    .b(2'b00),
    .fci(\PWM0/sub1/c17 ),
    .f(\PWM0/n26 [18:17]),
    .fco(\PWM0/sub1/c19 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM0/sub1/u0|PWM0/sub1/ucin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM0/sub1/u20|PWM0/sub1/u19  (
    .a(pnumcnt0[20:19]),
    .b(2'b00),
    .fci(\PWM0/sub1/c19 ),
    .f(\PWM0/n26 [20:19]),
    .fco(\PWM0/sub1/c21 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM0/sub1/u0|PWM0/sub1/ucin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM0/sub1/u22|PWM0/sub1/u21  (
    .a(pnumcnt0[22:21]),
    .b(2'b00),
    .fci(\PWM0/sub1/c21 ),
    .f(\PWM0/n26 [22:21]),
    .fco(\PWM0/sub1/c23 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM0/sub1/u0|PWM0/sub1/ucin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM0/sub1/u23_al_u3468  (
    .a({open_n1535,pnumcnt0[23]}),
    .b({open_n1536,1'b0}),
    .fci(\PWM0/sub1/c23 ),
    .f({open_n1555,\PWM0/n26 [23]}));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM0/sub1/u0|PWM0/sub1/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM0/sub1/u2|PWM0/sub1/u1  (
    .a(pnumcnt0[2:1]),
    .b(2'b00),
    .fci(\PWM0/sub1/c1 ),
    .f(\PWM0/n26 [2:1]),
    .fco(\PWM0/sub1/c3 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM0/sub1/u0|PWM0/sub1/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM0/sub1/u4|PWM0/sub1/u3  (
    .a(pnumcnt0[4:3]),
    .b(2'b00),
    .fci(\PWM0/sub1/c3 ),
    .f(\PWM0/n26 [4:3]),
    .fco(\PWM0/sub1/c5 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM0/sub1/u0|PWM0/sub1/ucin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM0/sub1/u6|PWM0/sub1/u5  (
    .a(pnumcnt0[6:5]),
    .b(2'b00),
    .fci(\PWM0/sub1/c5 ),
    .f(\PWM0/n26 [6:5]),
    .fco(\PWM0/sub1/c7 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM0/sub1/u0|PWM0/sub1/ucin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM0/sub1/u8|PWM0/sub1/u7  (
    .a(pnumcnt0[8:7]),
    .b(2'b00),
    .fci(\PWM0/sub1/c7 ),
    .f(\PWM0/n26 [8:7]),
    .fco(\PWM0/sub1/c9 ));
  // src/OnePWM.v(26)
  // src/OnePWM.v(26)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*~(~D*B*~A))"),
    //.LUTF1("(C*~(~D*B*~A))"),
    //.LUTG0("(C*~(~D*B*~A))"),
    //.LUTG1("(C*~(~D*B*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000010110000),
    .INIT_LUTF1(16'b1111000010110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \PWM1/State_reg|PWME/State_reg  (
    .a({_al_u3010_o,_al_u3049_o}),
    .b({\PWM1/n0_lutinv ,\PWME/n0_lutinv }),
    .c({_al_u3011_o,_al_u3050_o}),
    .clk(clk100m),
    .d({pwm_start_stop[17],pwm_start_stop[30]}),
    .sr(rstn),
    .q({pwm_state_read[1],pwm_state_read[14]}));  // src/OnePWM.v(26)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[0]  (
    .i(\PWM1/RemaTxNum[0]_keep ),
    .o(pnumcnt1[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[10]  (
    .i(\PWM1/RemaTxNum[10]_keep ),
    .o(pnumcnt1[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[11]  (
    .i(\PWM1/RemaTxNum[11]_keep ),
    .o(pnumcnt1[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[12]  (
    .i(\PWM1/RemaTxNum[12]_keep ),
    .o(pnumcnt1[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[13]  (
    .i(\PWM1/RemaTxNum[13]_keep ),
    .o(pnumcnt1[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[14]  (
    .i(\PWM1/RemaTxNum[14]_keep ),
    .o(pnumcnt1[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[15]  (
    .i(\PWM1/RemaTxNum[15]_keep ),
    .o(pnumcnt1[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[16]  (
    .i(\PWM1/RemaTxNum[16]_keep ),
    .o(pnumcnt1[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[17]  (
    .i(\PWM1/RemaTxNum[17]_keep ),
    .o(pnumcnt1[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[18]  (
    .i(\PWM1/RemaTxNum[18]_keep ),
    .o(pnumcnt1[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[19]  (
    .i(\PWM1/RemaTxNum[19]_keep ),
    .o(pnumcnt1[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[1]  (
    .i(\PWM1/RemaTxNum[1]_keep ),
    .o(pnumcnt1[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[20]  (
    .i(\PWM1/RemaTxNum[20]_keep ),
    .o(pnumcnt1[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[21]  (
    .i(\PWM1/RemaTxNum[21]_keep ),
    .o(pnumcnt1[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[22]  (
    .i(\PWM1/RemaTxNum[22]_keep ),
    .o(pnumcnt1[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[23]  (
    .i(\PWM1/RemaTxNum[23]_keep ),
    .o(pnumcnt1[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[2]  (
    .i(\PWM1/RemaTxNum[2]_keep ),
    .o(pnumcnt1[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[3]  (
    .i(\PWM1/RemaTxNum[3]_keep ),
    .o(pnumcnt1[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[4]  (
    .i(\PWM1/RemaTxNum[4]_keep ),
    .o(pnumcnt1[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[5]  (
    .i(\PWM1/RemaTxNum[5]_keep ),
    .o(pnumcnt1[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[6]  (
    .i(\PWM1/RemaTxNum[6]_keep ),
    .o(pnumcnt1[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[7]  (
    .i(\PWM1/RemaTxNum[7]_keep ),
    .o(pnumcnt1[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[8]  (
    .i(\PWM1/RemaTxNum[8]_keep ),
    .o(pnumcnt1[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[9]  (
    .i(\PWM1/RemaTxNum[9]_keep ),
    .o(pnumcnt1[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_dir  (
    .i(\PWM1/dir_keep ),
    .o(dir_pad[1]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[0]  (
    .i(\PWM1/pnumr[0]_keep ),
    .o(\PWM1/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[10]  (
    .i(\PWM1/pnumr[10]_keep ),
    .o(\PWM1/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[11]  (
    .i(\PWM1/pnumr[11]_keep ),
    .o(\PWM1/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[12]  (
    .i(\PWM1/pnumr[12]_keep ),
    .o(\PWM1/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[13]  (
    .i(\PWM1/pnumr[13]_keep ),
    .o(\PWM1/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[14]  (
    .i(\PWM1/pnumr[14]_keep ),
    .o(\PWM1/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[15]  (
    .i(\PWM1/pnumr[15]_keep ),
    .o(\PWM1/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[16]  (
    .i(\PWM1/pnumr[16]_keep ),
    .o(\PWM1/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[17]  (
    .i(\PWM1/pnumr[17]_keep ),
    .o(\PWM1/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[18]  (
    .i(\PWM1/pnumr[18]_keep ),
    .o(\PWM1/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[19]  (
    .i(\PWM1/pnumr[19]_keep ),
    .o(\PWM1/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[1]  (
    .i(\PWM1/pnumr[1]_keep ),
    .o(\PWM1/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[20]  (
    .i(\PWM1/pnumr[20]_keep ),
    .o(\PWM1/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[21]  (
    .i(\PWM1/pnumr[21]_keep ),
    .o(\PWM1/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[22]  (
    .i(\PWM1/pnumr[22]_keep ),
    .o(\PWM1/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[23]  (
    .i(\PWM1/pnumr[23]_keep ),
    .o(\PWM1/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[24]  (
    .i(\PWM1/pnumr[24]_keep ),
    .o(\PWM1/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[25]  (
    .i(\PWM1/pnumr[25]_keep ),
    .o(\PWM1/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[26]  (
    .i(\PWM1/pnumr[26]_keep ),
    .o(\PWM1/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[27]  (
    .i(\PWM1/pnumr[27]_keep ),
    .o(\PWM1/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[28]  (
    .i(\PWM1/pnumr[28]_keep ),
    .o(\PWM1/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[29]  (
    .i(\PWM1/pnumr[29]_keep ),
    .o(\PWM1/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[2]  (
    .i(\PWM1/pnumr[2]_keep ),
    .o(\PWM1/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[30]  (
    .i(\PWM1/pnumr[30]_keep ),
    .o(\PWM1/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[31]  (
    .i(\PWM1/pnumr[31]_keep ),
    .o(\PWM1/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[3]  (
    .i(\PWM1/pnumr[3]_keep ),
    .o(\PWM1/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[4]  (
    .i(\PWM1/pnumr[4]_keep ),
    .o(\PWM1/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[5]  (
    .i(\PWM1/pnumr[5]_keep ),
    .o(\PWM1/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[6]  (
    .i(\PWM1/pnumr[6]_keep ),
    .o(\PWM1/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[7]  (
    .i(\PWM1/pnumr[7]_keep ),
    .o(\PWM1/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[8]  (
    .i(\PWM1/pnumr[8]_keep ),
    .o(\PWM1/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[9]  (
    .i(\PWM1/pnumr[9]_keep ),
    .o(\PWM1/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pwm  (
    .i(\PWM1/pwm_keep ),
    .o(pwm_pad[1]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_stopreq  (
    .i(\PWM1/stopreq_keep ),
    .o(\PWM1/stopreq ));  // src/OnePWM.v(14)
  EF2_PHY_MSLICE #(
    //.LUT0("(D*~(C)*~((~0*~(B*A)))+D*C*~((~0*~(B*A)))+~(D)*C*(~0*~(B*A))+D*C*(~0*~(B*A)))"),
    //.LUT1("(D*~(C)*~((~1*~(B*A)))+D*C*~((~1*~(B*A)))+~(D)*C*(~1*~(B*A))+D*C*(~1*~(B*A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111100001110000),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/dir_reg  (
    .a({\PWM1/n24 ,\PWM1/n24 }),
    .b({\PWM1/n25_neg_lutinv ,\PWM1/n25_neg_lutinv }),
    .c({dir_pad[1],dir_pad[1]}),
    .clk(clk100m),
    .d({\PWM1/pnumr [31],\PWM1/pnumr [31]}),
    .mi({open_n1682,pwm_start_stop[17]}),
    .q({open_n1689,\PWM1/dir_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("~(~0*~(D*C*B*A))"),
    //.LUT1("~(~1*~(D*C*B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b1111111111111111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM1/pwm_reg  (
    .a({_al_u1383_o,_al_u1383_o}),
    .b({_al_u1389_o,_al_u1389_o}),
    .c({_al_u1391_o,_al_u1391_o}),
    .clk(clk100m),
    .d({_al_u1393_o,_al_u1393_o}),
    .mi({open_n1701,pwm_pad[1]}),
    .sr(\PWM1/u14_sel_is_1_o ),
    .q({open_n1707,\PWM1/pwm_keep }));  // src/OnePWM.v(45)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM1/reg0_b0|PWM1/reg0_b12  (
    .b({\PWM1/n12 [0],\PWM1/n12 [12]}),
    .c({freq1[0],freq1[12]}),
    .clk(clk100m),
    .d({\PWM1/n0_lutinv ,\PWM1/n0_lutinv }),
    .sr(\PWM1/n11 ),
    .q({\PWM1/FreCnt [0],\PWM1/FreCnt [12]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM1/reg0_b10|PWM1/reg0_b8  (
    .b({\PWM1/n12 [10],\PWM1/n12 [8]}),
    .c({freq1[10],freq1[8]}),
    .clk(clk100m),
    .d({\PWM1/n0_lutinv ,\PWM1/n0_lutinv }),
    .sr(\PWM1/n11 ),
    .q({\PWM1/FreCnt [10],\PWM1/FreCnt [8]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM1/reg0_b11|PWM1/reg0_b7  (
    .b({\PWM1/n12 [11],\PWM1/n12 [7]}),
    .c({freq1[11],freq1[7]}),
    .clk(clk100m),
    .d({\PWM1/n0_lutinv ,\PWM1/n0_lutinv }),
    .sr(\PWM1/n11 ),
    .q({\PWM1/FreCnt [11],\PWM1/FreCnt [7]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM1/reg0_b13|PWM1/reg0_b3  (
    .b({\PWM1/n12 [13],\PWM1/n12 [3]}),
    .c({freq1[13],freq1[3]}),
    .clk(clk100m),
    .d({\PWM1/n0_lutinv ,\PWM1/n0_lutinv }),
    .sr(\PWM1/n11 ),
    .q({\PWM1/FreCnt [13],\PWM1/FreCnt [3]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM1/reg0_b14|PWM1/reg0_b25  (
    .b({\PWM1/n12 [14],\PWM1/n12 [25]}),
    .c({freq1[14],freq1[25]}),
    .clk(clk100m),
    .d({\PWM1/n0_lutinv ,\PWM1/n0_lutinv }),
    .sr(\PWM1/n11 ),
    .q({\PWM1/FreCnt [14],\PWM1/FreCnt [25]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM1/reg0_b16|PWM1/reg0_b23  (
    .b({\PWM1/n12 [16],\PWM1/n12 [23]}),
    .c({freq1[16],freq1[23]}),
    .clk(clk100m),
    .d({\PWM1/n0_lutinv ,\PWM1/n0_lutinv }),
    .sr(\PWM1/n11 ),
    .q({\PWM1/FreCnt [16],\PWM1/FreCnt [23]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM1/reg0_b17|PWM1/reg0_b21  (
    .b({\PWM1/n12 [17],\PWM1/n12 [21]}),
    .c({freq1[17],freq1[21]}),
    .clk(clk100m),
    .d({\PWM1/n0_lutinv ,\PWM1/n0_lutinv }),
    .sr(\PWM1/n11 ),
    .q({\PWM1/FreCnt [17],\PWM1/FreCnt [21]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM1/reg0_b18|PWM1/reg0_b19  (
    .b({\PWM1/n12 [18],\PWM1/n12 [19]}),
    .c({freq1[18],freq1[19]}),
    .clk(clk100m),
    .d({\PWM1/n0_lutinv ,\PWM1/n0_lutinv }),
    .sr(\PWM1/n11 ),
    .q({\PWM1/FreCnt [18],\PWM1/FreCnt [19]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM1/reg0_b20|PWM1/reg0_b1  (
    .b({\PWM1/n12 [20],\PWM1/n12 [1]}),
    .c({freq1[20],freq1[1]}),
    .clk(clk100m),
    .d({\PWM1/n0_lutinv ,\PWM1/n0_lutinv }),
    .sr(\PWM1/n11 ),
    .q({\PWM1/FreCnt [20],\PWM1/FreCnt [1]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM1/reg0_b22|PWM1/reg0_b9  (
    .b({\PWM1/n12 [22],\PWM1/n12 [9]}),
    .c({freq1[22],freq1[9]}),
    .clk(clk100m),
    .d({\PWM1/n0_lutinv ,\PWM1/n0_lutinv }),
    .sr(\PWM1/n11 ),
    .q({\PWM1/FreCnt [22],\PWM1/FreCnt [9]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM1/reg0_b24|PWM1/reg0_b6  (
    .b({\PWM1/n12 [24],\PWM1/n12 [6]}),
    .c({freq1[24],freq1[6]}),
    .clk(clk100m),
    .d({\PWM1/n0_lutinv ,\PWM1/n0_lutinv }),
    .sr(\PWM1/n11 ),
    .q({\PWM1/FreCnt [24],\PWM1/FreCnt [6]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM1/reg0_b26|PWM1/reg0_b5  (
    .b({\PWM1/n12 [26],\PWM1/n12 [5]}),
    .c({freq1[26],freq1[5]}),
    .clk(clk100m),
    .d({\PWM1/n0_lutinv ,\PWM1/n0_lutinv }),
    .sr(\PWM1/n11 ),
    .q({\PWM1/FreCnt [26],\PWM1/FreCnt [5]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM1/reg0_b2|PWM1/reg0_b4  (
    .b({\PWM1/n12 [2],\PWM1/n12 [4]}),
    .c({freq1[2],freq1[4]}),
    .clk(clk100m),
    .d({\PWM1/n0_lutinv ,\PWM1/n0_lutinv }),
    .sr(\PWM1/n11 ),
    .q({\PWM1/FreCnt [2],\PWM1/FreCnt [4]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~A*~(0*~C)*~(D@B))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(~A*~(1*~C)*~(D@B))"),
    //.LUTG1("(C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100010000010001),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0100000000010000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg1_b11|PWM1/reg1_b23  (
    .a({open_n1996,_al_u1834_o}),
    .b({open_n1997,\PWM1/FreCnt [22]}),
    .c({\PWM1/FreCntr [11],\PWM1/FreCnt [3]}),
    .ce(\PWM1/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM1/FreCnt [10],\PWM1/FreCntr [23]}),
    .e({open_n1998,\PWM1/FreCntr [4]}),
    .mi({freq1[11],freq1[23]}),
    .f({_al_u1834_o,_al_u1835_o}),
    .q({\PWM1/FreCntr [11],\PWM1/FreCntr [23]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(~D*B))"),
    //.LUTF1("(~(D*~B)*~(C*~A))"),
    //.LUTG0("(A*~(1@C)*~(~D*B))"),
    //.LUTG1("(~(D*~B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101000000010),
    .INIT_LUTF1(16'b1000110010101111),
    .INIT_LUTG0(16'b1010000000100000),
    .INIT_LUTG1(16'b1000110010101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg1_b12|PWM1/reg1_b15  (
    .a({\PWM1/FreCnt [12],_al_u1824_o}),
    .b({\PWM1/FreCnt [15],\PWM1/FreCnt [12]}),
    .c({\PWM1/FreCntr [12],\PWM1/FreCnt [14]}),
    .ce(\PWM1/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM1/FreCntr [15],\PWM1/FreCntr [13]}),
    .e({open_n2015,\PWM1/FreCntr [15]}),
    .mi({freq1[12],freq1[15]}),
    .f({_al_u1387_o,_al_u1825_o}),
    .q({\PWM1/FreCntr [12],\PWM1/FreCntr [15]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(D*~B)*~(C*~A))"),
    //.LUTF1("(~(~D*B)*~(~C*A))"),
    //.LUTG0("(~(D*~B)*~(C*~A))"),
    //.LUTG1("(~(~D*B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000110010101111),
    .INIT_LUTF1(16'b1111010100110001),
    .INIT_LUTG0(16'b1000110010101111),
    .INIT_LUTG1(16'b1111010100110001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg1_b14|PWM1/reg1_b8  (
    .a({\PWM1/FreCnt [13],\PWM1/FreCnt [7]}),
    .b({\PWM1/FreCnt [7],\PWM1/FreCnt [8]}),
    .c({\PWM1/FreCntr [14],\PWM1/FreCntr [8]}),
    .ce(\PWM1/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM1/FreCntr [8],\PWM1/FreCntr [9]}),
    .mi({freq1[14],freq1[8]}),
    .f({_al_u1830_o,_al_u1845_o}),
    .q({\PWM1/FreCntr [14],\PWM1/FreCntr [8]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~B*~(0@C)*~(D*~A))"),
    //.LUTF1("(~(~D*B)*~(C*~A))"),
    //.LUTG0("(~B*~(1@C)*~(D*~A))"),
    //.LUTG1("(~(~D*B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000000011),
    .INIT_LUTF1(16'b1010111100100011),
    .INIT_LUTG0(16'b0010000000110000),
    .INIT_LUTG1(16'b1010111100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg1_b16|PWM1/reg1_b20  (
    .a({\PWM1/FreCnt [15],\PWM1/FreCnt [19]}),
    .b({\PWM1/FreCnt [19],\PWM1/FreCnt [26]}),
    .c({\PWM1/FreCntr [16],\PWM1/FreCnt [4]}),
    .ce(\PWM1/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM1/FreCntr [20],\PWM1/FreCntr [20]}),
    .e({open_n2050,\PWM1/FreCntr [5]}),
    .mi({freq1[16],freq1[20]}),
    .f({_al_u1843_o,_al_u1839_o}),
    .q({\PWM1/FreCntr [16],\PWM1/FreCntr [20]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*B*A*~(0@D))"),
    //.LUTF1("(D*~(C@B))"),
    //.LUTG0("(C*B*A*~(1@D))"),
    //.LUTG1("(D*~(C@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b1100001100000000),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b1100001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg1_b17|PWM1/reg1_b10  (
    .a({open_n2067,_al_u1825_o}),
    .b({\PWM1/FreCnt [16],_al_u1827_o}),
    .c({\PWM1/FreCntr [17],_al_u1828_o}),
    .ce(\PWM1/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({_al_u1826_o,\PWM1/FreCnt [9]}),
    .e({open_n2068,\PWM1/FreCntr [10]}),
    .mi({freq1[17],freq1[10]}),
    .f({_al_u1827_o,_al_u1829_o}),
    .q({\PWM1/FreCntr [17],\PWM1/FreCntr [10]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(~0*C)*~(D*~B))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(A*~(~1*C)*~(D*~B))"),
    //.LUTG1("(~C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000001010),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1000100010101010),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg1_b19|PWM1/reg1_b24  (
    .a({open_n2085,_al_u1830_o}),
    .b({open_n2086,\PWM1/FreCnt [18]}),
    .c({\PWM1/FreCntr [19],\PWM1/FreCnt [23]}),
    .ce(\PWM1/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM1/FreCnt [18],\PWM1/FreCntr [19]}),
    .e({open_n2087,\PWM1/FreCntr [24]}),
    .mi({freq1[19],freq1[24]}),
    .f({_al_u1836_o,_al_u1831_o}),
    .q({\PWM1/FreCntr [19],\PWM1/FreCntr [24]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(D*~B)*~(C*~A))"),
    //.LUT1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000110010101111),
    .INIT_LUT1(16'b1000010000100001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg1_b1|PWM1/reg1_b18  (
    .a({\PWM1/FreCnt [0],\PWM1/FreCnt [13]}),
    .b({\PWM1/FreCnt [11],\PWM1/FreCnt [17]}),
    .c({\PWM1/FreCntr [1],\PWM1/FreCntr [14]}),
    .ce(\PWM1/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM1/FreCntr [12],\PWM1/FreCntr [18]}),
    .mi({freq1[1],freq1[18]}),
    .f({_al_u1841_o,_al_u1828_o}),
    .q({\PWM1/FreCntr [1],\PWM1/FreCntr [18]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(~0*C)*~(D*~B))"),
    //.LUTF1("(A*~(~0*C)*~(~D*B))"),
    //.LUTG0("(A*~(~1*C)*~(D*~B))"),
    //.LUTG1("(A*~(~1*C)*~(~D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000001010),
    .INIT_LUTF1(16'b0000101000000010),
    .INIT_LUTG0(16'b1000100010101010),
    .INIT_LUTG1(16'b1010101000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg1_b22|PWM1/reg1_b26  (
    .a({_al_u1845_o,_al_u1843_o}),
    .b({\PWM1/FreCnt [21],\PWM1/FreCnt [25]}),
    .c({\PWM1/FreCnt [25],\PWM1/FreCnt [3]}),
    .ce(\PWM1/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM1/FreCntr [22],\PWM1/FreCntr [26]}),
    .e({\PWM1/FreCntr [26],\PWM1/FreCntr [4]}),
    .mi({freq1[22],freq1[26]}),
    .f({_al_u1846_o,_al_u1844_o}),
    .q({\PWM1/FreCntr [22],\PWM1/FreCntr [26]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(A*~(0@C)*~(D@B))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(A*~(1@C)*~(D@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b0000100000000010),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000000000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg1_b25|PWM1/reg1_b7  (
    .a({_al_u1839_o,_al_u1378_o}),
    .b({\PWM1/FreCnt [24],\PWM1/FreCnt [7]}),
    .c({\PWM1/FreCnt [6],\PWM1/FreCnt [9]}),
    .ce(\PWM1/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM1/FreCntr [25],\PWM1/FreCntr [7]}),
    .e({\PWM1/FreCntr [7],\PWM1/FreCntr [9]}),
    .mi({freq1[25],freq1[7]}),
    .f({_al_u1840_o,_al_u1379_o}),
    .q({\PWM1/FreCntr [25],\PWM1/FreCntr [7]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~A*~(~0*C)*~(D@B))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(~A*~(~1*C)*~(D@B))"),
    //.LUTG1("(C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010000000001),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0100010000010001),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg1_b2|PWM1/reg1_b6  (
    .a({open_n2150,_al_u1832_o}),
    .b({open_n2151,\PWM1/FreCnt [5]}),
    .c({\PWM1/FreCntr [2],\PWM1/FreCnt [8]}),
    .ce(\PWM1/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM1/FreCnt [1],\PWM1/FreCntr [6]}),
    .e({open_n2152,\PWM1/FreCntr [9]}),
    .mi({freq1[2],freq1[6]}),
    .f({_al_u1832_o,_al_u1833_o}),
    .q({\PWM1/FreCntr [2],\PWM1/FreCntr [6]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*B*A*~(0@D))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(C*B*A*~(1@D))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg1_b5|PWM1/reg1_b4  (
    .a({\PWM1/FreCnt [18],_al_u1379_o}),
    .b({\PWM1/FreCnt [5],_al_u1381_o}),
    .c({\PWM1/FreCntr [18],_al_u1382_o}),
    .ce(\PWM1/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM1/FreCntr [5],\PWM1/FreCnt [4]}),
    .e({open_n2169,\PWM1/FreCntr [4]}),
    .mi(freq1[5:4]),
    .f({_al_u1382_o,_al_u1383_o}),
    .q(\PWM1/FreCntr [5:4]));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg1_b9|PWM1/reg1_b0  (
    .b({_al_u775_o,open_n2188}),
    .c({_al_u777_o,\PWM1/n11 }),
    .ce(\PWM1/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({_al_u773_o,\PWM1/n0_lutinv }),
    .mi({freq1[9],freq1[0]}),
    .f({\PWM1/n0_lutinv ,\PWM1/mux3_b0_sel_is_3_o }),
    .q({\PWM1/FreCntr [9],\PWM1/FreCntr [0]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011100010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg2_b0|PWM1/reg2_b9  (
    .a({\PWM1/pnumr [0],\PWM1/pnumr [9]}),
    .b({pnum1[0],pnum1[32]}),
    .c({pnum1[32],pnum1[9]}),
    .clk(clk100m),
    .d({pwm_start_stop[17],pwm_start_stop[17]}),
    .q({\PWM1/pnumr[0]_keep ,\PWM1/pnumr[9]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg2_b10|PWM1/reg3_b10  (
    .a({\PWM1/pnumr [10],_al_u1817_o}),
    .b({pnum1[10],\PWM1/n24 }),
    .c({pnum1[32],pnumcnt1[10]}),
    .clk(clk100m),
    .d({pwm_start_stop[17],\PWM1/pnumr [10]}),
    .e({open_n2223,pwm_start_stop[17]}),
    .q({\PWM1/pnumr[10]_keep ,\PWM1/RemaTxNum[10]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011100010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg2_b11|PWM1/reg2_b6  (
    .a({\PWM1/pnumr [11],\PWM1/pnumr [6]}),
    .b({pnum1[11],pnum1[32]}),
    .c({pnum1[32],pnum1[6]}),
    .clk(clk100m),
    .d({pwm_start_stop[17],pwm_start_stop[17]}),
    .q({\PWM1/pnumr[11]_keep ,\PWM1/pnumr[6]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011100010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011100010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg2_b12|PWM1/reg2_b5  (
    .a({\PWM1/pnumr [12],\PWM1/pnumr [5]}),
    .b({pnum1[12],pnum1[32]}),
    .c({pnum1[32],pnum1[5]}),
    .clk(clk100m),
    .d({pwm_start_stop[17],pwm_start_stop[17]}),
    .q({\PWM1/pnumr[12]_keep ,\PWM1/pnumr[5]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg2_b13|PWM1/reg3_b13  (
    .a({\PWM1/pnumr [13],_al_u1811_o}),
    .b({pnum1[13],\PWM1/n24 }),
    .c({pnum1[32],pnumcnt1[13]}),
    .clk(clk100m),
    .d({pwm_start_stop[17],\PWM1/pnumr [13]}),
    .e({open_n2287,pwm_start_stop[17]}),
    .q({\PWM1/pnumr[13]_keep ,\PWM1/RemaTxNum[13]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg2_b14|PWM1/reg3_b14  (
    .a({\PWM1/pnumr [14],_al_u1809_o}),
    .b({pnum1[14],\PWM1/n24 }),
    .c({pnum1[32],pnumcnt1[14]}),
    .clk(clk100m),
    .d({pwm_start_stop[17],\PWM1/pnumr [14]}),
    .e({open_n2309,pwm_start_stop[17]}),
    .q({\PWM1/pnumr[14]_keep ,\PWM1/RemaTxNum[14]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg2_b15|PWM1/reg2_b23  (
    .a({\PWM1/pnumr [15],\PWM1/pnumr [23]}),
    .b({pnum1[15],pnum1[23]}),
    .c({pnum1[32],pnum1[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[17],pwm_start_stop[17]}),
    .q({\PWM1/pnumr[15]_keep ,\PWM1/pnumr[23]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg2_b16|PWM1/reg2_b22  (
    .a({\PWM1/pnumr [16],\PWM1/pnumr [22]}),
    .b({pnum1[16],pnum1[22]}),
    .c({pnum1[32],pnum1[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[17],pwm_start_stop[17]}),
    .q({\PWM1/pnumr[16]_keep ,\PWM1/pnumr[22]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg2_b17|PWM1/reg3_b17  (
    .a({\PWM1/pnumr [17],_al_u1803_o}),
    .b({pnum1[17],\PWM1/n24 }),
    .c({pnum1[32],pnumcnt1[17]}),
    .clk(clk100m),
    .d({pwm_start_stop[17],\PWM1/pnumr [17]}),
    .e({open_n2373,pwm_start_stop[17]}),
    .q({\PWM1/pnumr[17]_keep ,\PWM1/RemaTxNum[17]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg2_b18|PWM1/reg3_b18  (
    .a({\PWM1/pnumr [18],_al_u1801_o}),
    .b({pnum1[18],\PWM1/n24 }),
    .c({pnum1[32],pnumcnt1[18]}),
    .clk(clk100m),
    .d({pwm_start_stop[17],\PWM1/pnumr [18]}),
    .e({open_n2395,pwm_start_stop[17]}),
    .q({\PWM1/pnumr[18]_keep ,\PWM1/RemaTxNum[18]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg2_b19|PWM1/reg2_b2  (
    .a({\PWM1/pnumr [19],\PWM1/pnumr [2]}),
    .b({pnum1[19],pnum1[2]}),
    .c({pnum1[32],pnum1[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[17],pwm_start_stop[17]}),
    .q({\PWM1/pnumr[19]_keep ,\PWM1/pnumr[2]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg2_b1|PWM1/reg3_b1  (
    .a({\PWM1/pnumr [1],_al_u1819_o}),
    .b({pnum1[1],\PWM1/n24 }),
    .c({pnum1[32],pnumcnt1[1]}),
    .clk(clk100m),
    .d({pwm_start_stop[17],\PWM1/pnumr [1]}),
    .e({open_n2436,pwm_start_stop[17]}),
    .q({\PWM1/pnumr[1]_keep ,\PWM1/RemaTxNum[1]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg2_b20|PWM1/reg3_b20  (
    .a({\PWM1/pnumr [20],_al_u1795_o}),
    .b({pnum1[20],\PWM1/n24 }),
    .c({pnum1[32],pnumcnt1[20]}),
    .clk(clk100m),
    .d({pwm_start_stop[17],\PWM1/pnumr [20]}),
    .e({open_n2458,pwm_start_stop[17]}),
    .q({\PWM1/pnumr[20]_keep ,\PWM1/RemaTxNum[20]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg2_b21|PWM1/reg3_b21  (
    .a({\PWM1/pnumr [21],_al_u1793_o}),
    .b({pnum1[21],\PWM1/n24 }),
    .c({pnum1[32],pnumcnt1[21]}),
    .clk(clk100m),
    .d({pwm_start_stop[17],\PWM1/pnumr [21]}),
    .e({open_n2480,pwm_start_stop[17]}),
    .q({\PWM1/pnumr[21]_keep ,\PWM1/RemaTxNum[21]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg2_b24|PWM1/reg2_b31  (
    .a({\PWM1/pnumr [24],\PWM1/pnumr [31]}),
    .b({pnum1[24],pnum1[31]}),
    .c({pnum1[32],pnum1[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[17],pwm_start_stop[17]}),
    .q({\PWM1/pnumr[24]_keep ,\PWM1/pnumr[31]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg2_b25|PWM1/reg2_b30  (
    .a({\PWM1/pnumr [25],\PWM1/pnumr [30]}),
    .b({pnum1[25],pnum1[30]}),
    .c({pnum1[32],pnum1[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[17],pwm_start_stop[17]}),
    .q({\PWM1/pnumr[25]_keep ,\PWM1/pnumr[30]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg2_b26|PWM1/reg2_b29  (
    .a({\PWM1/pnumr [26],\PWM1/pnumr [29]}),
    .b({pnum1[26],pnum1[29]}),
    .c({pnum1[32],pnum1[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[17],pwm_start_stop[17]}),
    .q({\PWM1/pnumr[26]_keep ,\PWM1/pnumr[29]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg2_b27|PWM1/reg2_b28  (
    .a({\PWM1/pnumr [27],\PWM1/pnumr [28]}),
    .b({pnum1[27],pnum1[28]}),
    .c({pnum1[32],pnum1[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[17],pwm_start_stop[17]}),
    .q({\PWM1/pnumr[27]_keep ,\PWM1/pnumr[28]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg2_b3|PWM1/reg3_b3  (
    .a({\PWM1/pnumr [3],_al_u1787_o}),
    .b({pnum1[3],\PWM1/n24 }),
    .c({pnum1[32],pnumcnt1[3]}),
    .clk(clk100m),
    .d({pwm_start_stop[17],\PWM1/pnumr [3]}),
    .e({open_n2590,pwm_start_stop[17]}),
    .q({\PWM1/pnumr[3]_keep ,\PWM1/RemaTxNum[3]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg2_b4|PWM1/reg3_b4  (
    .a({\PWM1/pnumr [4],_al_u1785_o}),
    .b({pnum1[32],\PWM1/n24 }),
    .c({pnum1[4],pnumcnt1[4]}),
    .clk(clk100m),
    .d({pwm_start_stop[17],\PWM1/pnumr [4]}),
    .e({open_n2612,pwm_start_stop[17]}),
    .q({\PWM1/pnumr[4]_keep ,\PWM1/RemaTxNum[4]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg2_b7|PWM1/reg3_b7  (
    .a({\PWM1/pnumr [7],_al_u1779_o}),
    .b({pnum1[32],\PWM1/n24 }),
    .c({pnum1[7],pnumcnt1[7]}),
    .clk(clk100m),
    .d({pwm_start_stop[17],\PWM1/pnumr [7]}),
    .e({open_n2634,pwm_start_stop[17]}),
    .q({\PWM1/pnumr[7]_keep ,\PWM1/RemaTxNum[7]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg2_b8|PWM1/reg3_b8  (
    .a({\PWM1/pnumr [8],_al_u1777_o}),
    .b({pnum1[32],\PWM1/n24 }),
    .c({pnum1[8],pnumcnt1[8]}),
    .clk(clk100m),
    .d({pwm_start_stop[17],\PWM1/pnumr [8]}),
    .e({open_n2656,pwm_start_stop[17]}),
    .q({\PWM1/pnumr[8]_keep ,\PWM1/RemaTxNum[8]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg3_b0  (
    .a({_al_u1821_o,_al_u1821_o}),
    .b({\PWM1/n24 ,\PWM1/n24 }),
    .c({pnumcnt1[0],pnumcnt1[0]}),
    .clk(clk100m),
    .d({\PWM1/pnumr [0],\PWM1/pnumr [0]}),
    .mi({open_n2688,pwm_start_stop[17]}),
    .q({open_n2695,\PWM1/RemaTxNum[0]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg3_b11  (
    .a({_al_u1815_o,_al_u1815_o}),
    .b({\PWM1/n24 ,\PWM1/n24 }),
    .c({pnumcnt1[11],pnumcnt1[11]}),
    .clk(clk100m),
    .d({\PWM1/pnumr [11],\PWM1/pnumr [11]}),
    .mi({open_n2707,pwm_start_stop[17]}),
    .q({open_n2714,\PWM1/RemaTxNum[11]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg3_b12  (
    .a({_al_u1813_o,_al_u1813_o}),
    .b({\PWM1/n24 ,\PWM1/n24 }),
    .c({pnumcnt1[12],pnumcnt1[12]}),
    .clk(clk100m),
    .d({\PWM1/pnumr [12],\PWM1/pnumr [12]}),
    .mi({open_n2726,pwm_start_stop[17]}),
    .q({open_n2733,\PWM1/RemaTxNum[12]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg3_b15  (
    .a({_al_u1807_o,_al_u1807_o}),
    .b({\PWM1/n24 ,\PWM1/n24 }),
    .c({pnumcnt1[15],pnumcnt1[15]}),
    .clk(clk100m),
    .d({\PWM1/pnumr [15],\PWM1/pnumr [15]}),
    .mi({open_n2745,pwm_start_stop[17]}),
    .q({open_n2752,\PWM1/RemaTxNum[15]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg3_b16  (
    .a({_al_u1805_o,_al_u1805_o}),
    .b({\PWM1/n24 ,\PWM1/n24 }),
    .c({pnumcnt1[16],pnumcnt1[16]}),
    .clk(clk100m),
    .d({\PWM1/pnumr [16],\PWM1/pnumr [16]}),
    .mi({open_n2764,pwm_start_stop[17]}),
    .q({open_n2771,\PWM1/RemaTxNum[16]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg3_b19  (
    .a({_al_u1799_o,_al_u1799_o}),
    .b({\PWM1/n24 ,\PWM1/n24 }),
    .c({pnumcnt1[19],pnumcnt1[19]}),
    .clk(clk100m),
    .d({\PWM1/pnumr [19],\PWM1/pnumr [19]}),
    .mi({open_n2783,pwm_start_stop[17]}),
    .q({open_n2790,\PWM1/RemaTxNum[19]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg3_b2  (
    .a({_al_u1797_o,_al_u1797_o}),
    .b({\PWM1/n24 ,\PWM1/n24 }),
    .c({pnumcnt1[2],pnumcnt1[2]}),
    .clk(clk100m),
    .d({\PWM1/pnumr [2],\PWM1/pnumr [2]}),
    .mi({open_n2802,pwm_start_stop[17]}),
    .q({open_n2809,\PWM1/RemaTxNum[2]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg3_b22  (
    .a({_al_u1791_o,_al_u1791_o}),
    .b({\PWM1/n24 ,\PWM1/n24 }),
    .c({pnumcnt1[22],pnumcnt1[22]}),
    .clk(clk100m),
    .d({\PWM1/pnumr [22],\PWM1/pnumr [22]}),
    .mi({open_n2821,pwm_start_stop[17]}),
    .q({open_n2828,\PWM1/RemaTxNum[22]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg3_b23  (
    .a({_al_u1789_o,_al_u1789_o}),
    .b({\PWM1/n24 ,\PWM1/n24 }),
    .c({pnumcnt1[23],pnumcnt1[23]}),
    .clk(clk100m),
    .d({\PWM1/pnumr [23],\PWM1/pnumr [23]}),
    .mi({open_n2840,pwm_start_stop[17]}),
    .q({open_n2847,\PWM1/RemaTxNum[23]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg3_b5  (
    .a({_al_u1783_o,_al_u1783_o}),
    .b({\PWM1/n24 ,\PWM1/n24 }),
    .c({pnumcnt1[5],pnumcnt1[5]}),
    .clk(clk100m),
    .d({\PWM1/pnumr [5],\PWM1/pnumr [5]}),
    .mi({open_n2859,pwm_start_stop[17]}),
    .q({open_n2866,\PWM1/RemaTxNum[5]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg3_b6  (
    .a({_al_u1781_o,_al_u1781_o}),
    .b({\PWM1/n24 ,\PWM1/n24 }),
    .c({pnumcnt1[6],pnumcnt1[6]}),
    .clk(clk100m),
    .d({\PWM1/pnumr [6],\PWM1/pnumr [6]}),
    .mi({open_n2878,pwm_start_stop[17]}),
    .q({open_n2885,\PWM1/RemaTxNum[6]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/reg3_b9  (
    .a({_al_u1775_o,_al_u1775_o}),
    .b({\PWM1/n24 ,\PWM1/n24 }),
    .c({pnumcnt1[9],pnumcnt1[9]}),
    .clk(clk100m),
    .d({\PWM1/pnumr [9],\PWM1/pnumr [9]}),
    .mi({open_n2897,pwm_start_stop[17]}),
    .q({open_n2904,\PWM1/RemaTxNum[9]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_LSLICE #(
    //.MACRO("PWM1/sub0/ucin_al_u3370"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM1/sub0/u11_al_u3373  (
    .a({\PWM1/FreCnt [13],\PWM1/FreCnt [11]}),
    .b({\PWM1/FreCnt [14],\PWM1/FreCnt [12]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM1/sub0/c11 ),
    .f({\PWM1/n12 [13],\PWM1/n12 [11]}),
    .fco(\PWM1/sub0/c15 ),
    .fx({\PWM1/n12 [14],\PWM1/n12 [12]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM1/sub0/ucin_al_u3370"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM1/sub0/u15_al_u3374  (
    .a({\PWM1/FreCnt [17],\PWM1/FreCnt [15]}),
    .b({\PWM1/FreCnt [18],\PWM1/FreCnt [16]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM1/sub0/c15 ),
    .f({\PWM1/n12 [17],\PWM1/n12 [15]}),
    .fco(\PWM1/sub0/c19 ),
    .fx({\PWM1/n12 [18],\PWM1/n12 [16]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM1/sub0/ucin_al_u3370"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM1/sub0/u19_al_u3375  (
    .a({\PWM1/FreCnt [21],\PWM1/FreCnt [19]}),
    .b({\PWM1/FreCnt [22],\PWM1/FreCnt [20]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM1/sub0/c19 ),
    .f({\PWM1/n12 [21],\PWM1/n12 [19]}),
    .fco(\PWM1/sub0/c23 ),
    .fx({\PWM1/n12 [22],\PWM1/n12 [20]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM1/sub0/ucin_al_u3370"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM1/sub0/u23_al_u3376  (
    .a({\PWM1/FreCnt [25],\PWM1/FreCnt [23]}),
    .b({\PWM1/FreCnt [26],\PWM1/FreCnt [24]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM1/sub0/c23 ),
    .f({\PWM1/n12 [25],\PWM1/n12 [23]}),
    .fx({\PWM1/n12 [26],\PWM1/n12 [24]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM1/sub0/ucin_al_u3370"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM1/sub0/u3_al_u3371  (
    .a({\PWM1/FreCnt [5],\PWM1/FreCnt [3]}),
    .b({\PWM1/FreCnt [6],\PWM1/FreCnt [4]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM1/sub0/c3 ),
    .f({\PWM1/n12 [5],\PWM1/n12 [3]}),
    .fco(\PWM1/sub0/c7 ),
    .fx({\PWM1/n12 [6],\PWM1/n12 [4]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM1/sub0/ucin_al_u3370"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM1/sub0/u7_al_u3372  (
    .a({\PWM1/FreCnt [9],\PWM1/FreCnt [7]}),
    .b({\PWM1/FreCnt [10],\PWM1/FreCnt [8]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM1/sub0/c7 ),
    .f({\PWM1/n12 [9],\PWM1/n12 [7]}),
    .fco(\PWM1/sub0/c11 ),
    .fx({\PWM1/n12 [10],\PWM1/n12 [8]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM1/sub0/ucin_al_u3370"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h0005),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM1/sub0/ucin_al_u3370  (
    .a({\PWM1/FreCnt [1],1'b0}),
    .b({\PWM1/FreCnt [2],\PWM1/FreCnt [0]}),
    .c(2'b11),
    .d(2'b01),
    .e(2'b01),
    .f({\PWM1/n12 [1],open_n3031}),
    .fco(\PWM1/sub0/c3 ),
    .fx({\PWM1/n12 [2],\PWM1/n12 [0]}));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM1/sub1/u0|PWM1/sub1/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("SUB_CARRY"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000101),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM1/sub1/u0|PWM1/sub1/ucin  (
    .a({pnumcnt1[0],1'b0}),
    .b({1'b1,open_n3034}),
    .ce(\U_AHB/n10 ),
    .clk(clk100m),
    .mi({\U_AHB/h2h_hwdata [9],\U_AHB/h2h_hwdata [6]}),
    .f({\PWM1/n26 [0],open_n3050}),
    .fco(\PWM1/sub1/c1 ),
    .q({freq3[9],freq3[6]}));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM1/sub1/u0|PWM1/sub1/ucin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM1/sub1/u10|PWM1/sub1/u9  (
    .a(pnumcnt1[10:9]),
    .b(2'b00),
    .fci(\PWM1/sub1/c9 ),
    .f(\PWM1/n26 [10:9]),
    .fco(\PWM1/sub1/c11 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM1/sub1/u0|PWM1/sub1/ucin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM1/sub1/u12|PWM1/sub1/u11  (
    .a(pnumcnt1[12:11]),
    .b(2'b00),
    .fci(\PWM1/sub1/c11 ),
    .f(\PWM1/n26 [12:11]),
    .fco(\PWM1/sub1/c13 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM1/sub1/u0|PWM1/sub1/ucin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM1/sub1/u14|PWM1/sub1/u13  (
    .a(pnumcnt1[14:13]),
    .b(2'b00),
    .fci(\PWM1/sub1/c13 ),
    .f(\PWM1/n26 [14:13]),
    .fco(\PWM1/sub1/c15 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM1/sub1/u0|PWM1/sub1/ucin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM1/sub1/u16|PWM1/sub1/u15  (
    .a(pnumcnt1[16:15]),
    .b(2'b00),
    .fci(\PWM1/sub1/c15 ),
    .f(\PWM1/n26 [16:15]),
    .fco(\PWM1/sub1/c17 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM1/sub1/u0|PWM1/sub1/ucin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM1/sub1/u18|PWM1/sub1/u17  (
    .a(pnumcnt1[18:17]),
    .b(2'b00),
    .fci(\PWM1/sub1/c17 ),
    .f(\PWM1/n26 [18:17]),
    .fco(\PWM1/sub1/c19 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM1/sub1/u0|PWM1/sub1/ucin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM1/sub1/u20|PWM1/sub1/u19  (
    .a(pnumcnt1[20:19]),
    .b(2'b00),
    .fci(\PWM1/sub1/c19 ),
    .f(\PWM1/n26 [20:19]),
    .fco(\PWM1/sub1/c21 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM1/sub1/u0|PWM1/sub1/ucin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM1/sub1/u22|PWM1/sub1/u21  (
    .a(pnumcnt1[22:21]),
    .b(2'b00),
    .fci(\PWM1/sub1/c21 ),
    .f(\PWM1/n26 [22:21]),
    .fco(\PWM1/sub1/c23 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM1/sub1/u0|PWM1/sub1/ucin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM1/sub1/u23_al_u3469  (
    .a({open_n3207,pnumcnt1[23]}),
    .b({open_n3208,1'b0}),
    .fci(\PWM1/sub1/c23 ),
    .f({open_n3227,\PWM1/n26 [23]}));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM1/sub1/u0|PWM1/sub1/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM1/sub1/u2|PWM1/sub1/u1  (
    .a(pnumcnt1[2:1]),
    .b(2'b00),
    .fci(\PWM1/sub1/c1 ),
    .f(\PWM1/n26 [2:1]),
    .fco(\PWM1/sub1/c3 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM1/sub1/u0|PWM1/sub1/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM1/sub1/u4|PWM1/sub1/u3  (
    .a(pnumcnt1[4:3]),
    .b(2'b00),
    .fci(\PWM1/sub1/c3 ),
    .f(\PWM1/n26 [4:3]),
    .fco(\PWM1/sub1/c5 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM1/sub1/u0|PWM1/sub1/ucin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM1/sub1/u6|PWM1/sub1/u5  (
    .a(pnumcnt1[6:5]),
    .b(2'b00),
    .fci(\PWM1/sub1/c5 ),
    .f(\PWM1/n26 [6:5]),
    .fco(\PWM1/sub1/c7 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM1/sub1/u0|PWM1/sub1/ucin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM1/sub1/u8|PWM1/sub1/u7  (
    .a(pnumcnt1[8:7]),
    .b(2'b00),
    .fci(\PWM1/sub1/c7 ),
    .f(\PWM1/n26 [8:7]),
    .fco(\PWM1/sub1/c9 ));
  // src/OnePWM.v(26)
  // src/OnePWM.v(26)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*~(~D*B*~A))"),
    //.LUT1("(C*~(~D*B*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000010110000),
    .INIT_LUT1(16'b1111000010110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \PWM2/State_reg|PWMD/State_reg  (
    .a({_al_u3013_o,_al_u3046_o}),
    .b({\PWM2/n0_lutinv ,\PWMD/n0_lutinv }),
    .c({_al_u3014_o,_al_u3047_o}),
    .clk(clk100m),
    .d({pwm_start_stop[18],pwm_start_stop[29]}),
    .sr(rstn),
    .q({pwm_state_read[2],pwm_state_read[13]}));  // src/OnePWM.v(26)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[0]  (
    .i(\PWM2/RemaTxNum[0]_keep ),
    .o(pnumcnt2[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[10]  (
    .i(\PWM2/RemaTxNum[10]_keep ),
    .o(pnumcnt2[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[11]  (
    .i(\PWM2/RemaTxNum[11]_keep ),
    .o(pnumcnt2[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[12]  (
    .i(\PWM2/RemaTxNum[12]_keep ),
    .o(pnumcnt2[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[13]  (
    .i(\PWM2/RemaTxNum[13]_keep ),
    .o(pnumcnt2[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[14]  (
    .i(\PWM2/RemaTxNum[14]_keep ),
    .o(pnumcnt2[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[15]  (
    .i(\PWM2/RemaTxNum[15]_keep ),
    .o(pnumcnt2[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[16]  (
    .i(\PWM2/RemaTxNum[16]_keep ),
    .o(pnumcnt2[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[17]  (
    .i(\PWM2/RemaTxNum[17]_keep ),
    .o(pnumcnt2[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[18]  (
    .i(\PWM2/RemaTxNum[18]_keep ),
    .o(pnumcnt2[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[19]  (
    .i(\PWM2/RemaTxNum[19]_keep ),
    .o(pnumcnt2[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[1]  (
    .i(\PWM2/RemaTxNum[1]_keep ),
    .o(pnumcnt2[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[20]  (
    .i(\PWM2/RemaTxNum[20]_keep ),
    .o(pnumcnt2[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[21]  (
    .i(\PWM2/RemaTxNum[21]_keep ),
    .o(pnumcnt2[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[22]  (
    .i(\PWM2/RemaTxNum[22]_keep ),
    .o(pnumcnt2[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[23]  (
    .i(\PWM2/RemaTxNum[23]_keep ),
    .o(pnumcnt2[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[2]  (
    .i(\PWM2/RemaTxNum[2]_keep ),
    .o(pnumcnt2[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[3]  (
    .i(\PWM2/RemaTxNum[3]_keep ),
    .o(pnumcnt2[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[4]  (
    .i(\PWM2/RemaTxNum[4]_keep ),
    .o(pnumcnt2[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[5]  (
    .i(\PWM2/RemaTxNum[5]_keep ),
    .o(pnumcnt2[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[6]  (
    .i(\PWM2/RemaTxNum[6]_keep ),
    .o(pnumcnt2[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[7]  (
    .i(\PWM2/RemaTxNum[7]_keep ),
    .o(pnumcnt2[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[8]  (
    .i(\PWM2/RemaTxNum[8]_keep ),
    .o(pnumcnt2[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[9]  (
    .i(\PWM2/RemaTxNum[9]_keep ),
    .o(pnumcnt2[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_dir  (
    .i(\PWM2/dir_keep ),
    .o(dir_pad[2]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[0]  (
    .i(\PWM2/pnumr[0]_keep ),
    .o(\PWM2/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[10]  (
    .i(\PWM2/pnumr[10]_keep ),
    .o(\PWM2/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[11]  (
    .i(\PWM2/pnumr[11]_keep ),
    .o(\PWM2/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[12]  (
    .i(\PWM2/pnumr[12]_keep ),
    .o(\PWM2/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[13]  (
    .i(\PWM2/pnumr[13]_keep ),
    .o(\PWM2/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[14]  (
    .i(\PWM2/pnumr[14]_keep ),
    .o(\PWM2/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[15]  (
    .i(\PWM2/pnumr[15]_keep ),
    .o(\PWM2/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[16]  (
    .i(\PWM2/pnumr[16]_keep ),
    .o(\PWM2/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[17]  (
    .i(\PWM2/pnumr[17]_keep ),
    .o(\PWM2/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[18]  (
    .i(\PWM2/pnumr[18]_keep ),
    .o(\PWM2/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[19]  (
    .i(\PWM2/pnumr[19]_keep ),
    .o(\PWM2/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[1]  (
    .i(\PWM2/pnumr[1]_keep ),
    .o(\PWM2/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[20]  (
    .i(\PWM2/pnumr[20]_keep ),
    .o(\PWM2/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[21]  (
    .i(\PWM2/pnumr[21]_keep ),
    .o(\PWM2/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[22]  (
    .i(\PWM2/pnumr[22]_keep ),
    .o(\PWM2/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[23]  (
    .i(\PWM2/pnumr[23]_keep ),
    .o(\PWM2/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[24]  (
    .i(\PWM2/pnumr[24]_keep ),
    .o(\PWM2/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[25]  (
    .i(\PWM2/pnumr[25]_keep ),
    .o(\PWM2/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[26]  (
    .i(\PWM2/pnumr[26]_keep ),
    .o(\PWM2/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[27]  (
    .i(\PWM2/pnumr[27]_keep ),
    .o(\PWM2/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[28]  (
    .i(\PWM2/pnumr[28]_keep ),
    .o(\PWM2/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[29]  (
    .i(\PWM2/pnumr[29]_keep ),
    .o(\PWM2/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[2]  (
    .i(\PWM2/pnumr[2]_keep ),
    .o(\PWM2/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[30]  (
    .i(\PWM2/pnumr[30]_keep ),
    .o(\PWM2/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[31]  (
    .i(\PWM2/pnumr[31]_keep ),
    .o(\PWM2/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[3]  (
    .i(\PWM2/pnumr[3]_keep ),
    .o(\PWM2/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[4]  (
    .i(\PWM2/pnumr[4]_keep ),
    .o(\PWM2/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[5]  (
    .i(\PWM2/pnumr[5]_keep ),
    .o(\PWM2/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[6]  (
    .i(\PWM2/pnumr[6]_keep ),
    .o(\PWM2/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[7]  (
    .i(\PWM2/pnumr[7]_keep ),
    .o(\PWM2/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[8]  (
    .i(\PWM2/pnumr[8]_keep ),
    .o(\PWM2/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[9]  (
    .i(\PWM2/pnumr[9]_keep ),
    .o(\PWM2/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pwm  (
    .i(\PWM2/pwm_keep ),
    .o(pwm_pad[2]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_stopreq  (
    .i(\PWM2/stopreq_keep ),
    .o(\PWM2/stopreq ));  // src/OnePWM.v(14)
  EF2_PHY_MSLICE #(
    //.LUT0("~(~0*~(D*C*B*A))"),
    //.LUT1("~(~1*~(D*C*B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b1111111111111111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM2/pwm_reg  (
    .a({_al_u1400_o,_al_u1400_o}),
    .b({_al_u1407_o,_al_u1407_o}),
    .c({_al_u1409_o,_al_u1409_o}),
    .clk(clk100m),
    .d({_al_u1411_o,_al_u1411_o}),
    .mi({open_n3350,pwm_pad[2]}),
    .sr(\PWM2/u14_sel_is_1_o ),
    .q({open_n3356,\PWM2/pwm_keep }));  // src/OnePWM.v(45)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM2/reg0_b0|PWM2/reg0_b15  (
    .b({\PWM2/n12 [0],\PWM2/n12 [15]}),
    .c({freq2[0],freq2[15]}),
    .clk(clk100m),
    .d({\PWM2/n0_lutinv ,\PWM2/n0_lutinv }),
    .sr(\PWM2/n11 ),
    .q({\PWM2/FreCnt [0],\PWM2/FreCnt [15]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM2/reg0_b10|PWM2/reg0_b1  (
    .b({\PWM2/n12 [10],\PWM2/n12 [1]}),
    .c({freq2[10],freq2[1]}),
    .clk(clk100m),
    .d({\PWM2/n0_lutinv ,\PWM2/n0_lutinv }),
    .sr(\PWM2/n11 ),
    .q({\PWM2/FreCnt [10],\PWM2/FreCnt [1]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM2/reg0_b11|PWM2/reg0_b8  (
    .b({\PWM2/n12 [11],\PWM2/n12 [8]}),
    .c({freq2[11],freq2[8]}),
    .clk(clk100m),
    .d({\PWM2/n0_lutinv ,\PWM2/n0_lutinv }),
    .sr(\PWM2/n11 ),
    .q({\PWM2/FreCnt [11],\PWM2/FreCnt [8]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM2/reg0_b12|PWM2/reg0_b7  (
    .b({\PWM2/n12 [12],\PWM2/n12 [7]}),
    .c({freq2[12],freq2[7]}),
    .clk(clk100m),
    .d({\PWM2/n0_lutinv ,\PWM2/n0_lutinv }),
    .sr(\PWM2/n11 ),
    .q({\PWM2/FreCnt [12],\PWM2/FreCnt [7]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM2/reg0_b13|PWM2/reg0_b5  (
    .b({\PWM2/n12 [13],\PWM2/n12 [5]}),
    .c({freq2[13],freq2[5]}),
    .clk(clk100m),
    .d({\PWM2/n0_lutinv ,\PWM2/n0_lutinv }),
    .sr(\PWM2/n11 ),
    .q({\PWM2/FreCnt [13],\PWM2/FreCnt [5]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM2/reg0_b14|PWM2/reg0_b3  (
    .b({\PWM2/n12 [14],\PWM2/n12 [3]}),
    .c({freq2[14],freq2[3]}),
    .clk(clk100m),
    .d({\PWM2/n0_lutinv ,\PWM2/n0_lutinv }),
    .sr(\PWM2/n11 ),
    .q({\PWM2/FreCnt [14],\PWM2/FreCnt [3]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM2/reg0_b16|PWM2/reg0_b25  (
    .b({\PWM2/n12 [16],\PWM2/n12 [25]}),
    .c({freq2[16],freq2[25]}),
    .clk(clk100m),
    .d({\PWM2/n0_lutinv ,\PWM2/n0_lutinv }),
    .sr(\PWM2/n11 ),
    .q({\PWM2/FreCnt [16],\PWM2/FreCnt [25]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM2/reg0_b17|PWM2/reg0_b23  (
    .b({\PWM2/n12 [17],\PWM2/n12 [23]}),
    .c({freq2[17],freq2[23]}),
    .clk(clk100m),
    .d({\PWM2/n0_lutinv ,\PWM2/n0_lutinv }),
    .sr(\PWM2/n11 ),
    .q({\PWM2/FreCnt [17],\PWM2/FreCnt [23]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM2/reg0_b18|PWM2/reg0_b21  (
    .b({\PWM2/n12 [18],\PWM2/n12 [21]}),
    .c({freq2[18],freq2[21]}),
    .clk(clk100m),
    .d({\PWM2/n0_lutinv ,\PWM2/n0_lutinv }),
    .sr(\PWM2/n11 ),
    .q({\PWM2/FreCnt [18],\PWM2/FreCnt [21]}));  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM2/reg0_b2  (
    .b({open_n3551,\PWM2/n12 [2]}),
    .c({open_n3552,freq2[2]}),
    .clk(clk100m),
    .d({open_n3554,\PWM2/n0_lutinv }),
    .sr(\PWM2/n11 ),
    .q({open_n3572,\PWM2/FreCnt [2]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM2/reg0_b20|PWM2/reg0_b19  (
    .b(\PWM2/n12 [20:19]),
    .c(freq2[20:19]),
    .clk(clk100m),
    .d({\PWM2/n0_lutinv ,\PWM2/n0_lutinv }),
    .sr(\PWM2/n11 ),
    .q(\PWM2/FreCnt [20:19]));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM2/reg0_b22|PWM2/reg0_b9  (
    .b({\PWM2/n12 [22],\PWM2/n12 [9]}),
    .c({freq2[22],freq2[9]}),
    .clk(clk100m),
    .d({\PWM2/n0_lutinv ,\PWM2/n0_lutinv }),
    .sr(\PWM2/n11 ),
    .q({\PWM2/FreCnt [22],\PWM2/FreCnt [9]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM2/reg0_b24|PWM2/reg0_b6  (
    .b({\PWM2/n12 [24],\PWM2/n12 [6]}),
    .c({freq2[24],freq2[6]}),
    .clk(clk100m),
    .d({\PWM2/n0_lutinv ,\PWM2/n0_lutinv }),
    .sr(\PWM2/n11 ),
    .q({\PWM2/FreCnt [24],\PWM2/FreCnt [6]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM2/reg0_b26|PWM2/reg0_b4  (
    .b({\PWM2/n12 [26],\PWM2/n12 [4]}),
    .c({freq2[26],freq2[4]}),
    .clk(clk100m),
    .d({\PWM2/n0_lutinv ,\PWM2/n0_lutinv }),
    .sr(\PWM2/n11 ),
    .q({\PWM2/FreCnt [26],\PWM2/FreCnt [4]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*~C)*~(D*~B))"),
    //.LUTF1("(A*~(~0*C)*~(D*~B))"),
    //.LUTG0("(A*~(1*~C)*~(D*~B))"),
    //.LUTG1("(A*~(~1*C)*~(D*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000100010101010),
    .INIT_LUTF1(16'b0000100000001010),
    .INIT_LUTG0(16'b1000000010100000),
    .INIT_LUTG1(16'b1000100010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg1_b11|PWM2/reg1_b26  (
    .a({_al_u1909_o,_al_u1905_o}),
    .b({\PWM2/FreCnt [10],\PWM2/FreCnt [17]}),
    .c({\PWM2/FreCnt [25],\PWM2/FreCnt [25]}),
    .ce(\PWM2/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM2/FreCntr [11],\PWM2/FreCntr [18]}),
    .e({\PWM2/FreCntr [26],\PWM2/FreCntr [26]}),
    .mi({freq2[11],freq2[26]}),
    .f({_al_u1910_o,_al_u1906_o}),
    .q({\PWM2/FreCntr [11],\PWM2/FreCntr [26]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D@C)*~(0@B))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(A*~(D@C)*~(1@B))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010000000000010),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000000000001000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg1_b14|PWM2/reg1_b10  (
    .a({\PWM2/FreCnt [14],_al_u1914_o}),
    .b({\PWM2/FreCnt [25],\PWM2/FreCnt [13]}),
    .c({\PWM2/FreCntr [14],\PWM2/FreCnt [9]}),
    .ce(\PWM2/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM2/FreCntr [25],\PWM2/FreCntr [10]}),
    .e({open_n3681,\PWM2/FreCntr [14]}),
    .mi({freq2[14],freq2[10]}),
    .f({_al_u1408_o,_al_u1915_o}),
    .q({\PWM2/FreCntr [14],\PWM2/FreCntr [10]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~D*B)*~(~C*A))"),
    //.LUTF1("(~(~D*B)*~(~C*A))"),
    //.LUTG0("(~(~D*B)*~(~C*A))"),
    //.LUTG1("(~(~D*B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111010100110001),
    .INIT_LUTF1(16'b1111010100110001),
    .INIT_LUTG0(16'b1111010100110001),
    .INIT_LUTG1(16'b1111010100110001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg1_b18|PWM2/reg1_b2  (
    .a({\PWM2/FreCnt [17],\PWM2/FreCnt [1]}),
    .b({\PWM2/FreCnt [3],\PWM2/FreCnt [23]}),
    .c({\PWM2/FreCntr [18],\PWM2/FreCntr [2]}),
    .ce(\PWM2/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM2/FreCntr [4],\PWM2/FreCntr [24]}),
    .mi({freq2[18],freq2[2]}),
    .f({_al_u1924_o,_al_u1916_o}),
    .q({\PWM2/FreCntr [18],\PWM2/FreCntr [2]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg1_b1|PWM2/reg1_b19  (
    .a({\PWM2/FreCnt [0],_al_u1410_o}),
    .b({\PWM2/FreCnt [18],\PWM2/FreCnt [19]}),
    .c({\PWM2/FreCntr [1],\PWM2/FreCnt [2]}),
    .ce(\PWM2/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM2/FreCntr [19],\PWM2/FreCntr [19]}),
    .e({open_n3716,\PWM2/FreCntr [2]}),
    .mi({freq2[1],freq2[19]}),
    .f({_al_u1920_o,_al_u1411_o}),
    .q({\PWM2/FreCntr [1],\PWM2/FreCntr [19]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~A*~(0@C)*~(~D*B))"),
    //.LUTF1("(~A*~(0*~C)*~(D@B))"),
    //.LUTG0("(~A*~(1@C)*~(~D*B))"),
    //.LUTG1("(~A*~(1*~C)*~(D@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010100000001),
    .INIT_LUTF1(16'b0100010000010001),
    .INIT_LUTG0(16'b0101000000010000),
    .INIT_LUTG1(16'b0100000000010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg1_b21|PWM2/reg1_b24  (
    .a({_al_u1913_o,_al_u1404_o}),
    .b({\PWM2/FreCnt [20],\PWM2/FreCnt [12]}),
    .c({\PWM2/FreCnt [23],\PWM2/FreCnt [24]}),
    .ce(\PWM2/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM2/FreCntr [21],\PWM2/FreCntr [12]}),
    .e({\PWM2/FreCntr [24],\PWM2/FreCntr [24]}),
    .mi({freq2[21],freq2[24]}),
    .f({_al_u1914_o,_al_u1405_o}),
    .q({\PWM2/FreCntr [21],\PWM2/FreCntr [24]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*~C)*~(~D*B))"),
    //.LUTF1("(~(D*~B)*~(~C*A))"),
    //.LUTG0("(A*~(1*~C)*~(~D*B))"),
    //.LUTG1("(~(D*~B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101000100010),
    .INIT_LUTF1(16'b1100010011110101),
    .INIT_LUTG0(16'b1010000000100000),
    .INIT_LUTG1(16'b1100010011110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg1_b22|PWM2/reg1_b16  (
    .a({\PWM2/FreCnt [21],_al_u1916_o}),
    .b({\PWM2/FreCnt [5],\PWM2/FreCnt [15]}),
    .c({\PWM2/FreCntr [22],\PWM2/FreCnt [21]}),
    .ce(\PWM2/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM2/FreCntr [6],\PWM2/FreCntr [16]}),
    .e({open_n3749,\PWM2/FreCntr [22]}),
    .mi({freq2[22],freq2[16]}),
    .f({_al_u1907_o,_al_u1917_o}),
    .q({\PWM2/FreCntr [22],\PWM2/FreCntr [16]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~C*~(0@B)*~(~D*A))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(~C*~(1@B)*~(~D*A))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001100000001),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b0000110000000100),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg1_b23|PWM2/reg1_b12  (
    .a({\PWM2/FreCnt [22],\PWM2/FreCnt [11]}),
    .b(\PWM2/FreCnt [23:22]),
    .c({\PWM2/FreCntr [22],\PWM2/FreCnt [26]}),
    .ce(\PWM2/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM2/FreCntr [23],\PWM2/FreCntr [12]}),
    .e({open_n3766,\PWM2/FreCntr [23]}),
    .mi({freq2[23],freq2[12]}),
    .f({_al_u1395_o,_al_u1926_o}),
    .q({\PWM2/FreCntr [23],\PWM2/FreCntr [12]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg1_b3|PWM2/reg1_b15  (
    .a({\PWM2/FreCnt [10],_al_u1922_o}),
    .b({\PWM2/FreCnt [3],\PWM2/FreCnt [14]}),
    .c({\PWM2/FreCntr [10],\PWM2/FreCnt [2]}),
    .ce(\PWM2/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM2/FreCntr [3],\PWM2/FreCntr [15]}),
    .e({open_n3783,\PWM2/FreCntr [3]}),
    .mi({freq2[3],freq2[15]}),
    .f({_al_u1402_o,_al_u1923_o}),
    .q({\PWM2/FreCntr [3],\PWM2/FreCntr [15]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(D@B)*~(C@A))"),
    //.LUTF1("(D*~(C@B))"),
    //.LUTG0("(~(D@B)*~(C@A))"),
    //.LUTG1("(D*~(C@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000010000100001),
    .INIT_LUTF1(16'b1100001100000000),
    .INIT_LUTG0(16'b1000010000100001),
    .INIT_LUTG1(16'b1100001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg1_b5|PWM2/reg1_b25  (
    .a({open_n3800,\PWM2/FreCnt [24]}),
    .b({\PWM2/FreCnt [4],\PWM2/FreCnt [6]}),
    .c({\PWM2/FreCntr [5],\PWM2/FreCntr [25]}),
    .ce(\PWM2/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({_al_u1920_o,\PWM2/FreCntr [7]}),
    .mi({freq2[5],freq2[25]}),
    .f({_al_u1921_o,_al_u1922_o}),
    .q({\PWM2/FreCntr [5],\PWM2/FreCntr [25]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*B*A*~(0@D))"),
    //.LUTF1("(~(~D*B)*~(C*~A))"),
    //.LUTG0("(C*B*A*~(1@D))"),
    //.LUTG1("(~(~D*B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b1010111100100011),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b1010111100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg1_b6|PWM2/reg1_b17  (
    .a({\PWM2/FreCnt [1],_al_u1908_o}),
    .b({\PWM2/FreCnt [5],_al_u1910_o}),
    .c({\PWM2/FreCntr [2],_al_u1911_o}),
    .ce(\PWM2/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM2/FreCntr [6],\PWM2/FreCnt [16]}),
    .e({open_n3819,\PWM2/FreCntr [17]}),
    .mi({freq2[6],freq2[17]}),
    .f({_al_u1911_o,_al_u1912_o}),
    .q({\PWM2/FreCntr [6],\PWM2/FreCntr [17]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~D*B)*~(C*~A))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(~(~D*B)*~(C*~A))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010111100100011),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1010111100100011),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg1_b7|PWM2/reg1_b4  (
    .a({\PWM2/FreCnt [6],\PWM2/FreCnt [3]}),
    .b({\PWM2/FreCnt [7],\PWM2/FreCnt [7]}),
    .c({\PWM2/FreCntr [6],\PWM2/FreCntr [4]}),
    .ce(\PWM2/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM2/FreCntr [7],\PWM2/FreCntr [8]}),
    .mi({freq2[7],freq2[4]}),
    .f({_al_u1397_o,_al_u1909_o}),
    .q({\PWM2/FreCntr [7],\PWM2/FreCntr [4]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*B*A*~(0@D))"),
    //.LUTF1("(~(D*~B)*~(C*~A))"),
    //.LUTG0("(C*B*A*~(1@D))"),
    //.LUTG1("(~(D*~B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b1000110010101111),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b1000110010101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg1_b8|PWM2/reg1_b13  (
    .a({\PWM2/FreCnt [7],_al_u1915_o}),
    .b({\PWM2/FreCnt [8],_al_u1917_o}),
    .c({\PWM2/FreCntr [8],_al_u1918_o}),
    .ce(\PWM2/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM2/FreCntr [9],\PWM2/FreCnt [12]}),
    .e({open_n3854,\PWM2/FreCntr [13]}),
    .mi({freq2[8],freq2[13]}),
    .f({_al_u1918_o,_al_u1919_o}),
    .q({\PWM2/FreCntr [8],\PWM2/FreCntr [13]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(~0*C)*~(D*~B))"),
    //.LUTF1("(~(~D*B)*~(C*~A))"),
    //.LUTG0("(A*~(~1*C)*~(D*~B))"),
    //.LUTG1("(~(~D*B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000001010),
    .INIT_LUTF1(16'b1010111100100011),
    .INIT_LUTG0(16'b1000100010101010),
    .INIT_LUTG1(16'b1010111100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg1_b9|PWM2/reg1_b20  (
    .a({\PWM2/FreCnt [19],_al_u1924_o}),
    .b({\PWM2/FreCnt [8],\PWM2/FreCnt [11]}),
    .c({\PWM2/FreCntr [20],\PWM2/FreCnt [19]}),
    .ce(\PWM2/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM2/FreCntr [9],\PWM2/FreCntr [12]}),
    .e({open_n3871,\PWM2/FreCntr [20]}),
    .mi({freq2[9],freq2[20]}),
    .f({_al_u1905_o,_al_u1925_o}),
    .q({\PWM2/FreCntr [9],\PWM2/FreCntr [20]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011100010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011100010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg2_b0|PWM2/reg2_b7  (
    .a({\PWM2/pnumr [0],\PWM2/pnumr [7]}),
    .b({pnum2[0],pnum2[32]}),
    .c({pnum2[32],pnum2[7]}),
    .clk(clk100m),
    .d({pwm_start_stop[18],pwm_start_stop[18]}),
    .q({\PWM2/pnumr[0]_keep ,\PWM2/pnumr[7]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg2_b10|PWM2/reg3_b10  (
    .a({\PWM2/pnumr [10],_al_u1899_o}),
    .b({pnum2[10],\PWM2/n24 }),
    .c({pnum2[32],pnumcnt2[10]}),
    .clk(clk100m),
    .d({pwm_start_stop[18],\PWM2/pnumr [10]}),
    .e({open_n3912,pwm_start_stop[18]}),
    .q({\PWM2/pnumr[10]_keep ,\PWM2/RemaTxNum[10]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg2_b11|PWM2/reg3_b11  (
    .a({\PWM2/pnumr [11],_al_u1897_o}),
    .b({pnum2[11],\PWM2/n24 }),
    .c({pnum2[32],pnumcnt2[11]}),
    .clk(clk100m),
    .d({pwm_start_stop[18],\PWM2/pnumr [11]}),
    .e({open_n3934,pwm_start_stop[18]}),
    .q({\PWM2/pnumr[11]_keep ,\PWM2/RemaTxNum[11]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011100010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011100010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg2_b12|PWM2/reg2_b6  (
    .a({\PWM2/pnumr [12],\PWM2/pnumr [6]}),
    .b({pnum2[12],pnum2[32]}),
    .c({pnum2[32],pnum2[6]}),
    .clk(clk100m),
    .d({pwm_start_stop[18],pwm_start_stop[18]}),
    .q({\PWM2/pnumr[12]_keep ,\PWM2/pnumr[6]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg2_b13|PWM2/reg2_b3  (
    .a({\PWM2/pnumr [13],\PWM2/pnumr [3]}),
    .b({pnum2[13],pnum2[3]}),
    .c({pnum2[32],pnum2[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[18],pwm_start_stop[18]}),
    .q({\PWM2/pnumr[13]_keep ,\PWM2/pnumr[3]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg2_b14|PWM2/reg3_b14  (
    .a({\PWM2/pnumr [14],_al_u1891_o}),
    .b({pnum2[14],\PWM2/n24 }),
    .c({pnum2[32],pnumcnt2[14]}),
    .clk(clk100m),
    .d({pwm_start_stop[18],\PWM2/pnumr [14]}),
    .e({open_n3998,pwm_start_stop[18]}),
    .q({\PWM2/pnumr[14]_keep ,\PWM2/RemaTxNum[14]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg2_b15|PWM2/reg3_b15  (
    .a({\PWM2/pnumr [15],_al_u1889_o}),
    .b({pnum2[15],\PWM2/n24 }),
    .c({pnum2[32],pnumcnt2[15]}),
    .clk(clk100m),
    .d({pwm_start_stop[18],\PWM2/pnumr [15]}),
    .e({open_n4020,pwm_start_stop[18]}),
    .q({\PWM2/pnumr[15]_keep ,\PWM2/RemaTxNum[15]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg2_b16|PWM2/reg2_b23  (
    .a({\PWM2/pnumr [16],\PWM2/pnumr [23]}),
    .b({pnum2[16],pnum2[23]}),
    .c({pnum2[32],pnum2[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[18],pwm_start_stop[18]}),
    .q({\PWM2/pnumr[16]_keep ,\PWM2/pnumr[23]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg2_b17|PWM2/reg2_b20  (
    .a({\PWM2/pnumr [17],\PWM2/pnumr [20]}),
    .b({pnum2[17],pnum2[20]}),
    .c({pnum2[32],pnum2[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[18],pwm_start_stop[18]}),
    .q({\PWM2/pnumr[17]_keep ,\PWM2/pnumr[20]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg2_b18|PWM2/reg3_b18  (
    .a({\PWM2/pnumr [18],_al_u1883_o}),
    .b({pnum2[18],\PWM2/n24 }),
    .c({pnum2[32],pnumcnt2[18]}),
    .clk(clk100m),
    .d({pwm_start_stop[18],\PWM2/pnumr [18]}),
    .e({open_n4084,pwm_start_stop[18]}),
    .q({\PWM2/pnumr[18]_keep ,\PWM2/RemaTxNum[18]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg2_b19|PWM2/reg3_b19  (
    .a({\PWM2/pnumr [19],_al_u1881_o}),
    .b({pnum2[19],\PWM2/n24 }),
    .c({pnum2[32],pnumcnt2[19]}),
    .clk(clk100m),
    .d({pwm_start_stop[18],\PWM2/pnumr [19]}),
    .e({open_n4106,pwm_start_stop[18]}),
    .q({\PWM2/pnumr[19]_keep ,\PWM2/RemaTxNum[19]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg2_b1|PWM2/reg2_b2  (
    .a({\PWM2/pnumr [1],\PWM2/pnumr [2]}),
    .b({pnum2[1],pnum2[2]}),
    .c({pnum2[32],pnum2[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[18],pwm_start_stop[18]}),
    .q({\PWM2/pnumr[1]_keep ,\PWM2/pnumr[2]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg2_b21|PWM2/reg3_b21  (
    .a({\PWM2/pnumr [21],_al_u1875_o}),
    .b({pnum2[21],\PWM2/n24 }),
    .c({pnum2[32],pnumcnt2[21]}),
    .clk(clk100m),
    .d({pwm_start_stop[18],\PWM2/pnumr [21]}),
    .e({open_n4151,pwm_start_stop[18]}),
    .q({\PWM2/pnumr[21]_keep ,\PWM2/RemaTxNum[21]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg2_b22|PWM2/reg3_b22  (
    .a({\PWM2/pnumr [22],_al_u1873_o}),
    .b({pnum2[22],\PWM2/n24 }),
    .c({pnum2[32],pnumcnt2[22]}),
    .clk(clk100m),
    .d({pwm_start_stop[18],\PWM2/pnumr [22]}),
    .e({open_n4173,pwm_start_stop[18]}),
    .q({\PWM2/pnumr[22]_keep ,\PWM2/RemaTxNum[22]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg2_b24|PWM2/reg2_b30  (
    .a({\PWM2/pnumr [24],\PWM2/pnumr [30]}),
    .b({pnum2[24],pnum2[30]}),
    .c({pnum2[32],pnum2[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[18],pwm_start_stop[18]}),
    .q({\PWM2/pnumr[24]_keep ,\PWM2/pnumr[30]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg2_b25|PWM2/reg2_b29  (
    .a({\PWM2/pnumr [25],\PWM2/pnumr [29]}),
    .b({pnum2[25],pnum2[29]}),
    .c({pnum2[32],pnum2[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[18],pwm_start_stop[18]}),
    .q({\PWM2/pnumr[25]_keep ,\PWM2/pnumr[29]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg2_b26|PWM2/reg2_b28  (
    .a({\PWM2/pnumr [26],\PWM2/pnumr [28]}),
    .b({pnum2[26],pnum2[28]}),
    .c({pnum2[32],pnum2[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[18],pwm_start_stop[18]}),
    .q({\PWM2/pnumr[26]_keep ,\PWM2/pnumr[28]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~((~0*~(B*A)))+D*C*~((~0*~(B*A)))+~(D)*C*(~0*~(B*A))+D*C*(~0*~(B*A)))"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(D*~(C)*~((~1*~(B*A)))+D*C*~((~1*~(B*A)))+~(D)*C*(~1*~(B*A))+D*C*(~1*~(B*A)))"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111100001110000),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg2_b31|PWM2/dir_reg  (
    .a({\PWM2/pnumr [31],\PWM2/n24 }),
    .b({pnum2[31],\PWM2/n25_neg_lutinv }),
    .c({pnum2[32],dir_pad[2]}),
    .clk(clk100m),
    .d({pwm_start_stop[18],\PWM2/pnumr [31]}),
    .e({open_n4260,pwm_start_stop[18]}),
    .q({\PWM2/pnumr[31]_keep ,\PWM2/dir_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg2_b4|PWM2/reg3_b4  (
    .a({\PWM2/pnumr [4],_al_u1867_o}),
    .b({pnum2[32],\PWM2/n24 }),
    .c({pnum2[4],pnumcnt2[4]}),
    .clk(clk100m),
    .d({pwm_start_stop[18],\PWM2/pnumr [4]}),
    .e({open_n4282,pwm_start_stop[18]}),
    .q({\PWM2/pnumr[4]_keep ,\PWM2/RemaTxNum[4]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg2_b5|PWM2/reg3_b5  (
    .a({\PWM2/pnumr [5],_al_u1865_o}),
    .b({pnum2[32],\PWM2/n24 }),
    .c({pnum2[5],pnumcnt2[5]}),
    .clk(clk100m),
    .d({pwm_start_stop[18],\PWM2/pnumr [5]}),
    .e({open_n4304,pwm_start_stop[18]}),
    .q({\PWM2/pnumr[5]_keep ,\PWM2/RemaTxNum[5]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg2_b8|PWM2/reg3_b8  (
    .a({\PWM2/pnumr [8],_al_u1859_o}),
    .b({pnum2[32],\PWM2/n24 }),
    .c({pnum2[8],pnumcnt2[8]}),
    .clk(clk100m),
    .d({pwm_start_stop[18],\PWM2/pnumr [8]}),
    .e({open_n4326,pwm_start_stop[18]}),
    .q({\PWM2/pnumr[8]_keep ,\PWM2/RemaTxNum[8]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg2_b9|PWM2/reg3_b9  (
    .a({\PWM2/pnumr [9],_al_u1857_o}),
    .b({pnum2[32],\PWM2/n24 }),
    .c({pnum2[9],pnumcnt2[9]}),
    .clk(clk100m),
    .d({pwm_start_stop[18],\PWM2/pnumr [9]}),
    .e({open_n4348,pwm_start_stop[18]}),
    .q({\PWM2/pnumr[9]_keep ,\PWM2/RemaTxNum[9]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg3_b0  (
    .a({_al_u1903_o,_al_u1903_o}),
    .b({\PWM2/n24 ,\PWM2/n24 }),
    .c({pnumcnt2[0],pnumcnt2[0]}),
    .clk(clk100m),
    .d({\PWM2/pnumr [0],\PWM2/pnumr [0]}),
    .mi({open_n4380,pwm_start_stop[18]}),
    .q({open_n4387,\PWM2/RemaTxNum[0]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg3_b1  (
    .a({_al_u1901_o,_al_u1901_o}),
    .b({\PWM2/n24 ,\PWM2/n24 }),
    .c({pnumcnt2[1],pnumcnt2[1]}),
    .clk(clk100m),
    .d({\PWM2/pnumr [1],\PWM2/pnumr [1]}),
    .mi({open_n4399,pwm_start_stop[18]}),
    .q({open_n4406,\PWM2/RemaTxNum[1]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg3_b12  (
    .a({_al_u1895_o,_al_u1895_o}),
    .b({\PWM2/n24 ,\PWM2/n24 }),
    .c({pnumcnt2[12],pnumcnt2[12]}),
    .clk(clk100m),
    .d({\PWM2/pnumr [12],\PWM2/pnumr [12]}),
    .mi({open_n4418,pwm_start_stop[18]}),
    .q({open_n4425,\PWM2/RemaTxNum[12]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg3_b13  (
    .a({_al_u1893_o,_al_u1893_o}),
    .b({\PWM2/n24 ,\PWM2/n24 }),
    .c({pnumcnt2[13],pnumcnt2[13]}),
    .clk(clk100m),
    .d({\PWM2/pnumr [13],\PWM2/pnumr [13]}),
    .mi({open_n4437,pwm_start_stop[18]}),
    .q({open_n4444,\PWM2/RemaTxNum[13]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg3_b16  (
    .a({_al_u1887_o,_al_u1887_o}),
    .b({\PWM2/n24 ,\PWM2/n24 }),
    .c({pnumcnt2[16],pnumcnt2[16]}),
    .clk(clk100m),
    .d({\PWM2/pnumr [16],\PWM2/pnumr [16]}),
    .mi({open_n4456,pwm_start_stop[18]}),
    .q({open_n4463,\PWM2/RemaTxNum[16]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg3_b17  (
    .a({_al_u1885_o,_al_u1885_o}),
    .b({\PWM2/n24 ,\PWM2/n24 }),
    .c({pnumcnt2[17],pnumcnt2[17]}),
    .clk(clk100m),
    .d({\PWM2/pnumr [17],\PWM2/pnumr [17]}),
    .mi({open_n4475,pwm_start_stop[18]}),
    .q({open_n4482,\PWM2/RemaTxNum[17]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg3_b2  (
    .a({_al_u1879_o,_al_u1879_o}),
    .b({\PWM2/n24 ,\PWM2/n24 }),
    .c({pnumcnt2[2],pnumcnt2[2]}),
    .clk(clk100m),
    .d({\PWM2/pnumr [2],\PWM2/pnumr [2]}),
    .mi({open_n4494,pwm_start_stop[18]}),
    .q({open_n4501,\PWM2/RemaTxNum[2]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg3_b20  (
    .a({_al_u1877_o,_al_u1877_o}),
    .b({\PWM2/n24 ,\PWM2/n24 }),
    .c({pnumcnt2[20],pnumcnt2[20]}),
    .clk(clk100m),
    .d({\PWM2/pnumr [20],\PWM2/pnumr [20]}),
    .mi({open_n4513,pwm_start_stop[18]}),
    .q({open_n4520,\PWM2/RemaTxNum[20]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg3_b23  (
    .a({_al_u1871_o,_al_u1871_o}),
    .b({\PWM2/n24 ,\PWM2/n24 }),
    .c({pnumcnt2[23],pnumcnt2[23]}),
    .clk(clk100m),
    .d({\PWM2/pnumr [23],\PWM2/pnumr [23]}),
    .mi({open_n4532,pwm_start_stop[18]}),
    .q({open_n4539,\PWM2/RemaTxNum[23]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg3_b3  (
    .a({_al_u1869_o,_al_u1869_o}),
    .b({\PWM2/n24 ,\PWM2/n24 }),
    .c({pnumcnt2[3],pnumcnt2[3]}),
    .clk(clk100m),
    .d({\PWM2/pnumr [3],\PWM2/pnumr [3]}),
    .mi({open_n4551,pwm_start_stop[18]}),
    .q({open_n4558,\PWM2/RemaTxNum[3]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg3_b6  (
    .a({_al_u1863_o,_al_u1863_o}),
    .b({\PWM2/n24 ,\PWM2/n24 }),
    .c({pnumcnt2[6],pnumcnt2[6]}),
    .clk(clk100m),
    .d({\PWM2/pnumr [6],\PWM2/pnumr [6]}),
    .mi({open_n4570,pwm_start_stop[18]}),
    .q({open_n4577,\PWM2/RemaTxNum[6]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/reg3_b7  (
    .a({_al_u1861_o,_al_u1861_o}),
    .b({\PWM2/n24 ,\PWM2/n24 }),
    .c({pnumcnt2[7],pnumcnt2[7]}),
    .clk(clk100m),
    .d({\PWM2/pnumr [7],\PWM2/pnumr [7]}),
    .mi({open_n4589,pwm_start_stop[18]}),
    .q({open_n4596,\PWM2/RemaTxNum[7]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_LSLICE #(
    //.MACRO("PWM2/sub0/ucin_al_u3377"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM2/sub0/u11_al_u3380  (
    .a({\PWM2/FreCnt [13],\PWM2/FreCnt [11]}),
    .b({\PWM2/FreCnt [14],\PWM2/FreCnt [12]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM2/sub0/c11 ),
    .f({\PWM2/n12 [13],\PWM2/n12 [11]}),
    .fco(\PWM2/sub0/c15 ),
    .fx({\PWM2/n12 [14],\PWM2/n12 [12]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM2/sub0/ucin_al_u3377"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM2/sub0/u15_al_u3381  (
    .a({\PWM2/FreCnt [17],\PWM2/FreCnt [15]}),
    .b({\PWM2/FreCnt [18],\PWM2/FreCnt [16]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM2/sub0/c15 ),
    .f({\PWM2/n12 [17],\PWM2/n12 [15]}),
    .fco(\PWM2/sub0/c19 ),
    .fx({\PWM2/n12 [18],\PWM2/n12 [16]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM2/sub0/ucin_al_u3377"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM2/sub0/u19_al_u3382  (
    .a({\PWM2/FreCnt [21],\PWM2/FreCnt [19]}),
    .b({\PWM2/FreCnt [22],\PWM2/FreCnt [20]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM2/sub0/c19 ),
    .f({\PWM2/n12 [21],\PWM2/n12 [19]}),
    .fco(\PWM2/sub0/c23 ),
    .fx({\PWM2/n12 [22],\PWM2/n12 [20]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM2/sub0/ucin_al_u3377"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM2/sub0/u23_al_u3383  (
    .a({\PWM2/FreCnt [25],\PWM2/FreCnt [23]}),
    .b({\PWM2/FreCnt [26],\PWM2/FreCnt [24]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM2/sub0/c23 ),
    .f({\PWM2/n12 [25],\PWM2/n12 [23]}),
    .fx({\PWM2/n12 [26],\PWM2/n12 [24]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM2/sub0/ucin_al_u3377"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM2/sub0/u3_al_u3378  (
    .a({\PWM2/FreCnt [5],\PWM2/FreCnt [3]}),
    .b({\PWM2/FreCnt [6],\PWM2/FreCnt [4]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM2/sub0/c3 ),
    .f({\PWM2/n12 [5],\PWM2/n12 [3]}),
    .fco(\PWM2/sub0/c7 ),
    .fx({\PWM2/n12 [6],\PWM2/n12 [4]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM2/sub0/ucin_al_u3377"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM2/sub0/u7_al_u3379  (
    .a({\PWM2/FreCnt [9],\PWM2/FreCnt [7]}),
    .b({\PWM2/FreCnt [10],\PWM2/FreCnt [8]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM2/sub0/c7 ),
    .f({\PWM2/n12 [9],\PWM2/n12 [7]}),
    .fco(\PWM2/sub0/c11 ),
    .fx({\PWM2/n12 [10],\PWM2/n12 [8]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM2/sub0/ucin_al_u3377"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'h0005),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM2/sub0/ucin_al_u3377  (
    .a({\PWM2/FreCnt [1],1'b0}),
    .b({\PWM2/FreCnt [2],\PWM2/FreCnt [0]}),
    .c(2'b11),
    .ce(\U_AHB/n8 ),
    .clk(clk100m),
    .d(2'b01),
    .e(2'b01),
    .mi({open_n4707,\U_AHB/h2h_hwdata [2]}),
    .f({\PWM2/n12 [1],open_n4720}),
    .fco(\PWM2/sub0/c3 ),
    .fx({\PWM2/n12 [2],\PWM2/n12 [0]}),
    .q({open_n4721,freq2[2]}));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM2/sub1/u0|PWM2/sub1/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("SUB_CARRY"),
    .INIT_LUT0(16'b0000000000000101),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM2/sub1/u0|PWM2/sub1/ucin  (
    .a({pnumcnt2[0],1'b0}),
    .b({1'b1,open_n4722}),
    .f({\PWM2/n26 [0],open_n4742}),
    .fco(\PWM2/sub1/c1 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM2/sub1/u0|PWM2/sub1/ucin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM2/sub1/u10|PWM2/sub1/u9  (
    .a(pnumcnt2[10:9]),
    .b(2'b00),
    .fci(\PWM2/sub1/c9 ),
    .f(\PWM2/n26 [10:9]),
    .fco(\PWM2/sub1/c11 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM2/sub1/u0|PWM2/sub1/ucin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM2/sub1/u12|PWM2/sub1/u11  (
    .a(pnumcnt2[12:11]),
    .b(2'b00),
    .fci(\PWM2/sub1/c11 ),
    .f(\PWM2/n26 [12:11]),
    .fco(\PWM2/sub1/c13 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM2/sub1/u0|PWM2/sub1/ucin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM2/sub1/u14|PWM2/sub1/u13  (
    .a(pnumcnt2[14:13]),
    .b(2'b00),
    .fci(\PWM2/sub1/c13 ),
    .f(\PWM2/n26 [14:13]),
    .fco(\PWM2/sub1/c15 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM2/sub1/u0|PWM2/sub1/ucin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM2/sub1/u16|PWM2/sub1/u15  (
    .a(pnumcnt2[16:15]),
    .b(2'b00),
    .fci(\PWM2/sub1/c15 ),
    .f(\PWM2/n26 [16:15]),
    .fco(\PWM2/sub1/c17 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM2/sub1/u0|PWM2/sub1/ucin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM2/sub1/u18|PWM2/sub1/u17  (
    .a(pnumcnt2[18:17]),
    .b(2'b00),
    .fci(\PWM2/sub1/c17 ),
    .f(\PWM2/n26 [18:17]),
    .fco(\PWM2/sub1/c19 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM2/sub1/u0|PWM2/sub1/ucin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM2/sub1/u20|PWM2/sub1/u19  (
    .a(pnumcnt2[20:19]),
    .b(2'b00),
    .fci(\PWM2/sub1/c19 ),
    .f(\PWM2/n26 [20:19]),
    .fco(\PWM2/sub1/c21 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM2/sub1/u0|PWM2/sub1/ucin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM2/sub1/u22|PWM2/sub1/u21  (
    .a(pnumcnt2[22:21]),
    .b(2'b00),
    .fci(\PWM2/sub1/c21 ),
    .f(\PWM2/n26 [22:21]),
    .fco(\PWM2/sub1/c23 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM2/sub1/u0|PWM2/sub1/ucin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM2/sub1/u23_al_u3470  (
    .a({open_n4901,pnumcnt2[23]}),
    .b({open_n4902,1'b0}),
    .fci(\PWM2/sub1/c23 ),
    .f({open_n4921,\PWM2/n26 [23]}));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM2/sub1/u0|PWM2/sub1/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM2/sub1/u2|PWM2/sub1/u1  (
    .a(pnumcnt2[2:1]),
    .b(2'b00),
    .fci(\PWM2/sub1/c1 ),
    .f(\PWM2/n26 [2:1]),
    .fco(\PWM2/sub1/c3 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM2/sub1/u0|PWM2/sub1/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM2/sub1/u4|PWM2/sub1/u3  (
    .a(pnumcnt2[4:3]),
    .b(2'b00),
    .fci(\PWM2/sub1/c3 ),
    .f(\PWM2/n26 [4:3]),
    .fco(\PWM2/sub1/c5 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM2/sub1/u0|PWM2/sub1/ucin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM2/sub1/u6|PWM2/sub1/u5  (
    .a(pnumcnt2[6:5]),
    .b(2'b00),
    .fci(\PWM2/sub1/c5 ),
    .f(\PWM2/n26 [6:5]),
    .fco(\PWM2/sub1/c7 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM2/sub1/u0|PWM2/sub1/ucin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM2/sub1/u8|PWM2/sub1/u7  (
    .a(pnumcnt2[8:7]),
    .b(2'b00),
    .fci(\PWM2/sub1/c7 ),
    .f(\PWM2/n26 [8:7]),
    .fco(\PWM2/sub1/c9 ));
  // src/OnePWM.v(26)
  // src/OnePWM.v(26)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*~(~D*B*~A))"),
    //.LUT1("(C*~(~D*B*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000010110000),
    .INIT_LUT1(16'b1111000010110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \PWM3/State_reg|PWMC/State_reg  (
    .a({_al_u3016_o,_al_u3043_o}),
    .b({\PWM3/n0_lutinv ,\PWMC/n0_lutinv }),
    .c({_al_u3017_o,_al_u3044_o}),
    .clk(clk100m),
    .d({pwm_start_stop[19],pwm_start_stop[28]}),
    .sr(rstn),
    .q({pwm_state_read[3],pwm_state_read[12]}));  // src/OnePWM.v(26)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[0]  (
    .i(\PWM3/RemaTxNum[0]_keep ),
    .o(pnumcnt3[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[10]  (
    .i(\PWM3/RemaTxNum[10]_keep ),
    .o(pnumcnt3[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[11]  (
    .i(\PWM3/RemaTxNum[11]_keep ),
    .o(pnumcnt3[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[12]  (
    .i(\PWM3/RemaTxNum[12]_keep ),
    .o(pnumcnt3[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[13]  (
    .i(\PWM3/RemaTxNum[13]_keep ),
    .o(pnumcnt3[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[14]  (
    .i(\PWM3/RemaTxNum[14]_keep ),
    .o(pnumcnt3[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[15]  (
    .i(\PWM3/RemaTxNum[15]_keep ),
    .o(pnumcnt3[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[16]  (
    .i(\PWM3/RemaTxNum[16]_keep ),
    .o(pnumcnt3[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[17]  (
    .i(\PWM3/RemaTxNum[17]_keep ),
    .o(pnumcnt3[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[18]  (
    .i(\PWM3/RemaTxNum[18]_keep ),
    .o(pnumcnt3[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[19]  (
    .i(\PWM3/RemaTxNum[19]_keep ),
    .o(pnumcnt3[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[1]  (
    .i(\PWM3/RemaTxNum[1]_keep ),
    .o(pnumcnt3[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[20]  (
    .i(\PWM3/RemaTxNum[20]_keep ),
    .o(pnumcnt3[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[21]  (
    .i(\PWM3/RemaTxNum[21]_keep ),
    .o(pnumcnt3[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[22]  (
    .i(\PWM3/RemaTxNum[22]_keep ),
    .o(pnumcnt3[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[23]  (
    .i(\PWM3/RemaTxNum[23]_keep ),
    .o(pnumcnt3[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[2]  (
    .i(\PWM3/RemaTxNum[2]_keep ),
    .o(pnumcnt3[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[3]  (
    .i(\PWM3/RemaTxNum[3]_keep ),
    .o(pnumcnt3[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[4]  (
    .i(\PWM3/RemaTxNum[4]_keep ),
    .o(pnumcnt3[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[5]  (
    .i(\PWM3/RemaTxNum[5]_keep ),
    .o(pnumcnt3[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[6]  (
    .i(\PWM3/RemaTxNum[6]_keep ),
    .o(pnumcnt3[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[7]  (
    .i(\PWM3/RemaTxNum[7]_keep ),
    .o(pnumcnt3[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[8]  (
    .i(\PWM3/RemaTxNum[8]_keep ),
    .o(pnumcnt3[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[9]  (
    .i(\PWM3/RemaTxNum[9]_keep ),
    .o(pnumcnt3[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_dir  (
    .i(\PWM3/dir_keep ),
    .o(dir_pad[3]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[0]  (
    .i(\PWM3/pnumr[0]_keep ),
    .o(\PWM3/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[10]  (
    .i(\PWM3/pnumr[10]_keep ),
    .o(\PWM3/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[11]  (
    .i(\PWM3/pnumr[11]_keep ),
    .o(\PWM3/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[12]  (
    .i(\PWM3/pnumr[12]_keep ),
    .o(\PWM3/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[13]  (
    .i(\PWM3/pnumr[13]_keep ),
    .o(\PWM3/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[14]  (
    .i(\PWM3/pnumr[14]_keep ),
    .o(\PWM3/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[15]  (
    .i(\PWM3/pnumr[15]_keep ),
    .o(\PWM3/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[16]  (
    .i(\PWM3/pnumr[16]_keep ),
    .o(\PWM3/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[17]  (
    .i(\PWM3/pnumr[17]_keep ),
    .o(\PWM3/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[18]  (
    .i(\PWM3/pnumr[18]_keep ),
    .o(\PWM3/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[19]  (
    .i(\PWM3/pnumr[19]_keep ),
    .o(\PWM3/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[1]  (
    .i(\PWM3/pnumr[1]_keep ),
    .o(\PWM3/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[20]  (
    .i(\PWM3/pnumr[20]_keep ),
    .o(\PWM3/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[21]  (
    .i(\PWM3/pnumr[21]_keep ),
    .o(\PWM3/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[22]  (
    .i(\PWM3/pnumr[22]_keep ),
    .o(\PWM3/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[23]  (
    .i(\PWM3/pnumr[23]_keep ),
    .o(\PWM3/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[24]  (
    .i(\PWM3/pnumr[24]_keep ),
    .o(\PWM3/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[25]  (
    .i(\PWM3/pnumr[25]_keep ),
    .o(\PWM3/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[26]  (
    .i(\PWM3/pnumr[26]_keep ),
    .o(\PWM3/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[27]  (
    .i(\PWM3/pnumr[27]_keep ),
    .o(\PWM3/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[28]  (
    .i(\PWM3/pnumr[28]_keep ),
    .o(\PWM3/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[29]  (
    .i(\PWM3/pnumr[29]_keep ),
    .o(\PWM3/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[2]  (
    .i(\PWM3/pnumr[2]_keep ),
    .o(\PWM3/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[30]  (
    .i(\PWM3/pnumr[30]_keep ),
    .o(\PWM3/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[31]  (
    .i(\PWM3/pnumr[31]_keep ),
    .o(\PWM3/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[3]  (
    .i(\PWM3/pnumr[3]_keep ),
    .o(\PWM3/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[4]  (
    .i(\PWM3/pnumr[4]_keep ),
    .o(\PWM3/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[5]  (
    .i(\PWM3/pnumr[5]_keep ),
    .o(\PWM3/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[6]  (
    .i(\PWM3/pnumr[6]_keep ),
    .o(\PWM3/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[7]  (
    .i(\PWM3/pnumr[7]_keep ),
    .o(\PWM3/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[8]  (
    .i(\PWM3/pnumr[8]_keep ),
    .o(\PWM3/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[9]  (
    .i(\PWM3/pnumr[9]_keep ),
    .o(\PWM3/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pwm  (
    .i(\PWM3/pwm_keep ),
    .o(pwm_pad[3]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_stopreq  (
    .i(\PWM3/stopreq_keep ),
    .o(\PWM3/stopreq ));  // src/OnePWM.v(14)
  EF2_PHY_MSLICE #(
    //.LUT0("~(~0*~(D*C*B*A))"),
    //.LUT1("~(~1*~(D*C*B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b1111111111111111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM3/pwm_reg  (
    .a({_al_u1418_o,_al_u1418_o}),
    .b({_al_u1424_o,_al_u1424_o}),
    .c({_al_u1426_o,_al_u1426_o}),
    .clk(clk100m),
    .d({_al_u1428_o,_al_u1428_o}),
    .mi({open_n5044,pwm_pad[3]}),
    .sr(\PWM3/u14_sel_is_1_o ),
    .q({open_n5050,\PWM3/pwm_keep }));  // src/OnePWM.v(45)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM3/reg0_b0|PWM3/reg0_b12  (
    .b({\PWM3/n12 [0],\PWM3/n12 [12]}),
    .c({freq3[0],freq3[12]}),
    .clk(clk100m),
    .d({\PWM3/n0_lutinv ,\PWM3/n0_lutinv }),
    .sr(\PWM3/n11 ),
    .q({\PWM3/FreCnt [0],\PWM3/FreCnt [12]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM3/reg0_b10|PWM3/reg0_b9  (
    .b(\PWM3/n12 [10:9]),
    .c(freq3[10:9]),
    .clk(clk100m),
    .d({\PWM3/n0_lutinv ,\PWM3/n0_lutinv }),
    .sr(\PWM3/n11 ),
    .q(\PWM3/FreCnt [10:9]));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM3/reg0_b11|PWM3/reg0_b7  (
    .b({\PWM3/n12 [11],\PWM3/n12 [7]}),
    .c({freq3[11],freq3[7]}),
    .clk(clk100m),
    .d({\PWM3/n0_lutinv ,\PWM3/n0_lutinv }),
    .sr(\PWM3/n11 ),
    .q({\PWM3/FreCnt [11],\PWM3/FreCnt [7]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM3/reg0_b13|PWM3/reg0_b3  (
    .b({\PWM3/n12 [13],\PWM3/n12 [3]}),
    .c({freq3[13],freq3[3]}),
    .clk(clk100m),
    .d({\PWM3/n0_lutinv ,\PWM3/n0_lutinv }),
    .sr(\PWM3/n11 ),
    .q({\PWM3/FreCnt [13],\PWM3/FreCnt [3]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM3/reg0_b14|PWM3/reg0_b25  (
    .b({\PWM3/n12 [14],\PWM3/n12 [25]}),
    .c({freq3[14],freq3[25]}),
    .clk(clk100m),
    .d({\PWM3/n0_lutinv ,\PWM3/n0_lutinv }),
    .sr(\PWM3/n11 ),
    .q({\PWM3/FreCnt [14],\PWM3/FreCnt [25]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM3/reg0_b16|PWM3/reg0_b21  (
    .b({\PWM3/n12 [16],\PWM3/n12 [21]}),
    .c({freq3[16],freq3[21]}),
    .clk(clk100m),
    .d({\PWM3/n0_lutinv ,\PWM3/n0_lutinv }),
    .sr(\PWM3/n11 ),
    .q({\PWM3/FreCnt [16],\PWM3/FreCnt [21]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM3/reg0_b17|PWM3/reg0_b19  (
    .b({\PWM3/n12 [17],\PWM3/n12 [19]}),
    .c({freq3[17],freq3[19]}),
    .clk(clk100m),
    .d({\PWM3/n0_lutinv ,\PWM3/n0_lutinv }),
    .sr(\PWM3/n11 ),
    .q({\PWM3/FreCnt [17],\PWM3/FreCnt [19]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM3/reg0_b18|PWM3/reg0_b1  (
    .b({\PWM3/n12 [18],\PWM3/n12 [1]}),
    .c({freq3[18],freq3[1]}),
    .clk(clk100m),
    .d({\PWM3/n0_lutinv ,\PWM3/n0_lutinv }),
    .sr(\PWM3/n11 ),
    .q({\PWM3/FreCnt [18],\PWM3/FreCnt [1]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM3/reg0_b20|PWM3/reg0_b8  (
    .b({\PWM3/n12 [20],\PWM3/n12 [8]}),
    .c({freq3[20],freq3[8]}),
    .clk(clk100m),
    .d({\PWM3/n0_lutinv ,\PWM3/n0_lutinv }),
    .sr(\PWM3/n11 ),
    .q({\PWM3/FreCnt [20],\PWM3/FreCnt [8]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM3/reg0_b22|PWM3/reg0_b6  (
    .b({\PWM3/n12 [22],\PWM3/n12 [6]}),
    .c({freq3[22],freq3[6]}),
    .clk(clk100m),
    .d({\PWM3/n0_lutinv ,\PWM3/n0_lutinv }),
    .sr(\PWM3/n11 ),
    .q({\PWM3/FreCnt [22],\PWM3/FreCnt [6]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM3/reg0_b23|PWM3/reg0_b5  (
    .b({\PWM3/n12 [23],\PWM3/n12 [5]}),
    .c({freq3[23],freq3[5]}),
    .clk(clk100m),
    .d({\PWM3/n0_lutinv ,\PWM3/n0_lutinv }),
    .sr(\PWM3/n11 ),
    .q({\PWM3/FreCnt [23],\PWM3/FreCnt [5]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM3/reg0_b24|PWM3/reg0_b4  (
    .b({\PWM3/n12 [24],\PWM3/n12 [4]}),
    .c({freq3[24],freq3[4]}),
    .clk(clk100m),
    .d({\PWM3/n0_lutinv ,\PWM3/n0_lutinv }),
    .sr(\PWM3/n11 ),
    .q({\PWM3/FreCnt [24],\PWM3/FreCnt [4]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM3/reg0_b2|PWM3/reg0_b26  (
    .b({\PWM3/n12 [2],\PWM3/n12 [26]}),
    .c({freq3[2],freq3[26]}),
    .clk(clk100m),
    .d({\PWM3/n0_lutinv ,\PWM3/n0_lutinv }),
    .sr(\PWM3/n11 ),
    .q({\PWM3/FreCnt [2],\PWM3/FreCnt [26]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~A*~(~D*C)*~(0@B))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(~A*~(~D*C)*~(1@B))"),
    //.LUTG1("(C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0001000100000001),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0100010000000100),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg1_b10|PWM3/reg1_b21  (
    .a({open_n5335,_al_u1996_o}),
    .b({open_n5336,\PWM3/FreCnt [20]}),
    .c({\PWM3/FreCntr [10],\PWM3/FreCnt [9]}),
    .ce(\PWM3/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM3/FreCnt [9],\PWM3/FreCntr [10]}),
    .e({open_n5337,\PWM3/FreCntr [21]}),
    .mi({freq3[10],freq3[21]}),
    .f({_al_u1998_o,_al_u1997_o}),
    .q({\PWM3/FreCntr [10],\PWM3/FreCntr [21]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(B*A*~(D@C))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(B*A*~(D@C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1000000000001000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg1_b11|PWM3/reg1_b0  (
    .a({_al_u1993_o,open_n5354}),
    .b({_al_u1994_o,open_n5355}),
    .c({\PWM3/FreCnt [10],\PWM3/n11 }),
    .ce(\PWM3/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM3/FreCntr [11],\PWM3/n0_lutinv }),
    .mi({freq3[11],freq3[0]}),
    .f({_al_u1995_o,\PWM3/mux3_b0_sel_is_3_o }),
    .q({\PWM3/FreCntr [11],\PWM3/FreCntr [0]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~D*B)*~(C@A))"),
    //.LUTF1("(B*A*~(D@C))"),
    //.LUTG0("(~(~D*B)*~(C@A))"),
    //.LUTG1("(B*A*~(D@C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010010100100001),
    .INIT_LUTF1(16'b1000000000001000),
    .INIT_LUTG0(16'b1010010100100001),
    .INIT_LUTG1(16'b1000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg1_b12|PWM3/reg1_b7  (
    .a({_al_u2002_o,\PWM3/FreCnt [6]}),
    .b({_al_u2003_o,\PWM3/FreCnt [7]}),
    .c({\PWM3/FreCnt [11],\PWM3/FreCntr [7]}),
    .ce(\PWM3/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM3/FreCntr [12],\PWM3/FreCntr [8]}),
    .mi({freq3[12],freq3[7]}),
    .f({_al_u2004_o,_al_u1993_o}),
    .q({\PWM3/FreCntr [12],\PWM3/FreCntr [7]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(D@B)*~(C@A))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(~(D@B)*~(C@A))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000010000100001),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000010000100001),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg1_b15|PWM3/reg1_b25  (
    .a({\PWM3/FreCnt [14],\PWM3/FreCnt [2]}),
    .b({\PWM3/FreCnt [24],\PWM3/FreCnt [25]}),
    .c({\PWM3/FreCntr [15],\PWM3/FreCntr [2]}),
    .ce(\PWM3/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM3/FreCntr [25],\PWM3/FreCntr [25]}),
    .mi({freq3[15],freq3[25]}),
    .f({_al_u1987_o,_al_u1427_o}),
    .q({\PWM3/FreCntr [15],\PWM3/FreCntr [25]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~A*~(0@C)*~(D*~B))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~A*~(1@C)*~(D*~B))"),
    //.LUTG1("(~C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010000000101),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0100000001010000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg1_b17|PWM3/reg1_b19  (
    .a({open_n5410,_al_u1998_o}),
    .b({open_n5411,\PWM3/FreCnt [16]}),
    .c({\PWM3/FreCntr [17],\PWM3/FreCnt [18]}),
    .ce(\PWM3/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM3/FreCnt [16],\PWM3/FreCntr [17]}),
    .e({open_n5412,\PWM3/FreCntr [19]}),
    .mi({freq3[17],freq3[19]}),
    .f({_al_u2005_o,_al_u1999_o}),
    .q({\PWM3/FreCntr [17],\PWM3/FreCntr [19]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(D@B)*~(C@A))"),
    //.LUT1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000010000100001),
    .INIT_LUT1(16'b1000010000100001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg1_b1|PWM3/reg1_b23  (
    .a({\PWM3/FreCnt [0],\PWM3/FreCnt [22]}),
    .b({\PWM3/FreCnt [22],\PWM3/FreCnt [23]}),
    .c({\PWM3/FreCntr [1],\PWM3/FreCntr [22]}),
    .ce(\PWM3/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM3/FreCntr [23],\PWM3/FreCntr [23]}),
    .mi({freq3[1],freq3[23]}),
    .f({_al_u1985_o,_al_u1415_o}),
    .q({\PWM3/FreCntr [1],\PWM3/FreCntr [23]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~A*~(~0*C)*~(D@B))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(~A*~(~1*C)*~(D@B))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010000000001),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b0100010000010001),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg1_b20|PWM3/reg1_b18  (
    .a({\PWM3/FreCnt [20],_al_u2005_o}),
    .b({\PWM3/FreCnt [26],\PWM3/FreCnt [17]}),
    .c({\PWM3/FreCntr [20],\PWM3/FreCnt [19]}),
    .ce(\PWM3/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM3/FreCntr [26],\PWM3/FreCntr [18]}),
    .e({open_n5443,\PWM3/FreCntr [20]}),
    .mi({freq3[20],freq3[18]}),
    .f({_al_u1417_o,_al_u2006_o}),
    .q({\PWM3/FreCntr [20],\PWM3/FreCntr [18]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~B*~(0@C)*~(~D*A))"),
    //.LUTF1("(~(D*~B)*~(~C*A))"),
    //.LUTG0("(~B*~(1@C)*~(~D*A))"),
    //.LUTG1("(~(D*~B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001100000001),
    .INIT_LUTF1(16'b1100010011110101),
    .INIT_LUTG0(16'b0011000000010000),
    .INIT_LUTG1(16'b1100010011110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg1_b22|PWM3/reg1_b9  (
    .a({\PWM3/FreCnt [15],\PWM3/FreCnt [21]}),
    .b({\PWM3/FreCnt [21],\PWM3/FreCnt [26]}),
    .c({\PWM3/FreCntr [16],\PWM3/FreCnt [8]}),
    .ce(\PWM3/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM3/FreCntr [22],\PWM3/FreCntr [22]}),
    .e({open_n5460,\PWM3/FreCntr [9]}),
    .mi({freq3[22],freq3[9]}),
    .f({_al_u2001_o,_al_u1991_o}),
    .q({\PWM3/FreCntr [22],\PWM3/FreCntr [9]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~A*~(0@C)*~(D*~B))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(~A*~(1@C)*~(D*~B))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010000000101),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b0100000001010000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg1_b24|PWM3/reg1_b16  (
    .a({\PWM3/FreCnt [0],_al_u2007_o}),
    .b({\PWM3/FreCnt [24],\PWM3/FreCnt [15]}),
    .c({\PWM3/FreCntr [0],\PWM3/FreCnt [23]}),
    .ce(\PWM3/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM3/FreCntr [24],\PWM3/FreCntr [16]}),
    .e({open_n5477,\PWM3/FreCntr [24]}),
    .mi({freq3[24],freq3[16]}),
    .f({_al_u1421_o,_al_u2008_o}),
    .q({\PWM3/FreCntr [24],\PWM3/FreCntr [16]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(D*~B)*~(C*~A))"),
    //.LUT1("(~(~D*B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000110010101111),
    .INIT_LUT1(16'b1010111100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg1_b26|PWM3/reg1_b4  (
    .a({\PWM3/FreCnt [25],\PWM3/FreCnt [1]}),
    .b({\PWM3/FreCnt [3],\PWM3/FreCnt [3]}),
    .c({\PWM3/FreCntr [26],\PWM3/FreCntr [2]}),
    .ce(\PWM3/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM3/FreCntr [4],\PWM3/FreCntr [4]}),
    .mi({freq3[26],freq3[4]}),
    .f({_al_u2003_o,_al_u1989_o}),
    .q({\PWM3/FreCntr [26],\PWM3/FreCntr [4]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(~C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg1_b2|PWM3/reg1_b13  (
    .c({\PWM3/FreCntr [2],\PWM3/FreCntr [13]}),
    .ce(\PWM3/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM3/FreCnt [1],\PWM3/FreCnt [12]}),
    .mi({freq3[2],freq3[13]}),
    .f({_al_u2007_o,_al_u1996_o}),
    .q({\PWM3/FreCntr [2],\PWM3/FreCntr [13]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(D*~(C@B))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(D*~(C@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b1100001100000000),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1100001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg1_b6|PWM3/reg1_b5  (
    .a({open_n5526,_al_u1987_o}),
    .b({\PWM3/FreCnt [6],\PWM3/FreCnt [4]}),
    .c({\PWM3/FreCntr [6],\PWM3/FreCnt [5]}),
    .ce(\PWM3/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({_al_u1419_o,\PWM3/FreCntr [5]}),
    .e({open_n5527,\PWM3/FreCntr [6]}),
    .mi(freq3[6:5]),
    .f({_al_u1420_o,_al_u1988_o}),
    .q(\PWM3/FreCntr [6:5]));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*~C)*~(D*~B))"),
    //.LUTF1("(~(D*~B)*~(~C*A))"),
    //.LUTG0("(A*~(1*~C)*~(D*~B))"),
    //.LUTG1("(~(D*~B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000100010101010),
    .INIT_LUTF1(16'b1100010011110101),
    .INIT_LUTG0(16'b1000000010100000),
    .INIT_LUTG1(16'b1100010011110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg1_b8|PWM3/reg1_b14  (
    .a({\PWM3/FreCnt [13],_al_u2001_o}),
    .b({\PWM3/FreCnt [7],\PWM3/FreCnt [13]}),
    .c({\PWM3/FreCntr [14],\PWM3/FreCnt [19]}),
    .ce(\PWM3/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM3/FreCntr [8],\PWM3/FreCntr [14]}),
    .e({open_n5544,\PWM3/FreCntr [20]}),
    .mi({freq3[8],freq3[14]}),
    .f({_al_u1994_o,_al_u2002_o}),
    .q({\PWM3/FreCntr [8],\PWM3/FreCntr [14]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011100010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011100010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg2_b0|PWM3/reg2_b8  (
    .a({\PWM3/pnumr [0],\PWM3/pnumr [8]}),
    .b({pnum3[0],pnum3[32]}),
    .c({pnum3[32],pnum3[8]}),
    .clk(clk100m),
    .d({pwm_start_stop[19],pwm_start_stop[19]}),
    .q({\PWM3/pnumr[0]_keep ,\PWM3/pnumr[8]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011100010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg2_b10|PWM3/reg2_b7  (
    .a({\PWM3/pnumr [10],\PWM3/pnumr [7]}),
    .b({pnum3[10],pnum3[32]}),
    .c({pnum3[32],pnum3[7]}),
    .clk(clk100m),
    .d({pwm_start_stop[19],pwm_start_stop[19]}),
    .q({\PWM3/pnumr[10]_keep ,\PWM3/pnumr[7]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg2_b11|PWM3/reg3_b11  (
    .a({\PWM3/pnumr [11],_al_u1977_o}),
    .b({pnum3[11],\PWM3/n24 }),
    .c({pnum3[32],pnumcnt3[11]}),
    .clk(clk100m),
    .d({pwm_start_stop[19],\PWM3/pnumr [11]}),
    .e({open_n5604,pwm_start_stop[19]}),
    .q({\PWM3/pnumr[11]_keep ,\PWM3/RemaTxNum[11]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg2_b12|PWM3/reg3_b12  (
    .a({\PWM3/pnumr [12],_al_u1975_o}),
    .b({pnum3[12],\PWM3/n24 }),
    .c({pnum3[32],pnumcnt3[12]}),
    .clk(clk100m),
    .d({pwm_start_stop[19],\PWM3/pnumr [12]}),
    .e({open_n5626,pwm_start_stop[19]}),
    .q({\PWM3/pnumr[12]_keep ,\PWM3/RemaTxNum[12]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011100010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg2_b13|PWM3/reg2_b4  (
    .a({\PWM3/pnumr [13],\PWM3/pnumr [4]}),
    .b({pnum3[13],pnum3[32]}),
    .c({pnum3[32],pnum3[4]}),
    .clk(clk100m),
    .d({pwm_start_stop[19],pwm_start_stop[19]}),
    .q({\PWM3/pnumr[13]_keep ,\PWM3/pnumr[4]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg2_b14|PWM3/reg2_b3  (
    .a({\PWM3/pnumr [14],\PWM3/pnumr [3]}),
    .b({pnum3[14],pnum3[3]}),
    .c({pnum3[32],pnum3[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[19],pwm_start_stop[19]}),
    .q({\PWM3/pnumr[14]_keep ,\PWM3/pnumr[3]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg2_b15|PWM3/reg3_b15  (
    .a({\PWM3/pnumr [15],_al_u1969_o}),
    .b({pnum3[15],\PWM3/n24 }),
    .c({pnum3[32],pnumcnt3[15]}),
    .clk(clk100m),
    .d({pwm_start_stop[19],\PWM3/pnumr [15]}),
    .e({open_n5690,pwm_start_stop[19]}),
    .q({\PWM3/pnumr[15]_keep ,\PWM3/RemaTxNum[15]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg2_b16|PWM3/reg3_b16  (
    .a({\PWM3/pnumr [16],_al_u1967_o}),
    .b({pnum3[16],\PWM3/n24 }),
    .c({pnum3[32],pnumcnt3[16]}),
    .clk(clk100m),
    .d({pwm_start_stop[19],\PWM3/pnumr [16]}),
    .e({open_n5712,pwm_start_stop[19]}),
    .q({\PWM3/pnumr[16]_keep ,\PWM3/RemaTxNum[16]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg2_b17|PWM3/reg2_b21  (
    .a({\PWM3/pnumr [17],\PWM3/pnumr [21]}),
    .b({pnum3[17],pnum3[21]}),
    .c({pnum3[32],pnum3[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[19],pwm_start_stop[19]}),
    .q({\PWM3/pnumr[17]_keep ,\PWM3/pnumr[21]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg2_b18|PWM3/reg2_b20  (
    .a({\PWM3/pnumr [18],\PWM3/pnumr [20]}),
    .b({pnum3[18],pnum3[20]}),
    .c({pnum3[32],pnum3[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[19],pwm_start_stop[19]}),
    .q({\PWM3/pnumr[18]_keep ,\PWM3/pnumr[20]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg2_b19|PWM3/reg3_b19  (
    .a({\PWM3/pnumr [19],_al_u1961_o}),
    .b({pnum3[19],\PWM3/n24 }),
    .c({pnum3[32],pnumcnt3[19]}),
    .clk(clk100m),
    .d({pwm_start_stop[19],\PWM3/pnumr [19]}),
    .e({open_n5776,pwm_start_stop[19]}),
    .q({\PWM3/pnumr[19]_keep ,\PWM3/RemaTxNum[19]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg2_b22|PWM3/reg3_b22  (
    .a({\PWM3/pnumr [22],_al_u1953_o}),
    .b({pnum3[22],\PWM3/n24 }),
    .c({pnum3[32],pnumcnt3[22]}),
    .clk(clk100m),
    .d({pwm_start_stop[19],\PWM3/pnumr [22]}),
    .e({open_n5798,pwm_start_stop[19]}),
    .q({\PWM3/pnumr[22]_keep ,\PWM3/RemaTxNum[22]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg2_b23|PWM3/reg3_b23  (
    .a({\PWM3/pnumr [23],_al_u1951_o}),
    .b({pnum3[23],\PWM3/n24 }),
    .c({pnum3[32],pnumcnt3[23]}),
    .clk(clk100m),
    .d({pwm_start_stop[19],\PWM3/pnumr [23]}),
    .e({open_n5820,pwm_start_stop[19]}),
    .q({\PWM3/pnumr[23]_keep ,\PWM3/RemaTxNum[23]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg2_b24|PWM3/reg2_b1  (
    .a({\PWM3/pnumr [24],\PWM3/pnumr [1]}),
    .b({pnum3[24],pnum3[1]}),
    .c({pnum3[32],pnum3[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[19],pwm_start_stop[19]}),
    .q({\PWM3/pnumr[24]_keep ,\PWM3/pnumr[1]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg2_b25|PWM3/reg2_b30  (
    .a({\PWM3/pnumr [25],\PWM3/pnumr [30]}),
    .b({pnum3[25],pnum3[30]}),
    .c({pnum3[32],pnum3[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[19],pwm_start_stop[19]}),
    .q({\PWM3/pnumr[25]_keep ,\PWM3/pnumr[30]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg2_b26|PWM3/reg2_b29  (
    .a({\PWM3/pnumr [26],\PWM3/pnumr [29]}),
    .b({pnum3[26],pnum3[29]}),
    .c({pnum3[32],pnum3[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[19],pwm_start_stop[19]}),
    .q({\PWM3/pnumr[26]_keep ,\PWM3/pnumr[29]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg2_b27|PWM3/reg2_b28  (
    .a({\PWM3/pnumr [27],\PWM3/pnumr [28]}),
    .b({pnum3[27],pnum3[28]}),
    .c({pnum3[32],pnum3[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[19],pwm_start_stop[19]}),
    .q({\PWM3/pnumr[27]_keep ,\PWM3/pnumr[28]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg2_b2|PWM3/reg3_b2  (
    .a({\PWM3/pnumr [2],_al_u1959_o}),
    .b({pnum3[2],\PWM3/n24 }),
    .c({pnum3[32],pnumcnt3[2]}),
    .clk(clk100m),
    .d({pwm_start_stop[19],\PWM3/pnumr [2]}),
    .e({open_n5926,pwm_start_stop[19]}),
    .q({\PWM3/pnumr[2]_keep ,\PWM3/RemaTxNum[2]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~((~0*~(B*A)))+D*C*~((~0*~(B*A)))+~(D)*C*(~0*~(B*A))+D*C*(~0*~(B*A)))"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(D*~(C)*~((~1*~(B*A)))+D*C*~((~1*~(B*A)))+~(D)*C*(~1*~(B*A))+D*C*(~1*~(B*A)))"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111100001110000),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg2_b31|PWM3/dir_reg  (
    .a({\PWM3/pnumr [31],\PWM3/n24 }),
    .b({pnum3[31],\PWM3/n25_neg_lutinv }),
    .c({pnum3[32],dir_pad[3]}),
    .clk(clk100m),
    .d({pwm_start_stop[19],\PWM3/pnumr [31]}),
    .e({open_n5948,pwm_start_stop[19]}),
    .q({\PWM3/pnumr[31]_keep ,\PWM3/dir_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg2_b5|PWM3/reg3_b5  (
    .a({\PWM3/pnumr [5],_al_u1945_o}),
    .b({pnum3[32],\PWM3/n24 }),
    .c({pnum3[5],pnumcnt3[5]}),
    .clk(clk100m),
    .d({pwm_start_stop[19],\PWM3/pnumr [5]}),
    .e({open_n5970,pwm_start_stop[19]}),
    .q({\PWM3/pnumr[5]_keep ,\PWM3/RemaTxNum[5]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg2_b6|PWM3/reg3_b6  (
    .a({\PWM3/pnumr [6],_al_u1943_o}),
    .b({pnum3[32],\PWM3/n24 }),
    .c({pnum3[6],pnumcnt3[6]}),
    .clk(clk100m),
    .d({pwm_start_stop[19],\PWM3/pnumr [6]}),
    .e({open_n5992,pwm_start_stop[19]}),
    .q({\PWM3/pnumr[6]_keep ,\PWM3/RemaTxNum[6]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg2_b9|PWM3/reg3_b9  (
    .a({\PWM3/pnumr [9],_al_u1937_o}),
    .b({pnum3[32],\PWM3/n24 }),
    .c({pnum3[9],pnumcnt3[9]}),
    .clk(clk100m),
    .d({pwm_start_stop[19],\PWM3/pnumr [9]}),
    .e({open_n6014,pwm_start_stop[19]}),
    .q({\PWM3/pnumr[9]_keep ,\PWM3/RemaTxNum[9]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg3_b1  (
    .a({_al_u1981_o,_al_u1981_o}),
    .b({\PWM3/n24 ,\PWM3/n24 }),
    .c({pnumcnt3[1],pnumcnt3[1]}),
    .clk(clk100m),
    .d({\PWM3/pnumr [1],\PWM3/pnumr [1]}),
    .mi({open_n6046,pwm_start_stop[19]}),
    .q({open_n6053,\PWM3/RemaTxNum[1]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg3_b10  (
    .a({_al_u1979_o,_al_u1979_o}),
    .b({\PWM3/n24 ,\PWM3/n24 }),
    .c({pnumcnt3[10],pnumcnt3[10]}),
    .clk(clk100m),
    .d({\PWM3/pnumr [10],\PWM3/pnumr [10]}),
    .mi({open_n6065,pwm_start_stop[19]}),
    .q({open_n6072,\PWM3/RemaTxNum[10]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg3_b13  (
    .a({_al_u1973_o,_al_u1973_o}),
    .b({\PWM3/n24 ,\PWM3/n24 }),
    .c({pnumcnt3[13],pnumcnt3[13]}),
    .clk(clk100m),
    .d({\PWM3/pnumr [13],\PWM3/pnumr [13]}),
    .mi({open_n6084,pwm_start_stop[19]}),
    .q({open_n6091,\PWM3/RemaTxNum[13]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg3_b14  (
    .a({_al_u1971_o,_al_u1971_o}),
    .b({\PWM3/n24 ,\PWM3/n24 }),
    .c({pnumcnt3[14],pnumcnt3[14]}),
    .clk(clk100m),
    .d({\PWM3/pnumr [14],\PWM3/pnumr [14]}),
    .mi({open_n6103,pwm_start_stop[19]}),
    .q({open_n6110,\PWM3/RemaTxNum[14]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg3_b17  (
    .a({_al_u1965_o,_al_u1965_o}),
    .b({\PWM3/n24 ,\PWM3/n24 }),
    .c({pnumcnt3[17],pnumcnt3[17]}),
    .clk(clk100m),
    .d({\PWM3/pnumr [17],\PWM3/pnumr [17]}),
    .mi({open_n6122,pwm_start_stop[19]}),
    .q({open_n6129,\PWM3/RemaTxNum[17]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg3_b18  (
    .a({_al_u1963_o,_al_u1963_o}),
    .b({\PWM3/n24 ,\PWM3/n24 }),
    .c({pnumcnt3[18],pnumcnt3[18]}),
    .clk(clk100m),
    .d({\PWM3/pnumr [18],\PWM3/pnumr [18]}),
    .mi({open_n6141,pwm_start_stop[19]}),
    .q({open_n6148,\PWM3/RemaTxNum[18]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg3_b20  (
    .a({_al_u1957_o,_al_u1957_o}),
    .b({\PWM3/n24 ,\PWM3/n24 }),
    .c({pnumcnt3[20],pnumcnt3[20]}),
    .clk(clk100m),
    .d({\PWM3/pnumr [20],\PWM3/pnumr [20]}),
    .mi({open_n6160,pwm_start_stop[19]}),
    .q({open_n6167,\PWM3/RemaTxNum[20]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg3_b21  (
    .a({_al_u1955_o,_al_u1955_o}),
    .b({\PWM3/n24 ,\PWM3/n24 }),
    .c({pnumcnt3[21],pnumcnt3[21]}),
    .clk(clk100m),
    .d({\PWM3/pnumr [21],\PWM3/pnumr [21]}),
    .mi({open_n6179,pwm_start_stop[19]}),
    .q({open_n6186,\PWM3/RemaTxNum[21]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg3_b3  (
    .a({_al_u1949_o,_al_u1949_o}),
    .b({\PWM3/n24 ,\PWM3/n24 }),
    .c({pnumcnt3[3],pnumcnt3[3]}),
    .clk(clk100m),
    .d({\PWM3/pnumr [3],\PWM3/pnumr [3]}),
    .mi({open_n6198,pwm_start_stop[19]}),
    .q({open_n6205,\PWM3/RemaTxNum[3]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg3_b4  (
    .a({_al_u1947_o,_al_u1947_o}),
    .b({\PWM3/n24 ,\PWM3/n24 }),
    .c({pnumcnt3[4],pnumcnt3[4]}),
    .clk(clk100m),
    .d({\PWM3/pnumr [4],\PWM3/pnumr [4]}),
    .mi({open_n6217,pwm_start_stop[19]}),
    .q({open_n6224,\PWM3/RemaTxNum[4]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg3_b7  (
    .a({_al_u1941_o,_al_u1941_o}),
    .b({\PWM3/n24 ,\PWM3/n24 }),
    .c({pnumcnt3[7],pnumcnt3[7]}),
    .clk(clk100m),
    .d({\PWM3/pnumr [7],\PWM3/pnumr [7]}),
    .mi({open_n6236,pwm_start_stop[19]}),
    .q({open_n6243,\PWM3/RemaTxNum[7]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/reg3_b8  (
    .a({_al_u1939_o,_al_u1939_o}),
    .b({\PWM3/n24 ,\PWM3/n24 }),
    .c({pnumcnt3[8],pnumcnt3[8]}),
    .clk(clk100m),
    .d({\PWM3/pnumr [8],\PWM3/pnumr [8]}),
    .mi({open_n6255,pwm_start_stop[19]}),
    .q({open_n6262,\PWM3/RemaTxNum[8]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_LSLICE #(
    //.MACRO("PWM3/sub0/ucin_al_u3384"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM3/sub0/u11_al_u3387  (
    .a({\PWM3/FreCnt [13],\PWM3/FreCnt [11]}),
    .b({\PWM3/FreCnt [14],\PWM3/FreCnt [12]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM3/sub0/c11 ),
    .f({\PWM3/n12 [13],\PWM3/n12 [11]}),
    .fco(\PWM3/sub0/c15 ),
    .fx({\PWM3/n12 [14],\PWM3/n12 [12]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM3/sub0/ucin_al_u3384"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM3/sub0/u15_al_u3388  (
    .a({\PWM3/FreCnt [17],\PWM3/FreCnt [15]}),
    .b({\PWM3/FreCnt [18],\PWM3/FreCnt [16]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM3/sub0/c15 ),
    .f({\PWM3/n12 [17],\PWM3/n12 [15]}),
    .fco(\PWM3/sub0/c19 ),
    .fx({\PWM3/n12 [18],\PWM3/n12 [16]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM3/sub0/ucin_al_u3384"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM3/sub0/u19_al_u3389  (
    .a({\PWM3/FreCnt [21],\PWM3/FreCnt [19]}),
    .b({\PWM3/FreCnt [22],\PWM3/FreCnt [20]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM3/sub0/c19 ),
    .f({\PWM3/n12 [21],\PWM3/n12 [19]}),
    .fco(\PWM3/sub0/c23 ),
    .fx({\PWM3/n12 [22],\PWM3/n12 [20]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM3/sub0/ucin_al_u3384"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM3/sub0/u23_al_u3390  (
    .a({\PWM3/FreCnt [25],\PWM3/FreCnt [23]}),
    .b({\PWM3/FreCnt [26],\PWM3/FreCnt [24]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM3/sub0/c23 ),
    .f({\PWM3/n12 [25],\PWM3/n12 [23]}),
    .fx({\PWM3/n12 [26],\PWM3/n12 [24]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM3/sub0/ucin_al_u3384"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM3/sub0/u3_al_u3385  (
    .a({\PWM3/FreCnt [5],\PWM3/FreCnt [3]}),
    .b({\PWM3/FreCnt [6],\PWM3/FreCnt [4]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM3/sub0/c3 ),
    .f({\PWM3/n12 [5],\PWM3/n12 [3]}),
    .fco(\PWM3/sub0/c7 ),
    .fx({\PWM3/n12 [6],\PWM3/n12 [4]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM3/sub0/ucin_al_u3384"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM3/sub0/u7_al_u3386  (
    .a({\PWM3/FreCnt [9],\PWM3/FreCnt [7]}),
    .b({\PWM3/FreCnt [10],\PWM3/FreCnt [8]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM3/sub0/c7 ),
    .f({\PWM3/n12 [9],\PWM3/n12 [7]}),
    .fco(\PWM3/sub0/c11 ),
    .fx({\PWM3/n12 [10],\PWM3/n12 [8]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM3/sub0/ucin_al_u3384"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'h0005),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM3/sub0/ucin_al_u3384  (
    .a({\PWM3/FreCnt [1],1'b0}),
    .b({\PWM3/FreCnt [2],\PWM3/FreCnt [0]}),
    .c(2'b11),
    .ce(\U_AHB/n10 ),
    .clk(clk100m),
    .d(2'b01),
    .e(2'b01),
    .mi({open_n6373,\U_AHB/h2h_hwdata [2]}),
    .f({\PWM3/n12 [1],open_n6386}),
    .fco(\PWM3/sub0/c3 ),
    .fx({\PWM3/n12 [2],\PWM3/n12 [0]}),
    .q({open_n6387,freq3[2]}));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM3/sub1/u0|PWM3/sub1/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("SUB_CARRY"),
    .INIT_LUT0(16'b0000000000000101),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM3/sub1/u0|PWM3/sub1/ucin  (
    .a({pnumcnt3[0],1'b0}),
    .b({1'b1,open_n6388}),
    .f({\PWM3/n26 [0],open_n6408}),
    .fco(\PWM3/sub1/c1 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM3/sub1/u0|PWM3/sub1/ucin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM3/sub1/u10|PWM3/sub1/u9  (
    .a(pnumcnt3[10:9]),
    .b(2'b00),
    .fci(\PWM3/sub1/c9 ),
    .f(\PWM3/n26 [10:9]),
    .fco(\PWM3/sub1/c11 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM3/sub1/u0|PWM3/sub1/ucin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM3/sub1/u12|PWM3/sub1/u11  (
    .a(pnumcnt3[12:11]),
    .b(2'b00),
    .fci(\PWM3/sub1/c11 ),
    .f(\PWM3/n26 [12:11]),
    .fco(\PWM3/sub1/c13 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM3/sub1/u0|PWM3/sub1/ucin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM3/sub1/u14|PWM3/sub1/u13  (
    .a(pnumcnt3[14:13]),
    .b(2'b00),
    .fci(\PWM3/sub1/c13 ),
    .f(\PWM3/n26 [14:13]),
    .fco(\PWM3/sub1/c15 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM3/sub1/u0|PWM3/sub1/ucin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM3/sub1/u16|PWM3/sub1/u15  (
    .a(pnumcnt3[16:15]),
    .b(2'b00),
    .fci(\PWM3/sub1/c15 ),
    .f(\PWM3/n26 [16:15]),
    .fco(\PWM3/sub1/c17 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM3/sub1/u0|PWM3/sub1/ucin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM3/sub1/u18|PWM3/sub1/u17  (
    .a(pnumcnt3[18:17]),
    .b(2'b00),
    .fci(\PWM3/sub1/c17 ),
    .f(\PWM3/n26 [18:17]),
    .fco(\PWM3/sub1/c19 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM3/sub1/u0|PWM3/sub1/ucin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM3/sub1/u20|PWM3/sub1/u19  (
    .a(pnumcnt3[20:19]),
    .b(2'b00),
    .fci(\PWM3/sub1/c19 ),
    .f(\PWM3/n26 [20:19]),
    .fco(\PWM3/sub1/c21 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM3/sub1/u0|PWM3/sub1/ucin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM3/sub1/u22|PWM3/sub1/u21  (
    .a(pnumcnt3[22:21]),
    .b(2'b00),
    .fci(\PWM3/sub1/c21 ),
    .f(\PWM3/n26 [22:21]),
    .fco(\PWM3/sub1/c23 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM3/sub1/u0|PWM3/sub1/ucin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM3/sub1/u23_al_u3471  (
    .a({open_n6567,pnumcnt3[23]}),
    .b({open_n6568,1'b0}),
    .fci(\PWM3/sub1/c23 ),
    .f({open_n6587,\PWM3/n26 [23]}));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM3/sub1/u0|PWM3/sub1/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM3/sub1/u2|PWM3/sub1/u1  (
    .a(pnumcnt3[2:1]),
    .b(2'b00),
    .fci(\PWM3/sub1/c1 ),
    .f(\PWM3/n26 [2:1]),
    .fco(\PWM3/sub1/c3 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM3/sub1/u0|PWM3/sub1/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM3/sub1/u4|PWM3/sub1/u3  (
    .a(pnumcnt3[4:3]),
    .b(2'b00),
    .fci(\PWM3/sub1/c3 ),
    .f(\PWM3/n26 [4:3]),
    .fco(\PWM3/sub1/c5 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM3/sub1/u0|PWM3/sub1/ucin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM3/sub1/u6|PWM3/sub1/u5  (
    .a(pnumcnt3[6:5]),
    .b(2'b00),
    .fci(\PWM3/sub1/c5 ),
    .f(\PWM3/n26 [6:5]),
    .fco(\PWM3/sub1/c7 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM3/sub1/u0|PWM3/sub1/ucin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM3/sub1/u8|PWM3/sub1/u7  (
    .a(pnumcnt3[8:7]),
    .b(2'b00),
    .fci(\PWM3/sub1/c7 ),
    .f(\PWM3/n26 [8:7]),
    .fco(\PWM3/sub1/c9 ));
  // src/OnePWM.v(26)
  // src/OnePWM.v(26)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*~(~D*B*~A))"),
    //.LUTF1("(C*~(~D*B*~A))"),
    //.LUTG0("(C*~(~D*B*~A))"),
    //.LUTG1("(C*~(~D*B*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000010110000),
    .INIT_LUTF1(16'b1111000010110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \PWM4/State_reg|PWMB/State_reg  (
    .a({_al_u3019_o,_al_u3040_o}),
    .b({\PWM4/n0_lutinv ,\PWMB/n0_lutinv }),
    .c({_al_u3020_o,_al_u3041_o}),
    .clk(clk100m),
    .d({pwm_start_stop[20],pwm_start_stop[27]}),
    .sr(rstn),
    .q({pwm_state_read[4],pwm_state_read[11]}));  // src/OnePWM.v(26)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[0]  (
    .i(\PWM4/RemaTxNum[0]_keep ),
    .o(pnumcnt4[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[10]  (
    .i(\PWM4/RemaTxNum[10]_keep ),
    .o(pnumcnt4[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[11]  (
    .i(\PWM4/RemaTxNum[11]_keep ),
    .o(pnumcnt4[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[12]  (
    .i(\PWM4/RemaTxNum[12]_keep ),
    .o(pnumcnt4[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[13]  (
    .i(\PWM4/RemaTxNum[13]_keep ),
    .o(pnumcnt4[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[14]  (
    .i(\PWM4/RemaTxNum[14]_keep ),
    .o(pnumcnt4[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[15]  (
    .i(\PWM4/RemaTxNum[15]_keep ),
    .o(pnumcnt4[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[16]  (
    .i(\PWM4/RemaTxNum[16]_keep ),
    .o(pnumcnt4[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[17]  (
    .i(\PWM4/RemaTxNum[17]_keep ),
    .o(pnumcnt4[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[18]  (
    .i(\PWM4/RemaTxNum[18]_keep ),
    .o(pnumcnt4[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[19]  (
    .i(\PWM4/RemaTxNum[19]_keep ),
    .o(pnumcnt4[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[1]  (
    .i(\PWM4/RemaTxNum[1]_keep ),
    .o(pnumcnt4[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[20]  (
    .i(\PWM4/RemaTxNum[20]_keep ),
    .o(pnumcnt4[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[21]  (
    .i(\PWM4/RemaTxNum[21]_keep ),
    .o(pnumcnt4[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[22]  (
    .i(\PWM4/RemaTxNum[22]_keep ),
    .o(pnumcnt4[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[23]  (
    .i(\PWM4/RemaTxNum[23]_keep ),
    .o(pnumcnt4[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[2]  (
    .i(\PWM4/RemaTxNum[2]_keep ),
    .o(pnumcnt4[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[3]  (
    .i(\PWM4/RemaTxNum[3]_keep ),
    .o(pnumcnt4[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[4]  (
    .i(\PWM4/RemaTxNum[4]_keep ),
    .o(pnumcnt4[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[5]  (
    .i(\PWM4/RemaTxNum[5]_keep ),
    .o(pnumcnt4[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[6]  (
    .i(\PWM4/RemaTxNum[6]_keep ),
    .o(pnumcnt4[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[7]  (
    .i(\PWM4/RemaTxNum[7]_keep ),
    .o(pnumcnt4[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[8]  (
    .i(\PWM4/RemaTxNum[8]_keep ),
    .o(pnumcnt4[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[9]  (
    .i(\PWM4/RemaTxNum[9]_keep ),
    .o(pnumcnt4[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_dir  (
    .i(\PWM4/dir_keep ),
    .o(dir_pad[4]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[0]  (
    .i(\PWM4/pnumr[0]_keep ),
    .o(\PWM4/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[10]  (
    .i(\PWM4/pnumr[10]_keep ),
    .o(\PWM4/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[11]  (
    .i(\PWM4/pnumr[11]_keep ),
    .o(\PWM4/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[12]  (
    .i(\PWM4/pnumr[12]_keep ),
    .o(\PWM4/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[13]  (
    .i(\PWM4/pnumr[13]_keep ),
    .o(\PWM4/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[14]  (
    .i(\PWM4/pnumr[14]_keep ),
    .o(\PWM4/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[15]  (
    .i(\PWM4/pnumr[15]_keep ),
    .o(\PWM4/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[16]  (
    .i(\PWM4/pnumr[16]_keep ),
    .o(\PWM4/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[17]  (
    .i(\PWM4/pnumr[17]_keep ),
    .o(\PWM4/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[18]  (
    .i(\PWM4/pnumr[18]_keep ),
    .o(\PWM4/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[19]  (
    .i(\PWM4/pnumr[19]_keep ),
    .o(\PWM4/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[1]  (
    .i(\PWM4/pnumr[1]_keep ),
    .o(\PWM4/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[20]  (
    .i(\PWM4/pnumr[20]_keep ),
    .o(\PWM4/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[21]  (
    .i(\PWM4/pnumr[21]_keep ),
    .o(\PWM4/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[22]  (
    .i(\PWM4/pnumr[22]_keep ),
    .o(\PWM4/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[23]  (
    .i(\PWM4/pnumr[23]_keep ),
    .o(\PWM4/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[24]  (
    .i(\PWM4/pnumr[24]_keep ),
    .o(\PWM4/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[25]  (
    .i(\PWM4/pnumr[25]_keep ),
    .o(\PWM4/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[26]  (
    .i(\PWM4/pnumr[26]_keep ),
    .o(\PWM4/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[27]  (
    .i(\PWM4/pnumr[27]_keep ),
    .o(\PWM4/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[28]  (
    .i(\PWM4/pnumr[28]_keep ),
    .o(\PWM4/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[29]  (
    .i(\PWM4/pnumr[29]_keep ),
    .o(\PWM4/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[2]  (
    .i(\PWM4/pnumr[2]_keep ),
    .o(\PWM4/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[30]  (
    .i(\PWM4/pnumr[30]_keep ),
    .o(\PWM4/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[31]  (
    .i(\PWM4/pnumr[31]_keep ),
    .o(\PWM4/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[3]  (
    .i(\PWM4/pnumr[3]_keep ),
    .o(\PWM4/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[4]  (
    .i(\PWM4/pnumr[4]_keep ),
    .o(\PWM4/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[5]  (
    .i(\PWM4/pnumr[5]_keep ),
    .o(\PWM4/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[6]  (
    .i(\PWM4/pnumr[6]_keep ),
    .o(\PWM4/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[7]  (
    .i(\PWM4/pnumr[7]_keep ),
    .o(\PWM4/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[8]  (
    .i(\PWM4/pnumr[8]_keep ),
    .o(\PWM4/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[9]  (
    .i(\PWM4/pnumr[9]_keep ),
    .o(\PWM4/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pwm  (
    .i(\PWM4/pwm_keep ),
    .o(pwm_pad[4]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_stopreq  (
    .i(\PWM4/stopreq_keep ),
    .o(\PWM4/stopreq ));  // src/OnePWM.v(14)
  EF2_PHY_MSLICE #(
    //.LUT0("(D*~(C)*~((~0*~(B*A)))+D*C*~((~0*~(B*A)))+~(D)*C*(~0*~(B*A))+D*C*(~0*~(B*A)))"),
    //.LUT1("(D*~(C)*~((~1*~(B*A)))+D*C*~((~1*~(B*A)))+~(D)*C*(~1*~(B*A))+D*C*(~1*~(B*A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111100001110000),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/dir_reg  (
    .a({\PWM4/n24 ,\PWM4/n24 }),
    .b({\PWM4/n25_neg_lutinv ,\PWM4/n25_neg_lutinv }),
    .c({dir_pad[4],dir_pad[4]}),
    .clk(clk100m),
    .d({\PWM4/pnumr [31],\PWM4/pnumr [31]}),
    .mi({open_n6714,pwm_start_stop[20]}),
    .q({open_n6721,\PWM4/dir_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("~(~0*~(D*C*B*A))"),
    //.LUT1("~(~1*~(D*C*B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b1111111111111111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM4/pwm_reg  (
    .a({_al_u1435_o,_al_u1435_o}),
    .b({_al_u1441_o,_al_u1441_o}),
    .c({_al_u1443_o,_al_u1443_o}),
    .clk(clk100m),
    .d({_al_u1445_o,_al_u1445_o}),
    .mi({open_n6733,pwm_pad[4]}),
    .sr(\PWM4/u14_sel_is_1_o ),
    .q({open_n6739,\PWM4/pwm_keep }));  // src/OnePWM.v(45)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM4/reg0_b0|PWM4/reg0_b15  (
    .b({\PWM4/n12 [0],\PWM4/n12 [15]}),
    .c({freq4[0],freq4[15]}),
    .clk(clk100m),
    .d({\PWM4/n0_lutinv ,\PWM4/n0_lutinv }),
    .sr(\PWM4/n11 ),
    .q({\PWM4/FreCnt [0],\PWM4/FreCnt [15]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM4/reg0_b10|PWM4/reg0_b12  (
    .b({\PWM4/n12 [10],\PWM4/n12 [12]}),
    .c({freq4[10],freq4[12]}),
    .clk(clk100m),
    .d({\PWM4/n0_lutinv ,\PWM4/n0_lutinv }),
    .sr(\PWM4/n11 ),
    .q({\PWM4/FreCnt [10],\PWM4/FreCnt [12]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM4/reg0_b11|PWM4/reg0_b8  (
    .b({\PWM4/n12 [11],\PWM4/n12 [8]}),
    .c({freq4[11],freq4[8]}),
    .clk(clk100m),
    .d({\PWM4/n0_lutinv ,\PWM4/n0_lutinv }),
    .sr(\PWM4/n11 ),
    .q({\PWM4/FreCnt [11],\PWM4/FreCnt [8]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM4/reg0_b13|PWM4/reg0_b7  (
    .b({\PWM4/n12 [13],\PWM4/n12 [7]}),
    .c({freq4[13],freq4[7]}),
    .clk(clk100m),
    .d({\PWM4/n0_lutinv ,\PWM4/n0_lutinv }),
    .sr(\PWM4/n11 ),
    .q({\PWM4/FreCnt [13],\PWM4/FreCnt [7]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM4/reg0_b14|PWM4/reg0_b6  (
    .b({\PWM4/n12 [14],\PWM4/n12 [6]}),
    .c({freq4[14],freq4[6]}),
    .clk(clk100m),
    .d({\PWM4/n0_lutinv ,\PWM4/n0_lutinv }),
    .sr(\PWM4/n11 ),
    .q({\PWM4/FreCnt [14],\PWM4/FreCnt [6]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM4/reg0_b16|PWM4/reg0_b5  (
    .b({\PWM4/n12 [16],\PWM4/n12 [5]}),
    .c({freq4[16],freq4[5]}),
    .clk(clk100m),
    .d({\PWM4/n0_lutinv ,\PWM4/n0_lutinv }),
    .sr(\PWM4/n11 ),
    .q({\PWM4/FreCnt [16],\PWM4/FreCnt [5]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM4/reg0_b17|PWM4/reg0_b3  (
    .b({\PWM4/n12 [17],\PWM4/n12 [3]}),
    .c({freq4[17],freq4[3]}),
    .clk(clk100m),
    .d({\PWM4/n0_lutinv ,\PWM4/n0_lutinv }),
    .sr(\PWM4/n11 ),
    .q({\PWM4/FreCnt [17],\PWM4/FreCnt [3]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM4/reg0_b18|PWM4/reg0_b25  (
    .b({\PWM4/n12 [18],\PWM4/n12 [25]}),
    .c({freq4[18],freq4[25]}),
    .clk(clk100m),
    .d({\PWM4/n0_lutinv ,\PWM4/n0_lutinv }),
    .sr(\PWM4/n11 ),
    .q({\PWM4/FreCnt [18],\PWM4/FreCnt [25]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM4/reg0_b19|PWM4/reg0_b23  (
    .b({\PWM4/n12 [19],\PWM4/n12 [23]}),
    .c({freq4[19],freq4[23]}),
    .clk(clk100m),
    .d({\PWM4/n0_lutinv ,\PWM4/n0_lutinv }),
    .sr(\PWM4/n11 ),
    .q({\PWM4/FreCnt [19],\PWM4/FreCnt [23]}));  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM4/reg0_b2  (
    .b({open_n6934,\PWM4/n12 [2]}),
    .c({open_n6935,freq4[2]}),
    .clk(clk100m),
    .d({open_n6937,\PWM4/n0_lutinv }),
    .sr(\PWM4/n11 ),
    .q({open_n6955,\PWM4/FreCnt [2]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM4/reg0_b20|PWM4/reg0_b1  (
    .b({\PWM4/n12 [20],\PWM4/n12 [1]}),
    .c({freq4[20],freq4[1]}),
    .clk(clk100m),
    .d({\PWM4/n0_lutinv ,\PWM4/n0_lutinv }),
    .sr(\PWM4/n11 ),
    .q({\PWM4/FreCnt [20],\PWM4/FreCnt [1]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM4/reg0_b21|PWM4/reg0_b9  (
    .b({\PWM4/n12 [21],\PWM4/n12 [9]}),
    .c({freq4[21],freq4[9]}),
    .clk(clk100m),
    .d({\PWM4/n0_lutinv ,\PWM4/n0_lutinv }),
    .sr(\PWM4/n11 ),
    .q({\PWM4/FreCnt [21],\PWM4/FreCnt [9]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM4/reg0_b22|PWM4/reg0_b4  (
    .b({\PWM4/n12 [22],\PWM4/n12 [4]}),
    .c({freq4[22],freq4[4]}),
    .clk(clk100m),
    .d({\PWM4/n0_lutinv ,\PWM4/n0_lutinv }),
    .sr(\PWM4/n11 ),
    .q({\PWM4/FreCnt [22],\PWM4/FreCnt [4]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM4/reg0_b24|PWM4/reg0_b26  (
    .b({\PWM4/n12 [24],\PWM4/n12 [26]}),
    .c({freq4[24],freq4[26]}),
    .clk(clk100m),
    .d({\PWM4/n0_lutinv ,\PWM4/n0_lutinv }),
    .sr(\PWM4/n11 ),
    .q({\PWM4/FreCnt [24],\PWM4/FreCnt [26]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~A*~(0@C)*~(D*~B))"),
    //.LUTF1("(A*~(0@C)*~(D@B))"),
    //.LUTG0("(~A*~(1@C)*~(D*~B))"),
    //.LUTG1("(A*~(1@C)*~(D@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010000000101),
    .INIT_LUTF1(16'b0000100000000010),
    .INIT_LUTG0(16'b0100000001010000),
    .INIT_LUTG1(16'b1000000000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg1_b10|PWM4/reg1_b1  (
    .a({_al_u1444_o,_al_u2089_o}),
    .b(\PWM4/FreCnt [1:0]),
    .c(\PWM4/FreCnt [10:9]),
    .ce(\PWM4/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM4/FreCntr [1],\PWM4/FreCntr [1]}),
    .e({\PWM4/FreCntr [10],\PWM4/FreCntr [10]}),
    .mi({freq4[10],freq4[1]}),
    .f({_al_u1445_o,_al_u2090_o}),
    .q({\PWM4/FreCntr [10],\PWM4/FreCntr [1]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(~0*C)*~(D*~B))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(A*~(~1*C)*~(D*~B))"),
    //.LUTG1("(~C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000001010),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1000100010101010),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg1_b14|PWM4/reg1_b4  (
    .a({open_n7064,_al_u2084_o}),
    .b({open_n7065,\PWM4/FreCnt [13]}),
    .c({\PWM4/FreCntr [14],\PWM4/FreCnt [3]}),
    .ce(\PWM4/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM4/FreCnt [13],\PWM4/FreCntr [14]}),
    .e({open_n7066,\PWM4/FreCntr [4]}),
    .mi({freq4[14],freq4[4]}),
    .f({_al_u2087_o,_al_u2085_o}),
    .q({\PWM4/FreCntr [14],\PWM4/FreCntr [4]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg1_b15|PWM4/reg1_b5  (
    .a({\PWM4/FreCnt [14],_al_u1430_o}),
    .b({\PWM4/FreCnt [4],\PWM4/FreCnt [18]}),
    .c({\PWM4/FreCntr [15],\PWM4/FreCnt [5]}),
    .ce(\PWM4/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM4/FreCntr [5],\PWM4/FreCntr [18]}),
    .e({open_n7083,\PWM4/FreCntr [5]}),
    .mi({freq4[15],freq4[5]}),
    .f({_al_u2076_o,_al_u1431_o}),
    .q({\PWM4/FreCntr [15],\PWM4/FreCntr [5]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~(~D*B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111010100110001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg1_b16|PWM4/reg1_b0  (
    .a({\PWM4/FreCnt [15],open_n7100}),
    .b({\PWM4/FreCnt [7],open_n7101}),
    .c({\PWM4/FreCntr [16],\PWM4/n11 }),
    .ce(\PWM4/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM4/FreCntr [8],\PWM4/n0_lutinv }),
    .mi({freq4[16],freq4[0]}),
    .f({_al_u2084_o,\PWM4/mux3_b0_sel_is_3_o }),
    .q({\PWM4/FreCntr [16],\PWM4/FreCntr [0]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(B*A*~(D@C))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(B*A*~(D@C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b1000000000001000),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg1_b17|PWM4/reg1_b8  (
    .a({_al_u2068_o,_al_u1432_o}),
    .b({_al_u2069_o,\PWM4/FreCnt [17]}),
    .c({\PWM4/FreCnt [16],\PWM4/FreCnt [8]}),
    .ce(\PWM4/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM4/FreCntr [17],\PWM4/FreCntr [17]}),
    .e({open_n7116,\PWM4/FreCntr [8]}),
    .mi({freq4[17],freq4[8]}),
    .f({_al_u2070_o,_al_u1433_o}),
    .q({\PWM4/FreCntr [17],\PWM4/FreCntr [8]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~D*B)*~(C*~A))"),
    //.LUT1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111100100011),
    .INIT_LUT1(16'b1000010000100001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg1_b19|PWM4/reg1_b20  (
    .a({\PWM4/FreCnt [18],\PWM4/FreCnt [15]}),
    .b({\PWM4/FreCnt [2],\PWM4/FreCnt [19]}),
    .c({\PWM4/FreCntr [19],\PWM4/FreCntr [16]}),
    .ce(\PWM4/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM4/FreCntr [3],\PWM4/FreCntr [20]}),
    .mi({freq4[19],freq4[20]}),
    .f({_al_u2078_o,_al_u2073_o}),
    .q({\PWM4/FreCntr [19],\PWM4/FreCntr [20]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(D@B)*~(C@A))"),
    //.LUT1("(D*~(C@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000010000100001),
    .INIT_LUT1(16'b1100001100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg1_b21|PWM4/reg1_b3  (
    .a({open_n7147,\PWM4/FreCnt [2]}),
    .b({\PWM4/FreCnt [20],\PWM4/FreCnt [3]}),
    .c({\PWM4/FreCntr [21],\PWM4/FreCntr [2]}),
    .ce(\PWM4/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({_al_u2076_o,\PWM4/FreCntr [3]}),
    .mi({freq4[21],freq4[3]}),
    .f({_al_u2077_o,_al_u1444_o}),
    .q({\PWM4/FreCntr [21],\PWM4/FreCntr [3]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg1_b23|PWM4/reg1_b22  (
    .a({\PWM4/FreCnt [22],_al_u2078_o}),
    .b({\PWM4/FreCnt [23],\PWM4/FreCnt [21]}),
    .c({\PWM4/FreCntr [22],\PWM4/FreCnt [22]}),
    .ce(\PWM4/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d(\PWM4/FreCntr [23:22]),
    .e({open_n7162,\PWM4/FreCntr [23]}),
    .mi(freq4[23:22]),
    .f({_al_u1432_o,_al_u2079_o}),
    .q(\PWM4/FreCntr [23:22]));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*~C)*~(D@B))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(A*~(1*~C)*~(D@B))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000100000100010),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg1_b24|PWM4/reg1_b12  (
    .a({\PWM4/FreCnt [0],_al_u2085_o}),
    .b({\PWM4/FreCnt [24],\PWM4/FreCnt [11]}),
    .c({\PWM4/FreCntr [0],\PWM4/FreCnt [23]}),
    .ce(\PWM4/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM4/FreCntr [24],\PWM4/FreCntr [12]}),
    .e({open_n7179,\PWM4/FreCntr [24]}),
    .mi({freq4[24],freq4[12]}),
    .f({_al_u1438_o,_al_u2086_o}),
    .q({\PWM4/FreCntr [24],\PWM4/FreCntr [12]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*~C)*~(D*~B))"),
    //.LUTF1("(A*~(~0*C)*~(~D*B))"),
    //.LUTG0("(A*~(1*~C)*~(D*~B))"),
    //.LUTG1("(A*~(~1*C)*~(~D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000100010101010),
    .INIT_LUTF1(16'b0000101000000010),
    .INIT_LUTG0(16'b1000000010100000),
    .INIT_LUTG1(16'b1010101000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg1_b26|PWM4/reg1_b6  (
    .a({_al_u2067_o,_al_u2071_o}),
    .b({\PWM4/FreCnt [25],\PWM4/FreCnt [5]}),
    .c({\PWM4/FreCnt [5],\PWM4/FreCnt [7]}),
    .ce(\PWM4/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM4/FreCntr [26],\PWM4/FreCntr [6]}),
    .e({\PWM4/FreCntr [6],\PWM4/FreCntr [8]}),
    .mi({freq4[26],freq4[6]}),
    .f({_al_u2068_o,_al_u2072_o}),
    .q({\PWM4/FreCntr [26],\PWM4/FreCntr [6]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*~C)*~(~D*B))"),
    //.LUTF1("(~(~D*B)*~(C*~A))"),
    //.LUTG0("(A*~(1*~C)*~(~D*B))"),
    //.LUTG1("(~(~D*B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101000100010),
    .INIT_LUTF1(16'b1010111100100011),
    .INIT_LUTG0(16'b1010000000100000),
    .INIT_LUTG1(16'b1010111100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg1_b2|PWM4/reg1_b18  (
    .a({\PWM4/FreCnt [1],_al_u2080_o}),
    .b({\PWM4/FreCnt [23],\PWM4/FreCnt [17]}),
    .c({\PWM4/FreCntr [2],\PWM4/FreCnt [3]}),
    .ce(\PWM4/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM4/FreCntr [24],\PWM4/FreCntr [18]}),
    .e({open_n7212,\PWM4/FreCntr [4]}),
    .mi({freq4[2],freq4[18]}),
    .f({_al_u2080_o,_al_u2081_o}),
    .q({\PWM4/FreCntr [2],\PWM4/FreCntr [18]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~A*~(~0*C)*~(D@B))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(~A*~(~1*C)*~(D@B))"),
    //.LUTG1("(C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010000000001),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0100010000010001),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg1_b7|PWM4/reg1_b25  (
    .a({open_n7229,_al_u2087_o}),
    .b({open_n7230,\PWM4/FreCnt [24]}),
    .c({\PWM4/FreCntr [7],\PWM4/FreCnt [6]}),
    .ce(\PWM4/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM4/FreCnt [6],\PWM4/FreCntr [25]}),
    .e({open_n7231,\PWM4/FreCntr [7]}),
    .mi({freq4[7],freq4[25]}),
    .f({_al_u2089_o,_al_u2088_o}),
    .q({\PWM4/FreCntr [7],\PWM4/FreCntr [25]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*~C)*~(D*~B))"),
    //.LUTF1("(~(~D*B)*~(~C*A))"),
    //.LUTG0("(A*~(1*~C)*~(D*~B))"),
    //.LUTG1("(~(~D*B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000100010101010),
    .INIT_LUTF1(16'b1111010100110001),
    .INIT_LUTG0(16'b1000000010100000),
    .INIT_LUTG1(16'b1111010100110001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg1_b9|PWM4/reg1_b13  (
    .a({\PWM4/FreCnt [0],_al_u2073_o}),
    .b({\PWM4/FreCnt [8],\PWM4/FreCnt [12]}),
    .c({\PWM4/FreCntr [1],\PWM4/FreCnt [8]}),
    .ce(\PWM4/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM4/FreCntr [9],\PWM4/FreCntr [13]}),
    .e({open_n7248,\PWM4/FreCntr [9]}),
    .mi({freq4[9],freq4[13]}),
    .f({_al_u2071_o,_al_u2074_o}),
    .q({\PWM4/FreCntr [9],\PWM4/FreCntr [13]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg2_b0|PWM4/reg3_b0  (
    .a({\PWM4/pnumr [0],_al_u2065_o}),
    .b({pnum4[0],\PWM4/n24 }),
    .c({pnum4[32],pnumcnt4[0]}),
    .clk(clk100m),
    .d({pwm_start_stop[20],\PWM4/pnumr [0]}),
    .e({open_n7266,pwm_start_stop[20]}),
    .q({\PWM4/pnumr[0]_keep ,\PWM4/RemaTxNum[0]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011100010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg2_b10|PWM4/reg2_b9  (
    .a(\PWM4/pnumr [10:9]),
    .b({pnum4[10],pnum4[32]}),
    .c({pnum4[32],pnum4[9]}),
    .clk(clk100m),
    .d({pwm_start_stop[20],pwm_start_stop[20]}),
    .q({\PWM4/pnumr[10]_keep ,\PWM4/pnumr[9]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011100010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011100010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg2_b11|PWM4/reg2_b8  (
    .a({\PWM4/pnumr [11],\PWM4/pnumr [8]}),
    .b({pnum4[11],pnum4[32]}),
    .c({pnum4[32],pnum4[8]}),
    .clk(clk100m),
    .d({pwm_start_stop[20],pwm_start_stop[20]}),
    .q({\PWM4/pnumr[11]_keep ,\PWM4/pnumr[8]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg2_b12|PWM4/reg3_b12  (
    .a({\PWM4/pnumr [12],_al_u2057_o}),
    .b({pnum4[12],\PWM4/n24 }),
    .c({pnum4[32],pnumcnt4[12]}),
    .clk(clk100m),
    .d({pwm_start_stop[20],\PWM4/pnumr [12]}),
    .e({open_n7330,pwm_start_stop[20]}),
    .q({\PWM4/pnumr[12]_keep ,\PWM4/RemaTxNum[12]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg2_b13|PWM4/reg3_b13  (
    .a({\PWM4/pnumr [13],_al_u2055_o}),
    .b({pnum4[13],\PWM4/n24 }),
    .c({pnum4[32],pnumcnt4[13]}),
    .clk(clk100m),
    .d({pwm_start_stop[20],\PWM4/pnumr [13]}),
    .e({open_n7352,pwm_start_stop[20]}),
    .q({\PWM4/pnumr[13]_keep ,\PWM4/RemaTxNum[13]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011100010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011100010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg2_b14|PWM4/reg2_b5  (
    .a({\PWM4/pnumr [14],\PWM4/pnumr [5]}),
    .b({pnum4[14],pnum4[32]}),
    .c({pnum4[32],pnum4[5]}),
    .clk(clk100m),
    .d({pwm_start_stop[20],pwm_start_stop[20]}),
    .q({\PWM4/pnumr[14]_keep ,\PWM4/pnumr[5]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011100010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg2_b15|PWM4/reg2_b4  (
    .a({\PWM4/pnumr [15],\PWM4/pnumr [4]}),
    .b({pnum4[15],pnum4[32]}),
    .c({pnum4[32],pnum4[4]}),
    .clk(clk100m),
    .d({pwm_start_stop[20],pwm_start_stop[20]}),
    .q({\PWM4/pnumr[15]_keep ,\PWM4/pnumr[4]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg2_b16|PWM4/reg3_b16  (
    .a({\PWM4/pnumr [16],_al_u2049_o}),
    .b({pnum4[16],\PWM4/n24 }),
    .c({pnum4[32],pnumcnt4[16]}),
    .clk(clk100m),
    .d({pwm_start_stop[20],\PWM4/pnumr [16]}),
    .e({open_n7416,pwm_start_stop[20]}),
    .q({\PWM4/pnumr[16]_keep ,\PWM4/RemaTxNum[16]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg2_b17|PWM4/reg3_b17  (
    .a({\PWM4/pnumr [17],_al_u2047_o}),
    .b({pnum4[17],\PWM4/n24 }),
    .c({pnum4[32],pnumcnt4[17]}),
    .clk(clk100m),
    .d({pwm_start_stop[20],\PWM4/pnumr [17]}),
    .e({open_n7438,pwm_start_stop[20]}),
    .q({\PWM4/pnumr[17]_keep ,\PWM4/RemaTxNum[17]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg2_b18|PWM4/reg2_b22  (
    .a({\PWM4/pnumr [18],\PWM4/pnumr [22]}),
    .b({pnum4[18],pnum4[22]}),
    .c({pnum4[32],pnum4[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[20],pwm_start_stop[20]}),
    .q({\PWM4/pnumr[18]_keep ,\PWM4/pnumr[22]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg2_b19|PWM4/reg2_b21  (
    .a({\PWM4/pnumr [19],\PWM4/pnumr [21]}),
    .b({pnum4[19],pnum4[21]}),
    .c({pnum4[32],pnum4[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[20],pwm_start_stop[20]}),
    .q({\PWM4/pnumr[19]_keep ,\PWM4/pnumr[21]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg2_b1|PWM4/reg3_b1  (
    .a({\PWM4/pnumr [1],_al_u2063_o}),
    .b({pnum4[1],\PWM4/n24 }),
    .c({pnum4[32],pnumcnt4[1]}),
    .clk(clk100m),
    .d({pwm_start_stop[20],\PWM4/pnumr [1]}),
    .e({open_n7502,pwm_start_stop[20]}),
    .q({\PWM4/pnumr[1]_keep ,\PWM4/RemaTxNum[1]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg2_b20|PWM4/reg3_b20  (
    .a({\PWM4/pnumr [20],_al_u2039_o}),
    .b({pnum4[20],\PWM4/n24 }),
    .c({pnum4[32],pnumcnt4[20]}),
    .clk(clk100m),
    .d({pwm_start_stop[20],\PWM4/pnumr [20]}),
    .e({open_n7524,pwm_start_stop[20]}),
    .q({\PWM4/pnumr[20]_keep ,\PWM4/RemaTxNum[20]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg2_b23|PWM4/reg3_b23  (
    .a({\PWM4/pnumr [23],_al_u2033_o}),
    .b({pnum4[23],\PWM4/n24 }),
    .c({pnum4[32],pnumcnt4[23]}),
    .clk(clk100m),
    .d({pwm_start_stop[20],\PWM4/pnumr [23]}),
    .e({open_n7546,pwm_start_stop[20]}),
    .q({\PWM4/pnumr[23]_keep ,\PWM4/RemaTxNum[23]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg2_b24|PWM4/reg2_b31  (
    .a({\PWM4/pnumr [24],\PWM4/pnumr [31]}),
    .b({pnum4[24],pnum4[31]}),
    .c({pnum4[32],pnum4[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[20],pwm_start_stop[20]}),
    .q({\PWM4/pnumr[24]_keep ,\PWM4/pnumr[31]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg2_b25|PWM4/reg2_b30  (
    .a({\PWM4/pnumr [25],\PWM4/pnumr [30]}),
    .b({pnum4[25],pnum4[30]}),
    .c({pnum4[32],pnum4[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[20],pwm_start_stop[20]}),
    .q({\PWM4/pnumr[25]_keep ,\PWM4/pnumr[30]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg2_b26|PWM4/reg2_b29  (
    .a({\PWM4/pnumr [26],\PWM4/pnumr [29]}),
    .b({pnum4[26],pnum4[29]}),
    .c({pnum4[32],pnum4[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[20],pwm_start_stop[20]}),
    .q({\PWM4/pnumr[26]_keep ,\PWM4/pnumr[29]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg2_b27|PWM4/reg2_b28  (
    .a({\PWM4/pnumr [27],\PWM4/pnumr [28]}),
    .b({pnum4[27],pnum4[28]}),
    .c({pnum4[32],pnum4[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[20],pwm_start_stop[20]}),
    .q({\PWM4/pnumr[27]_keep ,\PWM4/pnumr[28]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg2_b2|PWM4/reg3_b2  (
    .a({\PWM4/pnumr [2],_al_u2041_o}),
    .b({pnum4[2],\PWM4/n24 }),
    .c({pnum4[32],pnumcnt4[2]}),
    .clk(clk100m),
    .d({pwm_start_stop[20],\PWM4/pnumr [2]}),
    .e({open_n7648,pwm_start_stop[20]}),
    .q({\PWM4/pnumr[2]_keep ,\PWM4/RemaTxNum[2]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg2_b3|PWM4/reg3_b3  (
    .a({\PWM4/pnumr [3],_al_u2031_o}),
    .b({pnum4[3],\PWM4/n24 }),
    .c({pnum4[32],pnumcnt4[3]}),
    .clk(clk100m),
    .d({pwm_start_stop[20],\PWM4/pnumr [3]}),
    .e({open_n7670,pwm_start_stop[20]}),
    .q({\PWM4/pnumr[3]_keep ,\PWM4/RemaTxNum[3]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg2_b6|PWM4/reg3_b6  (
    .a({\PWM4/pnumr [6],_al_u2025_o}),
    .b({pnum4[32],\PWM4/n24 }),
    .c({pnum4[6],pnumcnt4[6]}),
    .clk(clk100m),
    .d({pwm_start_stop[20],\PWM4/pnumr [6]}),
    .e({open_n7692,pwm_start_stop[20]}),
    .q({\PWM4/pnumr[6]_keep ,\PWM4/RemaTxNum[6]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg2_b7|PWM4/reg3_b7  (
    .a({\PWM4/pnumr [7],_al_u2023_o}),
    .b({pnum4[32],\PWM4/n24 }),
    .c({pnum4[7],pnumcnt4[7]}),
    .clk(clk100m),
    .d({pwm_start_stop[20],\PWM4/pnumr [7]}),
    .e({open_n7714,pwm_start_stop[20]}),
    .q({\PWM4/pnumr[7]_keep ,\PWM4/RemaTxNum[7]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg3_b10  (
    .a({_al_u2061_o,_al_u2061_o}),
    .b({\PWM4/n24 ,\PWM4/n24 }),
    .c({pnumcnt4[10],pnumcnt4[10]}),
    .clk(clk100m),
    .d({\PWM4/pnumr [10],\PWM4/pnumr [10]}),
    .mi({open_n7746,pwm_start_stop[20]}),
    .q({open_n7753,\PWM4/RemaTxNum[10]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg3_b11  (
    .a({_al_u2059_o,_al_u2059_o}),
    .b({\PWM4/n24 ,\PWM4/n24 }),
    .c({pnumcnt4[11],pnumcnt4[11]}),
    .clk(clk100m),
    .d({\PWM4/pnumr [11],\PWM4/pnumr [11]}),
    .mi({open_n7765,pwm_start_stop[20]}),
    .q({open_n7772,\PWM4/RemaTxNum[11]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg3_b14  (
    .a({_al_u2053_o,_al_u2053_o}),
    .b({\PWM4/n24 ,\PWM4/n24 }),
    .c({pnumcnt4[14],pnumcnt4[14]}),
    .clk(clk100m),
    .d({\PWM4/pnumr [14],\PWM4/pnumr [14]}),
    .mi({open_n7784,pwm_start_stop[20]}),
    .q({open_n7791,\PWM4/RemaTxNum[14]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg3_b15  (
    .a({_al_u2051_o,_al_u2051_o}),
    .b({\PWM4/n24 ,\PWM4/n24 }),
    .c({pnumcnt4[15],pnumcnt4[15]}),
    .clk(clk100m),
    .d({\PWM4/pnumr [15],\PWM4/pnumr [15]}),
    .mi({open_n7803,pwm_start_stop[20]}),
    .q({open_n7810,\PWM4/RemaTxNum[15]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg3_b18  (
    .a({_al_u2045_o,_al_u2045_o}),
    .b({\PWM4/n24 ,\PWM4/n24 }),
    .c({pnumcnt4[18],pnumcnt4[18]}),
    .clk(clk100m),
    .d({\PWM4/pnumr [18],\PWM4/pnumr [18]}),
    .mi({open_n7822,pwm_start_stop[20]}),
    .q({open_n7829,\PWM4/RemaTxNum[18]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg3_b19  (
    .a({_al_u2043_o,_al_u2043_o}),
    .b({\PWM4/n24 ,\PWM4/n24 }),
    .c({pnumcnt4[19],pnumcnt4[19]}),
    .clk(clk100m),
    .d({\PWM4/pnumr [19],\PWM4/pnumr [19]}),
    .mi({open_n7841,pwm_start_stop[20]}),
    .q({open_n7848,\PWM4/RemaTxNum[19]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg3_b21  (
    .a({_al_u2037_o,_al_u2037_o}),
    .b({\PWM4/n24 ,\PWM4/n24 }),
    .c({pnumcnt4[21],pnumcnt4[21]}),
    .clk(clk100m),
    .d({\PWM4/pnumr [21],\PWM4/pnumr [21]}),
    .mi({open_n7860,pwm_start_stop[20]}),
    .q({open_n7867,\PWM4/RemaTxNum[21]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg3_b22  (
    .a({_al_u2035_o,_al_u2035_o}),
    .b({\PWM4/n24 ,\PWM4/n24 }),
    .c({pnumcnt4[22],pnumcnt4[22]}),
    .clk(clk100m),
    .d({\PWM4/pnumr [22],\PWM4/pnumr [22]}),
    .mi({open_n7879,pwm_start_stop[20]}),
    .q({open_n7886,\PWM4/RemaTxNum[22]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg3_b4  (
    .a({_al_u2029_o,_al_u2029_o}),
    .b({\PWM4/n24 ,\PWM4/n24 }),
    .c({pnumcnt4[4],pnumcnt4[4]}),
    .clk(clk100m),
    .d({\PWM4/pnumr [4],\PWM4/pnumr [4]}),
    .mi({open_n7898,pwm_start_stop[20]}),
    .q({open_n7905,\PWM4/RemaTxNum[4]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg3_b5  (
    .a({_al_u2027_o,_al_u2027_o}),
    .b({\PWM4/n24 ,\PWM4/n24 }),
    .c({pnumcnt4[5],pnumcnt4[5]}),
    .clk(clk100m),
    .d({\PWM4/pnumr [5],\PWM4/pnumr [5]}),
    .mi({open_n7917,pwm_start_stop[20]}),
    .q({open_n7924,\PWM4/RemaTxNum[5]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg3_b8  (
    .a({_al_u2021_o,_al_u2021_o}),
    .b({\PWM4/n24 ,\PWM4/n24 }),
    .c({pnumcnt4[8],pnumcnt4[8]}),
    .clk(clk100m),
    .d({\PWM4/pnumr [8],\PWM4/pnumr [8]}),
    .mi({open_n7936,pwm_start_stop[20]}),
    .q({open_n7943,\PWM4/RemaTxNum[8]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/reg3_b9  (
    .a({_al_u2019_o,_al_u2019_o}),
    .b({\PWM4/n24 ,\PWM4/n24 }),
    .c({pnumcnt4[9],pnumcnt4[9]}),
    .clk(clk100m),
    .d({\PWM4/pnumr [9],\PWM4/pnumr [9]}),
    .mi({open_n7955,pwm_start_stop[20]}),
    .q({open_n7962,\PWM4/RemaTxNum[9]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_LSLICE #(
    //.MACRO("PWM4/sub0/ucin_al_u3391"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM4/sub0/u11_al_u3394  (
    .a({\PWM4/FreCnt [13],\PWM4/FreCnt [11]}),
    .b({\PWM4/FreCnt [14],\PWM4/FreCnt [12]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM4/sub0/c11 ),
    .f({\PWM4/n12 [13],\PWM4/n12 [11]}),
    .fco(\PWM4/sub0/c15 ),
    .fx({\PWM4/n12 [14],\PWM4/n12 [12]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM4/sub0/ucin_al_u3391"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM4/sub0/u15_al_u3395  (
    .a({\PWM4/FreCnt [17],\PWM4/FreCnt [15]}),
    .b({\PWM4/FreCnt [18],\PWM4/FreCnt [16]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM4/sub0/c15 ),
    .f({\PWM4/n12 [17],\PWM4/n12 [15]}),
    .fco(\PWM4/sub0/c19 ),
    .fx({\PWM4/n12 [18],\PWM4/n12 [16]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM4/sub0/ucin_al_u3391"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM4/sub0/u19_al_u3396  (
    .a({\PWM4/FreCnt [21],\PWM4/FreCnt [19]}),
    .b({\PWM4/FreCnt [22],\PWM4/FreCnt [20]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM4/sub0/c19 ),
    .f({\PWM4/n12 [21],\PWM4/n12 [19]}),
    .fco(\PWM4/sub0/c23 ),
    .fx({\PWM4/n12 [22],\PWM4/n12 [20]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM4/sub0/ucin_al_u3391"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM4/sub0/u23_al_u3397  (
    .a({\PWM4/FreCnt [25],\PWM4/FreCnt [23]}),
    .b({\PWM4/FreCnt [26],\PWM4/FreCnt [24]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM4/sub0/c23 ),
    .f({\PWM4/n12 [25],\PWM4/n12 [23]}),
    .fx({\PWM4/n12 [26],\PWM4/n12 [24]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM4/sub0/ucin_al_u3391"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM4/sub0/u3_al_u3392  (
    .a({\PWM4/FreCnt [5],\PWM4/FreCnt [3]}),
    .b({\PWM4/FreCnt [6],\PWM4/FreCnt [4]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM4/sub0/c3 ),
    .f({\PWM4/n12 [5],\PWM4/n12 [3]}),
    .fco(\PWM4/sub0/c7 ),
    .fx({\PWM4/n12 [6],\PWM4/n12 [4]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM4/sub0/ucin_al_u3391"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM4/sub0/u7_al_u3393  (
    .a({\PWM4/FreCnt [9],\PWM4/FreCnt [7]}),
    .b({\PWM4/FreCnt [10],\PWM4/FreCnt [8]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM4/sub0/c7 ),
    .f({\PWM4/n12 [9],\PWM4/n12 [7]}),
    .fco(\PWM4/sub0/c11 ),
    .fx({\PWM4/n12 [10],\PWM4/n12 [8]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM4/sub0/ucin_al_u3391"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'h0005),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM4/sub0/ucin_al_u3391  (
    .a({\PWM4/FreCnt [1],1'b0}),
    .b({\PWM4/FreCnt [2],\PWM4/FreCnt [0]}),
    .c(2'b11),
    .ce(\U_AHB/n12 ),
    .clk(clk100m),
    .d(2'b01),
    .e(2'b01),
    .mi({open_n8073,\U_AHB/h2h_hwdata [2]}),
    .f({\PWM4/n12 [1],open_n8086}),
    .fco(\PWM4/sub0/c3 ),
    .fx({\PWM4/n12 [2],\PWM4/n12 [0]}),
    .q({open_n8087,freq4[2]}));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM4/sub1/u0|PWM4/sub1/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("SUB_CARRY"),
    .INIT_LUT0(16'b0000000000000101),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM4/sub1/u0|PWM4/sub1/ucin  (
    .a({pnumcnt4[0],1'b0}),
    .b({1'b1,open_n8088}),
    .f({\PWM4/n26 [0],open_n8108}),
    .fco(\PWM4/sub1/c1 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM4/sub1/u0|PWM4/sub1/ucin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM4/sub1/u10|PWM4/sub1/u9  (
    .a(pnumcnt4[10:9]),
    .b(2'b00),
    .fci(\PWM4/sub1/c9 ),
    .f(\PWM4/n26 [10:9]),
    .fco(\PWM4/sub1/c11 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM4/sub1/u0|PWM4/sub1/ucin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM4/sub1/u12|PWM4/sub1/u11  (
    .a(pnumcnt4[12:11]),
    .b(2'b00),
    .fci(\PWM4/sub1/c11 ),
    .f(\PWM4/n26 [12:11]),
    .fco(\PWM4/sub1/c13 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM4/sub1/u0|PWM4/sub1/ucin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM4/sub1/u14|PWM4/sub1/u13  (
    .a(pnumcnt4[14:13]),
    .b(2'b00),
    .fci(\PWM4/sub1/c13 ),
    .f(\PWM4/n26 [14:13]),
    .fco(\PWM4/sub1/c15 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM4/sub1/u0|PWM4/sub1/ucin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM4/sub1/u16|PWM4/sub1/u15  (
    .a(pnumcnt4[16:15]),
    .b(2'b00),
    .fci(\PWM4/sub1/c15 ),
    .f(\PWM4/n26 [16:15]),
    .fco(\PWM4/sub1/c17 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM4/sub1/u0|PWM4/sub1/ucin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM4/sub1/u18|PWM4/sub1/u17  (
    .a(pnumcnt4[18:17]),
    .b(2'b00),
    .fci(\PWM4/sub1/c17 ),
    .f(\PWM4/n26 [18:17]),
    .fco(\PWM4/sub1/c19 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM4/sub1/u0|PWM4/sub1/ucin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM4/sub1/u20|PWM4/sub1/u19  (
    .a(pnumcnt4[20:19]),
    .b(2'b00),
    .fci(\PWM4/sub1/c19 ),
    .f(\PWM4/n26 [20:19]),
    .fco(\PWM4/sub1/c21 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM4/sub1/u0|PWM4/sub1/ucin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM4/sub1/u22|PWM4/sub1/u21  (
    .a(pnumcnt4[22:21]),
    .b(2'b00),
    .fci(\PWM4/sub1/c21 ),
    .f(\PWM4/n26 [22:21]),
    .fco(\PWM4/sub1/c23 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM4/sub1/u0|PWM4/sub1/ucin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM4/sub1/u23_al_u3472  (
    .a({open_n8267,pnumcnt4[23]}),
    .b({open_n8268,1'b0}),
    .fci(\PWM4/sub1/c23 ),
    .f({open_n8287,\PWM4/n26 [23]}));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM4/sub1/u0|PWM4/sub1/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM4/sub1/u2|PWM4/sub1/u1  (
    .a(pnumcnt4[2:1]),
    .b(2'b00),
    .fci(\PWM4/sub1/c1 ),
    .f(\PWM4/n26 [2:1]),
    .fco(\PWM4/sub1/c3 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM4/sub1/u0|PWM4/sub1/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM4/sub1/u4|PWM4/sub1/u3  (
    .a(pnumcnt4[4:3]),
    .b(2'b00),
    .fci(\PWM4/sub1/c3 ),
    .f(\PWM4/n26 [4:3]),
    .fco(\PWM4/sub1/c5 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM4/sub1/u0|PWM4/sub1/ucin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM4/sub1/u6|PWM4/sub1/u5  (
    .a(pnumcnt4[6:5]),
    .b(2'b00),
    .fci(\PWM4/sub1/c5 ),
    .f(\PWM4/n26 [6:5]),
    .fco(\PWM4/sub1/c7 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM4/sub1/u0|PWM4/sub1/ucin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM4/sub1/u8|PWM4/sub1/u7  (
    .a(pnumcnt4[8:7]),
    .b(2'b00),
    .fci(\PWM4/sub1/c7 ),
    .f(\PWM4/n26 [8:7]),
    .fco(\PWM4/sub1/c9 ));
  // src/OnePWM.v(26)
  // src/OnePWM.v(26)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*~(~D*B*~A))"),
    //.LUTF1("(C*~(~D*B*~A))"),
    //.LUTG0("(C*~(~D*B*~A))"),
    //.LUTG1("(C*~(~D*B*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000010110000),
    .INIT_LUTF1(16'b1111000010110000),
    .INIT_LUTG0(16'b1111000010110000),
    .INIT_LUTG1(16'b1111000010110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \PWM5/State_reg|PWMA/State_reg  (
    .a({_al_u3022_o,_al_u3037_o}),
    .b({\PWM5/n0_lutinv ,\PWMA/n0_lutinv }),
    .c({_al_u3023_o,_al_u3038_o}),
    .clk(clk100m),
    .d({pwm_start_stop[21],pwm_start_stop[26]}),
    .sr(rstn),
    .q({pwm_state_read[5],pwm_state_read[10]}));  // src/OnePWM.v(26)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[0]  (
    .i(\PWM5/RemaTxNum[0]_keep ),
    .o(pnumcnt5[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[10]  (
    .i(\PWM5/RemaTxNum[10]_keep ),
    .o(pnumcnt5[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[11]  (
    .i(\PWM5/RemaTxNum[11]_keep ),
    .o(pnumcnt5[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[12]  (
    .i(\PWM5/RemaTxNum[12]_keep ),
    .o(pnumcnt5[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[13]  (
    .i(\PWM5/RemaTxNum[13]_keep ),
    .o(pnumcnt5[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[14]  (
    .i(\PWM5/RemaTxNum[14]_keep ),
    .o(pnumcnt5[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[15]  (
    .i(\PWM5/RemaTxNum[15]_keep ),
    .o(pnumcnt5[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[16]  (
    .i(\PWM5/RemaTxNum[16]_keep ),
    .o(pnumcnt5[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[17]  (
    .i(\PWM5/RemaTxNum[17]_keep ),
    .o(pnumcnt5[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[18]  (
    .i(\PWM5/RemaTxNum[18]_keep ),
    .o(pnumcnt5[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[19]  (
    .i(\PWM5/RemaTxNum[19]_keep ),
    .o(pnumcnt5[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[1]  (
    .i(\PWM5/RemaTxNum[1]_keep ),
    .o(pnumcnt5[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[20]  (
    .i(\PWM5/RemaTxNum[20]_keep ),
    .o(pnumcnt5[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[21]  (
    .i(\PWM5/RemaTxNum[21]_keep ),
    .o(pnumcnt5[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[22]  (
    .i(\PWM5/RemaTxNum[22]_keep ),
    .o(pnumcnt5[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[23]  (
    .i(\PWM5/RemaTxNum[23]_keep ),
    .o(pnumcnt5[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[2]  (
    .i(\PWM5/RemaTxNum[2]_keep ),
    .o(pnumcnt5[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[3]  (
    .i(\PWM5/RemaTxNum[3]_keep ),
    .o(pnumcnt5[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[4]  (
    .i(\PWM5/RemaTxNum[4]_keep ),
    .o(pnumcnt5[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[5]  (
    .i(\PWM5/RemaTxNum[5]_keep ),
    .o(pnumcnt5[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[6]  (
    .i(\PWM5/RemaTxNum[6]_keep ),
    .o(pnumcnt5[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[7]  (
    .i(\PWM5/RemaTxNum[7]_keep ),
    .o(pnumcnt5[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[8]  (
    .i(\PWM5/RemaTxNum[8]_keep ),
    .o(pnumcnt5[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[9]  (
    .i(\PWM5/RemaTxNum[9]_keep ),
    .o(pnumcnt5[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_dir  (
    .i(\PWM5/dir_keep ),
    .o(dir_pad[5]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[0]  (
    .i(\PWM5/pnumr[0]_keep ),
    .o(\PWM5/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[10]  (
    .i(\PWM5/pnumr[10]_keep ),
    .o(\PWM5/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[11]  (
    .i(\PWM5/pnumr[11]_keep ),
    .o(\PWM5/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[12]  (
    .i(\PWM5/pnumr[12]_keep ),
    .o(\PWM5/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[13]  (
    .i(\PWM5/pnumr[13]_keep ),
    .o(\PWM5/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[14]  (
    .i(\PWM5/pnumr[14]_keep ),
    .o(\PWM5/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[15]  (
    .i(\PWM5/pnumr[15]_keep ),
    .o(\PWM5/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[16]  (
    .i(\PWM5/pnumr[16]_keep ),
    .o(\PWM5/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[17]  (
    .i(\PWM5/pnumr[17]_keep ),
    .o(\PWM5/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[18]  (
    .i(\PWM5/pnumr[18]_keep ),
    .o(\PWM5/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[19]  (
    .i(\PWM5/pnumr[19]_keep ),
    .o(\PWM5/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[1]  (
    .i(\PWM5/pnumr[1]_keep ),
    .o(\PWM5/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[20]  (
    .i(\PWM5/pnumr[20]_keep ),
    .o(\PWM5/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[21]  (
    .i(\PWM5/pnumr[21]_keep ),
    .o(\PWM5/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[22]  (
    .i(\PWM5/pnumr[22]_keep ),
    .o(\PWM5/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[23]  (
    .i(\PWM5/pnumr[23]_keep ),
    .o(\PWM5/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[24]  (
    .i(\PWM5/pnumr[24]_keep ),
    .o(\PWM5/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[25]  (
    .i(\PWM5/pnumr[25]_keep ),
    .o(\PWM5/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[26]  (
    .i(\PWM5/pnumr[26]_keep ),
    .o(\PWM5/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[27]  (
    .i(\PWM5/pnumr[27]_keep ),
    .o(\PWM5/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[28]  (
    .i(\PWM5/pnumr[28]_keep ),
    .o(\PWM5/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[29]  (
    .i(\PWM5/pnumr[29]_keep ),
    .o(\PWM5/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[2]  (
    .i(\PWM5/pnumr[2]_keep ),
    .o(\PWM5/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[30]  (
    .i(\PWM5/pnumr[30]_keep ),
    .o(\PWM5/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[31]  (
    .i(\PWM5/pnumr[31]_keep ),
    .o(\PWM5/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[3]  (
    .i(\PWM5/pnumr[3]_keep ),
    .o(\PWM5/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[4]  (
    .i(\PWM5/pnumr[4]_keep ),
    .o(\PWM5/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[5]  (
    .i(\PWM5/pnumr[5]_keep ),
    .o(\PWM5/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[6]  (
    .i(\PWM5/pnumr[6]_keep ),
    .o(\PWM5/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[7]  (
    .i(\PWM5/pnumr[7]_keep ),
    .o(\PWM5/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[8]  (
    .i(\PWM5/pnumr[8]_keep ),
    .o(\PWM5/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[9]  (
    .i(\PWM5/pnumr[9]_keep ),
    .o(\PWM5/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pwm  (
    .i(\PWM5/pwm_keep ),
    .o(pwm_pad[5]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_stopreq  (
    .i(\PWM5/stopreq_keep ),
    .o(\PWM5/stopreq ));  // src/OnePWM.v(14)
  EF2_PHY_MSLICE #(
    //.LUT0("(D*~(C)*~((~0*~(B*A)))+D*C*~((~0*~(B*A)))+~(D)*C*(~0*~(B*A))+D*C*(~0*~(B*A)))"),
    //.LUT1("(D*~(C)*~((~1*~(B*A)))+D*C*~((~1*~(B*A)))+~(D)*C*(~1*~(B*A))+D*C*(~1*~(B*A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111100001110000),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/dir_reg  (
    .a({\PWM5/n24 ,\PWM5/n24 }),
    .b({\PWM5/n25_neg_lutinv ,\PWM5/n25_neg_lutinv }),
    .c({dir_pad[5],dir_pad[5]}),
    .clk(clk100m),
    .d({\PWM5/pnumr [31],\PWM5/pnumr [31]}),
    .mi({open_n8414,pwm_start_stop[21]}),
    .q({open_n8421,\PWM5/dir_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("~(~0*~(D*C*B*A))"),
    //.LUT1("~(~1*~(D*C*B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b1111111111111111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM5/pwm_reg  (
    .a({_al_u1452_o,_al_u1452_o}),
    .b({_al_u1458_o,_al_u1458_o}),
    .c({_al_u1460_o,_al_u1460_o}),
    .clk(clk100m),
    .d({_al_u1462_o,_al_u1462_o}),
    .mi({open_n8433,pwm_pad[5]}),
    .sr(\PWM5/u14_sel_is_1_o ),
    .q({open_n8439,\PWM5/pwm_keep }));  // src/OnePWM.v(45)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM5/reg0_b0|PWM5/reg0_b15  (
    .b({\PWM5/n12 [0],\PWM5/n12 [15]}),
    .c({freq5[0],freq5[15]}),
    .clk(clk100m),
    .d({\PWM5/n0_lutinv ,\PWM5/n0_lutinv }),
    .sr(\PWM5/n11 ),
    .q({\PWM5/FreCnt [0],\PWM5/FreCnt [15]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM5/reg0_b10|PWM5/reg0_b12  (
    .b({\PWM5/n12 [10],\PWM5/n12 [12]}),
    .c({freq5[10],freq5[12]}),
    .clk(clk100m),
    .d({\PWM5/n0_lutinv ,\PWM5/n0_lutinv }),
    .sr(\PWM5/n11 ),
    .q({\PWM5/FreCnt [10],\PWM5/FreCnt [12]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM5/reg0_b11|PWM5/reg0_b8  (
    .b({\PWM5/n12 [11],\PWM5/n12 [8]}),
    .c({freq5[11],freq5[8]}),
    .clk(clk100m),
    .d({\PWM5/n0_lutinv ,\PWM5/n0_lutinv }),
    .sr(\PWM5/n11 ),
    .q({\PWM5/FreCnt [11],\PWM5/FreCnt [8]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM5/reg0_b13|PWM5/reg0_b7  (
    .b({\PWM5/n12 [13],\PWM5/n12 [7]}),
    .c({freq5[13],freq5[7]}),
    .clk(clk100m),
    .d({\PWM5/n0_lutinv ,\PWM5/n0_lutinv }),
    .sr(\PWM5/n11 ),
    .q({\PWM5/FreCnt [13],\PWM5/FreCnt [7]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM5/reg0_b14|PWM5/reg0_b5  (
    .b({\PWM5/n12 [14],\PWM5/n12 [5]}),
    .c({freq5[14],freq5[5]}),
    .clk(clk100m),
    .d({\PWM5/n0_lutinv ,\PWM5/n0_lutinv }),
    .sr(\PWM5/n11 ),
    .q({\PWM5/FreCnt [14],\PWM5/FreCnt [5]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM5/reg0_b16|PWM5/reg0_b3  (
    .b({\PWM5/n12 [16],\PWM5/n12 [3]}),
    .c({freq5[16],freq5[3]}),
    .clk(clk100m),
    .d({\PWM5/n0_lutinv ,\PWM5/n0_lutinv }),
    .sr(\PWM5/n11 ),
    .q({\PWM5/FreCnt [16],\PWM5/FreCnt [3]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM5/reg0_b17|PWM5/reg0_b25  (
    .b({\PWM5/n12 [17],\PWM5/n12 [25]}),
    .c({freq5[17],freq5[25]}),
    .clk(clk100m),
    .d({\PWM5/n0_lutinv ,\PWM5/n0_lutinv }),
    .sr(\PWM5/n11 ),
    .q({\PWM5/FreCnt [17],\PWM5/FreCnt [25]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM5/reg0_b18|PWM5/reg0_b23  (
    .b({\PWM5/n12 [18],\PWM5/n12 [23]}),
    .c({freq5[18],freq5[23]}),
    .clk(clk100m),
    .d({\PWM5/n0_lutinv ,\PWM5/n0_lutinv }),
    .sr(\PWM5/n11 ),
    .q({\PWM5/FreCnt [18],\PWM5/FreCnt [23]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM5/reg0_b19|PWM5/reg0_b22  (
    .b({\PWM5/n12 [19],\PWM5/n12 [22]}),
    .c({freq5[19],freq5[22]}),
    .clk(clk100m),
    .d({\PWM5/n0_lutinv ,\PWM5/n0_lutinv }),
    .sr(\PWM5/n11 ),
    .q({\PWM5/FreCnt [19],\PWM5/FreCnt [22]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM5/reg0_b1|PWM5/reg0_b21  (
    .b({\PWM5/n12 [1],\PWM5/n12 [21]}),
    .c({freq5[1],freq5[21]}),
    .clk(clk100m),
    .d({\PWM5/n0_lutinv ,\PWM5/n0_lutinv }),
    .sr(\PWM5/n11 ),
    .q({\PWM5/FreCnt [1],\PWM5/FreCnt [21]}));  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM5/reg0_b2  (
    .b({open_n8666,\PWM5/n12 [2]}),
    .c({open_n8667,freq5[2]}),
    .clk(clk100m),
    .d({open_n8669,\PWM5/n0_lutinv }),
    .sr(\PWM5/n11 ),
    .q({open_n8687,\PWM5/FreCnt [2]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM5/reg0_b20|PWM5/reg0_b9  (
    .b({\PWM5/n12 [20],\PWM5/n12 [9]}),
    .c({freq5[20],freq5[9]}),
    .clk(clk100m),
    .d({\PWM5/n0_lutinv ,\PWM5/n0_lutinv }),
    .sr(\PWM5/n11 ),
    .q({\PWM5/FreCnt [20],\PWM5/FreCnt [9]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM5/reg0_b24|PWM5/reg0_b6  (
    .b({\PWM5/n12 [24],\PWM5/n12 [6]}),
    .c({freq5[24],freq5[6]}),
    .clk(clk100m),
    .d({\PWM5/n0_lutinv ,\PWM5/n0_lutinv }),
    .sr(\PWM5/n11 ),
    .q({\PWM5/FreCnt [24],\PWM5/FreCnt [6]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM5/reg0_b26|PWM5/reg0_b4  (
    .b({\PWM5/n12 [26],\PWM5/n12 [4]}),
    .c({freq5[26],freq5[4]}),
    .clk(clk100m),
    .d({\PWM5/n0_lutinv ,\PWM5/n0_lutinv }),
    .sr(\PWM5/n11 ),
    .q({\PWM5/FreCnt [26],\PWM5/FreCnt [4]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~(D*~B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1100010011110101),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg1_b11|PWM5/reg1_b0  (
    .a({\PWM5/FreCnt [10],open_n8756}),
    .b({\PWM5/FreCnt [5],open_n8757}),
    .c({\PWM5/FreCntr [11],\PWM5/n11 }),
    .ce(\PWM5/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM5/FreCntr [6],\PWM5/n0_lutinv }),
    .mi({freq5[11],freq5[0]}),
    .f({_al_u2167_o,\PWM5/mux3_b0_sel_is_3_o }),
    .q({\PWM5/FreCntr [11],\PWM5/FreCntr [0]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~D*B)*~(C*~A))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(~(~D*B)*~(C*~A))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010111100100011),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1010111100100011),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg1_b12|PWM5/reg1_b16  (
    .a({\PWM5/FreCnt [11],\PWM5/FreCnt [15]}),
    .b({\PWM5/FreCnt [6],\PWM5/FreCnt [19]}),
    .c({\PWM5/FreCntr [12],\PWM5/FreCntr [16]}),
    .ce(\PWM5/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM5/FreCntr [7],\PWM5/FreCntr [20]}),
    .mi({freq5[12],freq5[16]}),
    .f({_al_u2151_o,_al_u2169_o}),
    .q({\PWM5/FreCntr [12],\PWM5/FreCntr [16]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(~0*C)*~(~D*B))"),
    //.LUTF1("(A*~(0*~C)*~(D*~B))"),
    //.LUTG0("(A*~(~1*C)*~(~D*B))"),
    //.LUTG1("(A*~(1*~C)*~(D*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101000000010),
    .INIT_LUTF1(16'b1000100010101010),
    .INIT_LUTG0(16'b1010101000100010),
    .INIT_LUTG1(16'b1000000010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg1_b14|PWM5/reg1_b24  (
    .a({_al_u2171_o,_al_u2160_o}),
    .b({\PWM5/FreCnt [13],\PWM5/FreCnt [13]}),
    .c({\PWM5/FreCnt [17],\PWM5/FreCnt [23]}),
    .ce(\PWM5/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM5/FreCntr [14],\PWM5/FreCntr [14]}),
    .e({\PWM5/FreCntr [18],\PWM5/FreCntr [24]}),
    .mi({freq5[14],freq5[24]}),
    .f({_al_u2172_o,_al_u2161_o}),
    .q({\PWM5/FreCntr [14],\PWM5/FreCntr [24]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg1_b17|PWM5/reg1_b19  (
    .a({\PWM5/FreCnt [16],_al_u1455_o}),
    .b({\PWM5/FreCnt [18],\PWM5/FreCnt [13]}),
    .c({\PWM5/FreCntr [17],\PWM5/FreCnt [19]}),
    .ce(\PWM5/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM5/FreCntr [19],\PWM5/FreCntr [13]}),
    .e({open_n8806,\PWM5/FreCntr [19]}),
    .mi({freq5[17],freq5[19]}),
    .f({_al_u2162_o,_al_u1456_o}),
    .q({\PWM5/FreCntr [17],\PWM5/FreCntr [19]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~D*B)*~(C*~A))"),
    //.LUT1("(D*~(C@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111100100011),
    .INIT_LUT1(16'b1100001100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg1_b1|PWM5/reg1_b13  (
    .a({open_n8823,\PWM5/FreCnt [10]}),
    .b({\PWM5/FreCnt [0],\PWM5/FreCnt [12]}),
    .c({\PWM5/FreCntr [1],\PWM5/FreCntr [11]}),
    .ce(\PWM5/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({_al_u2151_o,\PWM5/FreCntr [13]}),
    .mi({freq5[1],freq5[13]}),
    .f({_al_u2152_o,_al_u2165_o}),
    .q({\PWM5/FreCntr [1],\PWM5/FreCntr [13]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~A*~(0*~C)*~(D@B))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(~A*~(1*~C)*~(D@B))"),
    //.LUTG1("(C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100010000010001),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0100000000010000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg1_b20|PWM5/reg1_b15  (
    .a({open_n8838,_al_u2155_o}),
    .b({open_n8839,\PWM5/FreCnt [14]}),
    .c({\PWM5/FreCntr [20],\PWM5/FreCnt [22]}),
    .ce(\PWM5/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM5/FreCnt [19],\PWM5/FreCntr [15]}),
    .e({open_n8840,\PWM5/FreCntr [23]}),
    .mi({freq5[20],freq5[15]}),
    .f({_al_u2155_o,_al_u2156_o}),
    .q({\PWM5/FreCntr [20],\PWM5/FreCntr [15]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D@C)*~(0@B))"),
    //.LUTF1("(C*B*A*~(0@D))"),
    //.LUTG0("(A*~(D@C)*~(1@B))"),
    //.LUTG1("(C*B*A*~(1@D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010000000000010),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b1000000000001000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg1_b21|PWM5/reg1_b10  (
    .a({_al_u1454_o,_al_u2162_o}),
    .b({_al_u1456_o,\PWM5/FreCnt [20]}),
    .c({_al_u1457_o,\PWM5/FreCnt [9]}),
    .ce(\PWM5/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM5/FreCnt [21],\PWM5/FreCntr [10]}),
    .e({\PWM5/FreCntr [21],\PWM5/FreCntr [21]}),
    .mi({freq5[21],freq5[10]}),
    .f({_al_u1458_o,_al_u2163_o}),
    .q({\PWM5/FreCntr [21],\PWM5/FreCntr [10]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(~0*C)*~(~D*B))"),
    //.LUTF1("(~(D*~B)*~(C*~A))"),
    //.LUTG0("(A*~(~1*C)*~(~D*B))"),
    //.LUTG1("(~(D*~B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101000000010),
    .INIT_LUTF1(16'b1000110010101111),
    .INIT_LUTG0(16'b1010101000100010),
    .INIT_LUTG1(16'b1000110010101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg1_b22|PWM5/reg1_b18  (
    .a({\PWM5/FreCnt [12],_al_u2153_o}),
    .b({\PWM5/FreCnt [21],\PWM5/FreCnt [17]}),
    .c({\PWM5/FreCntr [13],\PWM5/FreCnt [21]}),
    .ce(\PWM5/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM5/FreCntr [22],\PWM5/FreCntr [18]}),
    .e({open_n8873,\PWM5/FreCntr [22]}),
    .mi({freq5[22],freq5[18]}),
    .f({_al_u2158_o,_al_u2154_o}),
    .q({\PWM5/FreCntr [22],\PWM5/FreCntr [18]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(A*~(0@C)*~(D@B))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(A*~(1@C)*~(D@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b0000100000000010),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000000000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg1_b25|PWM5/reg1_b5  (
    .a({_al_u2149_o,_al_u1447_o}),
    .b({\PWM5/FreCnt [24],\PWM5/FreCnt [18]}),
    .c({\PWM5/FreCnt [4],\PWM5/FreCnt [5]}),
    .ce(\PWM5/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM5/FreCntr [25],\PWM5/FreCntr [18]}),
    .e({\PWM5/FreCntr [5],\PWM5/FreCntr [5]}),
    .mi({freq5[25],freq5[5]}),
    .f({_al_u2150_o,_al_u1448_o}),
    .q({\PWM5/FreCntr [25],\PWM5/FreCntr [5]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(~0*C)*~(D*~B))"),
    //.LUTF1("(A*~(0*~C)*~(~D*B))"),
    //.LUTG0("(A*~(~1*C)*~(D*~B))"),
    //.LUTG1("(A*~(1*~C)*~(~D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000001010),
    .INIT_LUTF1(16'b1010101000100010),
    .INIT_LUTG0(16'b1000100010101010),
    .INIT_LUTG1(16'b1010000000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg1_b26|PWM5/reg1_b4  (
    .a({_al_u2169_o,_al_u2165_o}),
    .b({\PWM5/FreCnt [25],\PWM5/FreCnt [25]}),
    .c({\PWM5/FreCnt [3],\PWM5/FreCnt [3]}),
    .ce(\PWM5/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM5/FreCntr [26],\PWM5/FreCntr [26]}),
    .e({\PWM5/FreCntr [4],\PWM5/FreCntr [4]}),
    .mi({freq5[26],freq5[4]}),
    .f({_al_u2170_o,_al_u2166_o}),
    .q({\PWM5/FreCntr [26],\PWM5/FreCntr [4]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~C*~(~D*B)*~(0@A))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(~C*~(~D*B)*~(1@A))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010100000001),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b0000101000000010),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg1_b3|PWM5/reg1_b23  (
    .a({\PWM5/FreCnt [2],\PWM5/FreCnt [2]}),
    .b({\PWM5/FreCnt [3],\PWM5/FreCnt [22]}),
    .c({\PWM5/FreCntr [2],\PWM5/FreCnt [26]}),
    .ce(\PWM5/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM5/FreCntr [3],\PWM5/FreCntr [23]}),
    .e({open_n8922,\PWM5/FreCntr [3]}),
    .mi({freq5[3],freq5[23]}),
    .f({_al_u1461_o,_al_u2149_o}),
    .q({\PWM5/FreCntr [3],\PWM5/FreCntr [23]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(D*~B)*~(C*~A))"),
    //.LUTF1("(~(~D*B)*~(~C*A))"),
    //.LUTG0("(~(D*~B)*~(C*~A))"),
    //.LUTG1("(~(~D*B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000110010101111),
    .INIT_LUTF1(16'b1111010100110001),
    .INIT_LUTG0(16'b1000110010101111),
    .INIT_LUTG1(16'b1111010100110001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg1_b6|PWM5/reg1_b8  (
    .a({\PWM5/FreCnt [5],\PWM5/FreCnt [7]}),
    .b({\PWM5/FreCnt [7],\PWM5/FreCnt [8]}),
    .c({\PWM5/FreCntr [6],\PWM5/FreCntr [8]}),
    .ce(\PWM5/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM5/FreCntr [8],\PWM5/FreCntr [9]}),
    .mi({freq5[6],freq5[8]}),
    .f({_al_u2160_o,_al_u2153_o}),
    .q({\PWM5/FreCntr [6],\PWM5/FreCntr [8]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(D*~B)*~(~C*A))"),
    //.LUT1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100010011110101),
    .INIT_LUT1(16'b1000010000100001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg1_b7|PWM5/reg1_b2  (
    .a({\PWM5/FreCnt [7],\PWM5/FreCnt [1]}),
    .b({\PWM5/FreCnt [9],\PWM5/FreCnt [23]}),
    .c({\PWM5/FreCntr [7],\PWM5/FreCntr [2]}),
    .ce(\PWM5/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM5/FreCntr [9],\PWM5/FreCntr [24]}),
    .mi({freq5[7],freq5[2]}),
    .f({_al_u1459_o,_al_u2171_o}),
    .q({\PWM5/FreCntr [7],\PWM5/FreCntr [2]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011100010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011100010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg2_b0|PWM5/reg2_b9  (
    .a({\PWM5/pnumr [0],\PWM5/pnumr [9]}),
    .b({pnum5[0],pnum5[32]}),
    .c({pnum5[32],pnum5[9]}),
    .clk(clk100m),
    .d({pwm_start_stop[21],pwm_start_stop[21]}),
    .q({\PWM5/pnumr[0]_keep ,\PWM5/pnumr[9]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg2_b10|PWM5/reg3_b10  (
    .a({\PWM5/pnumr [10],_al_u2143_o}),
    .b({pnum5[10],\PWM5/n24 }),
    .c({pnum5[32],pnumcnt5[10]}),
    .clk(clk100m),
    .d({pwm_start_stop[21],\PWM5/pnumr [10]}),
    .e({open_n8995,pwm_start_stop[21]}),
    .q({\PWM5/pnumr[10]_keep ,\PWM5/RemaTxNum[10]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011100010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg2_b11|PWM5/reg2_b6  (
    .a({\PWM5/pnumr [11],\PWM5/pnumr [6]}),
    .b({pnum5[11],pnum5[32]}),
    .c({pnum5[32],pnum5[6]}),
    .clk(clk100m),
    .d({pwm_start_stop[21],pwm_start_stop[21]}),
    .q({\PWM5/pnumr[11]_keep ,\PWM5/pnumr[6]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011100010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg2_b12|PWM5/reg2_b5  (
    .a({\PWM5/pnumr [12],\PWM5/pnumr [5]}),
    .b({pnum5[12],pnum5[32]}),
    .c({pnum5[32],pnum5[5]}),
    .clk(clk100m),
    .d({pwm_start_stop[21],pwm_start_stop[21]}),
    .q({\PWM5/pnumr[12]_keep ,\PWM5/pnumr[5]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg2_b13|PWM5/reg3_b13  (
    .a({\PWM5/pnumr [13],_al_u2137_o}),
    .b({pnum5[13],\PWM5/n24 }),
    .c({pnum5[32],pnumcnt5[13]}),
    .clk(clk100m),
    .d({pwm_start_stop[21],\PWM5/pnumr [13]}),
    .e({open_n9055,pwm_start_stop[21]}),
    .q({\PWM5/pnumr[13]_keep ,\PWM5/RemaTxNum[13]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg2_b14|PWM5/reg3_b14  (
    .a({\PWM5/pnumr [14],_al_u2135_o}),
    .b({pnum5[14],\PWM5/n24 }),
    .c({pnum5[32],pnumcnt5[14]}),
    .clk(clk100m),
    .d({pwm_start_stop[21],\PWM5/pnumr [14]}),
    .e({open_n9077,pwm_start_stop[21]}),
    .q({\PWM5/pnumr[14]_keep ,\PWM5/RemaTxNum[14]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg2_b15|PWM5/reg2_b23  (
    .a({\PWM5/pnumr [15],\PWM5/pnumr [23]}),
    .b({pnum5[15],pnum5[23]}),
    .c({pnum5[32],pnum5[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[21],pwm_start_stop[21]}),
    .q({\PWM5/pnumr[15]_keep ,\PWM5/pnumr[23]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg2_b16|PWM5/reg2_b22  (
    .a({\PWM5/pnumr [16],\PWM5/pnumr [22]}),
    .b({pnum5[16],pnum5[22]}),
    .c({pnum5[32],pnum5[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[21],pwm_start_stop[21]}),
    .q({\PWM5/pnumr[16]_keep ,\PWM5/pnumr[22]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg2_b17|PWM5/reg3_b17  (
    .a({\PWM5/pnumr [17],_al_u2129_o}),
    .b({pnum5[17],\PWM5/n24 }),
    .c({pnum5[32],pnumcnt5[17]}),
    .clk(clk100m),
    .d({pwm_start_stop[21],\PWM5/pnumr [17]}),
    .e({open_n9145,pwm_start_stop[21]}),
    .q({\PWM5/pnumr[17]_keep ,\PWM5/RemaTxNum[17]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg2_b18|PWM5/reg3_b18  (
    .a({\PWM5/pnumr [18],_al_u2127_o}),
    .b({pnum5[18],\PWM5/n24 }),
    .c({pnum5[32],pnumcnt5[18]}),
    .clk(clk100m),
    .d({pwm_start_stop[21],\PWM5/pnumr [18]}),
    .e({open_n9167,pwm_start_stop[21]}),
    .q({\PWM5/pnumr[18]_keep ,\PWM5/RemaTxNum[18]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg2_b19|PWM5/reg2_b2  (
    .a({\PWM5/pnumr [19],\PWM5/pnumr [2]}),
    .b({pnum5[19],pnum5[2]}),
    .c({pnum5[32],pnum5[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[21],pwm_start_stop[21]}),
    .q({\PWM5/pnumr[19]_keep ,\PWM5/pnumr[2]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg2_b1|PWM5/reg3_b1  (
    .a({\PWM5/pnumr [1],_al_u2145_o}),
    .b({pnum5[1],\PWM5/n24 }),
    .c({pnum5[32],pnumcnt5[1]}),
    .clk(clk100m),
    .d({pwm_start_stop[21],\PWM5/pnumr [1]}),
    .e({open_n9208,pwm_start_stop[21]}),
    .q({\PWM5/pnumr[1]_keep ,\PWM5/RemaTxNum[1]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg2_b20|PWM5/reg3_b20  (
    .a({\PWM5/pnumr [20],_al_u2121_o}),
    .b({pnum5[20],\PWM5/n24 }),
    .c({pnum5[32],pnumcnt5[20]}),
    .clk(clk100m),
    .d({pwm_start_stop[21],\PWM5/pnumr [20]}),
    .e({open_n9230,pwm_start_stop[21]}),
    .q({\PWM5/pnumr[20]_keep ,\PWM5/RemaTxNum[20]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg2_b21|PWM5/reg3_b21  (
    .a({\PWM5/pnumr [21],_al_u2119_o}),
    .b({pnum5[21],\PWM5/n24 }),
    .c({pnum5[32],pnumcnt5[21]}),
    .clk(clk100m),
    .d({pwm_start_stop[21],\PWM5/pnumr [21]}),
    .e({open_n9252,pwm_start_stop[21]}),
    .q({\PWM5/pnumr[21]_keep ,\PWM5/RemaTxNum[21]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg2_b24|PWM5/reg2_b31  (
    .a({\PWM5/pnumr [24],\PWM5/pnumr [31]}),
    .b({pnum5[24],pnum5[31]}),
    .c({pnum5[32],pnum5[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[21],pwm_start_stop[21]}),
    .q({\PWM5/pnumr[24]_keep ,\PWM5/pnumr[31]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg2_b25|PWM5/reg2_b30  (
    .a({\PWM5/pnumr [25],\PWM5/pnumr [30]}),
    .b({pnum5[25],pnum5[30]}),
    .c({pnum5[32],pnum5[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[21],pwm_start_stop[21]}),
    .q({\PWM5/pnumr[25]_keep ,\PWM5/pnumr[30]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg2_b26|PWM5/reg2_b29  (
    .a({\PWM5/pnumr [26],\PWM5/pnumr [29]}),
    .b({pnum5[26],pnum5[29]}),
    .c({pnum5[32],pnum5[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[21],pwm_start_stop[21]}),
    .q({\PWM5/pnumr[26]_keep ,\PWM5/pnumr[29]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg2_b27|PWM5/reg2_b28  (
    .a({\PWM5/pnumr [27],\PWM5/pnumr [28]}),
    .b({pnum5[27],pnum5[28]}),
    .c({pnum5[32],pnum5[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[21],pwm_start_stop[21]}),
    .q({\PWM5/pnumr[27]_keep ,\PWM5/pnumr[28]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg2_b3|PWM5/reg3_b3  (
    .a({\PWM5/pnumr [3],_al_u2113_o}),
    .b({pnum5[3],\PWM5/n24 }),
    .c({pnum5[32],pnumcnt5[3]}),
    .clk(clk100m),
    .d({pwm_start_stop[21],\PWM5/pnumr [3]}),
    .e({open_n9354,pwm_start_stop[21]}),
    .q({\PWM5/pnumr[3]_keep ,\PWM5/RemaTxNum[3]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg2_b4|PWM5/reg3_b4  (
    .a({\PWM5/pnumr [4],_al_u2111_o}),
    .b({pnum5[32],\PWM5/n24 }),
    .c({pnum5[4],pnumcnt5[4]}),
    .clk(clk100m),
    .d({pwm_start_stop[21],\PWM5/pnumr [4]}),
    .e({open_n9376,pwm_start_stop[21]}),
    .q({\PWM5/pnumr[4]_keep ,\PWM5/RemaTxNum[4]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg2_b7|PWM5/reg3_b7  (
    .a({\PWM5/pnumr [7],_al_u2105_o}),
    .b({pnum5[32],\PWM5/n24 }),
    .c({pnum5[7],pnumcnt5[7]}),
    .clk(clk100m),
    .d({pwm_start_stop[21],\PWM5/pnumr [7]}),
    .e({open_n9398,pwm_start_stop[21]}),
    .q({\PWM5/pnumr[7]_keep ,\PWM5/RemaTxNum[7]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg2_b8|PWM5/reg3_b8  (
    .a({\PWM5/pnumr [8],_al_u2103_o}),
    .b({pnum5[32],\PWM5/n24 }),
    .c({pnum5[8],pnumcnt5[8]}),
    .clk(clk100m),
    .d({pwm_start_stop[21],\PWM5/pnumr [8]}),
    .e({open_n9420,pwm_start_stop[21]}),
    .q({\PWM5/pnumr[8]_keep ,\PWM5/RemaTxNum[8]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg3_b0  (
    .a({_al_u2147_o,_al_u2147_o}),
    .b({\PWM5/n24 ,\PWM5/n24 }),
    .c({pnumcnt5[0],pnumcnt5[0]}),
    .clk(clk100m),
    .d({\PWM5/pnumr [0],\PWM5/pnumr [0]}),
    .mi({open_n9452,pwm_start_stop[21]}),
    .q({open_n9459,\PWM5/RemaTxNum[0]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg3_b11  (
    .a({_al_u2141_o,_al_u2141_o}),
    .b({\PWM5/n24 ,\PWM5/n24 }),
    .c({pnumcnt5[11],pnumcnt5[11]}),
    .clk(clk100m),
    .d({\PWM5/pnumr [11],\PWM5/pnumr [11]}),
    .mi({open_n9471,pwm_start_stop[21]}),
    .q({open_n9478,\PWM5/RemaTxNum[11]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg3_b12  (
    .a({_al_u2139_o,_al_u2139_o}),
    .b({\PWM5/n24 ,\PWM5/n24 }),
    .c({pnumcnt5[12],pnumcnt5[12]}),
    .clk(clk100m),
    .d({\PWM5/pnumr [12],\PWM5/pnumr [12]}),
    .mi({open_n9490,pwm_start_stop[21]}),
    .q({open_n9497,\PWM5/RemaTxNum[12]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg3_b15  (
    .a({_al_u2133_o,_al_u2133_o}),
    .b({\PWM5/n24 ,\PWM5/n24 }),
    .c({pnumcnt5[15],pnumcnt5[15]}),
    .clk(clk100m),
    .d({\PWM5/pnumr [15],\PWM5/pnumr [15]}),
    .mi({open_n9509,pwm_start_stop[21]}),
    .q({open_n9516,\PWM5/RemaTxNum[15]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg3_b16  (
    .a({_al_u2131_o,_al_u2131_o}),
    .b({\PWM5/n24 ,\PWM5/n24 }),
    .c({pnumcnt5[16],pnumcnt5[16]}),
    .clk(clk100m),
    .d({\PWM5/pnumr [16],\PWM5/pnumr [16]}),
    .mi({open_n9528,pwm_start_stop[21]}),
    .q({open_n9535,\PWM5/RemaTxNum[16]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg3_b19  (
    .a({_al_u2125_o,_al_u2125_o}),
    .b({\PWM5/n24 ,\PWM5/n24 }),
    .c({pnumcnt5[19],pnumcnt5[19]}),
    .clk(clk100m),
    .d({\PWM5/pnumr [19],\PWM5/pnumr [19]}),
    .mi({open_n9547,pwm_start_stop[21]}),
    .q({open_n9554,\PWM5/RemaTxNum[19]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg3_b2  (
    .a({_al_u2123_o,_al_u2123_o}),
    .b({\PWM5/n24 ,\PWM5/n24 }),
    .c({pnumcnt5[2],pnumcnt5[2]}),
    .clk(clk100m),
    .d({\PWM5/pnumr [2],\PWM5/pnumr [2]}),
    .mi({open_n9566,pwm_start_stop[21]}),
    .q({open_n9573,\PWM5/RemaTxNum[2]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg3_b22  (
    .a({_al_u2117_o,_al_u2117_o}),
    .b({\PWM5/n24 ,\PWM5/n24 }),
    .c({pnumcnt5[22],pnumcnt5[22]}),
    .clk(clk100m),
    .d({\PWM5/pnumr [22],\PWM5/pnumr [22]}),
    .mi({open_n9585,pwm_start_stop[21]}),
    .q({open_n9592,\PWM5/RemaTxNum[22]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg3_b23  (
    .a({_al_u2115_o,_al_u2115_o}),
    .b({\PWM5/n24 ,\PWM5/n24 }),
    .c({pnumcnt5[23],pnumcnt5[23]}),
    .clk(clk100m),
    .d({\PWM5/pnumr [23],\PWM5/pnumr [23]}),
    .mi({open_n9604,pwm_start_stop[21]}),
    .q({open_n9611,\PWM5/RemaTxNum[23]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg3_b5  (
    .a({_al_u2109_o,_al_u2109_o}),
    .b({\PWM5/n24 ,\PWM5/n24 }),
    .c({pnumcnt5[5],pnumcnt5[5]}),
    .clk(clk100m),
    .d({\PWM5/pnumr [5],\PWM5/pnumr [5]}),
    .mi({open_n9623,pwm_start_stop[21]}),
    .q({open_n9630,\PWM5/RemaTxNum[5]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg3_b6  (
    .a({_al_u2107_o,_al_u2107_o}),
    .b({\PWM5/n24 ,\PWM5/n24 }),
    .c({pnumcnt5[6],pnumcnt5[6]}),
    .clk(clk100m),
    .d({\PWM5/pnumr [6],\PWM5/pnumr [6]}),
    .mi({open_n9642,pwm_start_stop[21]}),
    .q({open_n9649,\PWM5/RemaTxNum[6]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/reg3_b9  (
    .a({_al_u2101_o,_al_u2101_o}),
    .b({\PWM5/n24 ,\PWM5/n24 }),
    .c({pnumcnt5[9],pnumcnt5[9]}),
    .clk(clk100m),
    .d({\PWM5/pnumr [9],\PWM5/pnumr [9]}),
    .mi({open_n9661,pwm_start_stop[21]}),
    .q({open_n9668,\PWM5/RemaTxNum[9]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_LSLICE #(
    //.MACRO("PWM5/sub0/ucin_al_u3398"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM5/sub0/u11_al_u3401  (
    .a({\PWM5/FreCnt [13],\PWM5/FreCnt [11]}),
    .b({\PWM5/FreCnt [14],\PWM5/FreCnt [12]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM5/sub0/c11 ),
    .f({\PWM5/n12 [13],\PWM5/n12 [11]}),
    .fco(\PWM5/sub0/c15 ),
    .fx({\PWM5/n12 [14],\PWM5/n12 [12]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM5/sub0/ucin_al_u3398"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM5/sub0/u15_al_u3402  (
    .a({\PWM5/FreCnt [17],\PWM5/FreCnt [15]}),
    .b({\PWM5/FreCnt [18],\PWM5/FreCnt [16]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM5/sub0/c15 ),
    .f({\PWM5/n12 [17],\PWM5/n12 [15]}),
    .fco(\PWM5/sub0/c19 ),
    .fx({\PWM5/n12 [18],\PWM5/n12 [16]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM5/sub0/ucin_al_u3398"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM5/sub0/u19_al_u3403  (
    .a({\PWM5/FreCnt [21],\PWM5/FreCnt [19]}),
    .b({\PWM5/FreCnt [22],\PWM5/FreCnt [20]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM5/sub0/c19 ),
    .f({\PWM5/n12 [21],\PWM5/n12 [19]}),
    .fco(\PWM5/sub0/c23 ),
    .fx({\PWM5/n12 [22],\PWM5/n12 [20]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM5/sub0/ucin_al_u3398"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM5/sub0/u23_al_u3404  (
    .a({\PWM5/FreCnt [25],\PWM5/FreCnt [23]}),
    .b({\PWM5/FreCnt [26],\PWM5/FreCnt [24]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM5/sub0/c23 ),
    .f({\PWM5/n12 [25],\PWM5/n12 [23]}),
    .fx({\PWM5/n12 [26],\PWM5/n12 [24]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM5/sub0/ucin_al_u3398"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM5/sub0/u3_al_u3399  (
    .a({\PWM5/FreCnt [5],\PWM5/FreCnt [3]}),
    .b({\PWM5/FreCnt [6],\PWM5/FreCnt [4]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM5/sub0/c3 ),
    .f({\PWM5/n12 [5],\PWM5/n12 [3]}),
    .fco(\PWM5/sub0/c7 ),
    .fx({\PWM5/n12 [6],\PWM5/n12 [4]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM5/sub0/ucin_al_u3398"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM5/sub0/u7_al_u3400  (
    .a({\PWM5/FreCnt [9],\PWM5/FreCnt [7]}),
    .b({\PWM5/FreCnt [10],\PWM5/FreCnt [8]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM5/sub0/c7 ),
    .f({\PWM5/n12 [9],\PWM5/n12 [7]}),
    .fco(\PWM5/sub0/c11 ),
    .fx({\PWM5/n12 [10],\PWM5/n12 [8]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM5/sub0/ucin_al_u3398"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'h0005),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM5/sub0/ucin_al_u3398  (
    .a({\PWM5/FreCnt [1],1'b0}),
    .b({\PWM5/FreCnt [2],\PWM5/FreCnt [0]}),
    .c(2'b11),
    .ce(\U_AHB/n14 ),
    .clk(clk100m),
    .d(2'b01),
    .e(2'b01),
    .mi({open_n9779,\U_AHB/h2h_hwdata [2]}),
    .f({\PWM5/n12 [1],open_n9792}),
    .fco(\PWM5/sub0/c3 ),
    .fx({\PWM5/n12 [2],\PWM5/n12 [0]}),
    .q({open_n9793,freq5[2]}));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM5/sub1/u0|PWM5/sub1/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("SUB_CARRY"),
    .INIT_LUT0(16'b0000000000000101),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM5/sub1/u0|PWM5/sub1/ucin  (
    .a({pnumcnt5[0],1'b0}),
    .b({1'b1,open_n9794}),
    .f({\PWM5/n26 [0],open_n9814}),
    .fco(\PWM5/sub1/c1 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM5/sub1/u0|PWM5/sub1/ucin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM5/sub1/u10|PWM5/sub1/u9  (
    .a(pnumcnt5[10:9]),
    .b(2'b00),
    .fci(\PWM5/sub1/c9 ),
    .f(\PWM5/n26 [10:9]),
    .fco(\PWM5/sub1/c11 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM5/sub1/u0|PWM5/sub1/ucin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM5/sub1/u12|PWM5/sub1/u11  (
    .a(pnumcnt5[12:11]),
    .b(2'b00),
    .fci(\PWM5/sub1/c11 ),
    .f(\PWM5/n26 [12:11]),
    .fco(\PWM5/sub1/c13 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM5/sub1/u0|PWM5/sub1/ucin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM5/sub1/u14|PWM5/sub1/u13  (
    .a(pnumcnt5[14:13]),
    .b(2'b00),
    .fci(\PWM5/sub1/c13 ),
    .f(\PWM5/n26 [14:13]),
    .fco(\PWM5/sub1/c15 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM5/sub1/u0|PWM5/sub1/ucin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM5/sub1/u16|PWM5/sub1/u15  (
    .a(pnumcnt5[16:15]),
    .b(2'b00),
    .fci(\PWM5/sub1/c15 ),
    .f(\PWM5/n26 [16:15]),
    .fco(\PWM5/sub1/c17 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM5/sub1/u0|PWM5/sub1/ucin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM5/sub1/u18|PWM5/sub1/u17  (
    .a(pnumcnt5[18:17]),
    .b(2'b00),
    .fci(\PWM5/sub1/c17 ),
    .f(\PWM5/n26 [18:17]),
    .fco(\PWM5/sub1/c19 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM5/sub1/u0|PWM5/sub1/ucin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM5/sub1/u20|PWM5/sub1/u19  (
    .a(pnumcnt5[20:19]),
    .b(2'b00),
    .fci(\PWM5/sub1/c19 ),
    .f(\PWM5/n26 [20:19]),
    .fco(\PWM5/sub1/c21 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM5/sub1/u0|PWM5/sub1/ucin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM5/sub1/u22|PWM5/sub1/u21  (
    .a(pnumcnt5[22:21]),
    .b(2'b00),
    .fci(\PWM5/sub1/c21 ),
    .f(\PWM5/n26 [22:21]),
    .fco(\PWM5/sub1/c23 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM5/sub1/u0|PWM5/sub1/ucin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM5/sub1/u23_al_u3473  (
    .a({open_n9973,pnumcnt5[23]}),
    .b({open_n9974,1'b0}),
    .fci(\PWM5/sub1/c23 ),
    .f({open_n9993,\PWM5/n26 [23]}));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM5/sub1/u0|PWM5/sub1/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM5/sub1/u2|PWM5/sub1/u1  (
    .a(pnumcnt5[2:1]),
    .b(2'b00),
    .fci(\PWM5/sub1/c1 ),
    .f(\PWM5/n26 [2:1]),
    .fco(\PWM5/sub1/c3 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM5/sub1/u0|PWM5/sub1/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM5/sub1/u4|PWM5/sub1/u3  (
    .a(pnumcnt5[4:3]),
    .b(2'b00),
    .fci(\PWM5/sub1/c3 ),
    .f(\PWM5/n26 [4:3]),
    .fco(\PWM5/sub1/c5 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM5/sub1/u0|PWM5/sub1/ucin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM5/sub1/u6|PWM5/sub1/u5  (
    .a(pnumcnt5[6:5]),
    .b(2'b00),
    .fci(\PWM5/sub1/c5 ),
    .f(\PWM5/n26 [6:5]),
    .fco(\PWM5/sub1/c7 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM5/sub1/u0|PWM5/sub1/ucin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM5/sub1/u8|PWM5/sub1/u7  (
    .a(pnumcnt5[8:7]),
    .b(2'b00),
    .fci(\PWM5/sub1/c7 ),
    .f(\PWM5/n26 [8:7]),
    .fco(\PWM5/sub1/c9 ));
  // src/OnePWM.v(26)
  // src/OnePWM.v(26)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*~(~D*B*~A))"),
    //.LUT1("(C*~(~D*B*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000010110000),
    .INIT_LUT1(16'b1111000010110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \PWM6/State_reg|PWM9/State_reg  (
    .a({_al_u3025_o,_al_u3034_o}),
    .b({\PWM6/n0_lutinv ,\PWM9/n0_lutinv }),
    .c({_al_u3026_o,_al_u3035_o}),
    .clk(clk100m),
    .d({pwm_start_stop[22],pwm_start_stop[25]}),
    .sr(rstn),
    .q({pwm_state_read[6],pwm_state_read[9]}));  // src/OnePWM.v(26)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[0]  (
    .i(\PWM6/RemaTxNum[0]_keep ),
    .o(pnumcnt6[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[10]  (
    .i(\PWM6/RemaTxNum[10]_keep ),
    .o(pnumcnt6[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[11]  (
    .i(\PWM6/RemaTxNum[11]_keep ),
    .o(pnumcnt6[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[12]  (
    .i(\PWM6/RemaTxNum[12]_keep ),
    .o(pnumcnt6[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[13]  (
    .i(\PWM6/RemaTxNum[13]_keep ),
    .o(pnumcnt6[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[14]  (
    .i(\PWM6/RemaTxNum[14]_keep ),
    .o(pnumcnt6[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[15]  (
    .i(\PWM6/RemaTxNum[15]_keep ),
    .o(pnumcnt6[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[16]  (
    .i(\PWM6/RemaTxNum[16]_keep ),
    .o(pnumcnt6[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[17]  (
    .i(\PWM6/RemaTxNum[17]_keep ),
    .o(pnumcnt6[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[18]  (
    .i(\PWM6/RemaTxNum[18]_keep ),
    .o(pnumcnt6[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[19]  (
    .i(\PWM6/RemaTxNum[19]_keep ),
    .o(pnumcnt6[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[1]  (
    .i(\PWM6/RemaTxNum[1]_keep ),
    .o(pnumcnt6[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[20]  (
    .i(\PWM6/RemaTxNum[20]_keep ),
    .o(pnumcnt6[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[21]  (
    .i(\PWM6/RemaTxNum[21]_keep ),
    .o(pnumcnt6[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[22]  (
    .i(\PWM6/RemaTxNum[22]_keep ),
    .o(pnumcnt6[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[23]  (
    .i(\PWM6/RemaTxNum[23]_keep ),
    .o(pnumcnt6[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[2]  (
    .i(\PWM6/RemaTxNum[2]_keep ),
    .o(pnumcnt6[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[3]  (
    .i(\PWM6/RemaTxNum[3]_keep ),
    .o(pnumcnt6[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[4]  (
    .i(\PWM6/RemaTxNum[4]_keep ),
    .o(pnumcnt6[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[5]  (
    .i(\PWM6/RemaTxNum[5]_keep ),
    .o(pnumcnt6[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[6]  (
    .i(\PWM6/RemaTxNum[6]_keep ),
    .o(pnumcnt6[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[7]  (
    .i(\PWM6/RemaTxNum[7]_keep ),
    .o(pnumcnt6[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[8]  (
    .i(\PWM6/RemaTxNum[8]_keep ),
    .o(pnumcnt6[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[9]  (
    .i(\PWM6/RemaTxNum[9]_keep ),
    .o(pnumcnt6[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_dir  (
    .i(\PWM6/dir_keep ),
    .o(dir_pad[6]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[0]  (
    .i(\PWM6/pnumr[0]_keep ),
    .o(\PWM6/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[10]  (
    .i(\PWM6/pnumr[10]_keep ),
    .o(\PWM6/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[11]  (
    .i(\PWM6/pnumr[11]_keep ),
    .o(\PWM6/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[12]  (
    .i(\PWM6/pnumr[12]_keep ),
    .o(\PWM6/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[13]  (
    .i(\PWM6/pnumr[13]_keep ),
    .o(\PWM6/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[14]  (
    .i(\PWM6/pnumr[14]_keep ),
    .o(\PWM6/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[15]  (
    .i(\PWM6/pnumr[15]_keep ),
    .o(\PWM6/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[16]  (
    .i(\PWM6/pnumr[16]_keep ),
    .o(\PWM6/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[17]  (
    .i(\PWM6/pnumr[17]_keep ),
    .o(\PWM6/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[18]  (
    .i(\PWM6/pnumr[18]_keep ),
    .o(\PWM6/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[19]  (
    .i(\PWM6/pnumr[19]_keep ),
    .o(\PWM6/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[1]  (
    .i(\PWM6/pnumr[1]_keep ),
    .o(\PWM6/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[20]  (
    .i(\PWM6/pnumr[20]_keep ),
    .o(\PWM6/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[21]  (
    .i(\PWM6/pnumr[21]_keep ),
    .o(\PWM6/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[22]  (
    .i(\PWM6/pnumr[22]_keep ),
    .o(\PWM6/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[23]  (
    .i(\PWM6/pnumr[23]_keep ),
    .o(\PWM6/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[24]  (
    .i(\PWM6/pnumr[24]_keep ),
    .o(\PWM6/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[25]  (
    .i(\PWM6/pnumr[25]_keep ),
    .o(\PWM6/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[26]  (
    .i(\PWM6/pnumr[26]_keep ),
    .o(\PWM6/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[27]  (
    .i(\PWM6/pnumr[27]_keep ),
    .o(\PWM6/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[28]  (
    .i(\PWM6/pnumr[28]_keep ),
    .o(\PWM6/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[29]  (
    .i(\PWM6/pnumr[29]_keep ),
    .o(\PWM6/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[2]  (
    .i(\PWM6/pnumr[2]_keep ),
    .o(\PWM6/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[30]  (
    .i(\PWM6/pnumr[30]_keep ),
    .o(\PWM6/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[31]  (
    .i(\PWM6/pnumr[31]_keep ),
    .o(\PWM6/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[3]  (
    .i(\PWM6/pnumr[3]_keep ),
    .o(\PWM6/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[4]  (
    .i(\PWM6/pnumr[4]_keep ),
    .o(\PWM6/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[5]  (
    .i(\PWM6/pnumr[5]_keep ),
    .o(\PWM6/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[6]  (
    .i(\PWM6/pnumr[6]_keep ),
    .o(\PWM6/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[7]  (
    .i(\PWM6/pnumr[7]_keep ),
    .o(\PWM6/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[8]  (
    .i(\PWM6/pnumr[8]_keep ),
    .o(\PWM6/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[9]  (
    .i(\PWM6/pnumr[9]_keep ),
    .o(\PWM6/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pwm  (
    .i(\PWM6/pwm_keep ),
    .o(pwm_pad[6]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_stopreq  (
    .i(\PWM6/stopreq_keep ),
    .o(\PWM6/stopreq ));  // src/OnePWM.v(14)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM6/reg0_b0|PWM6/reg0_b8  (
    .b({\PWM6/n12 [0],\PWM6/n12 [8]}),
    .c({freq6[0],freq6[8]}),
    .clk(clk100m),
    .d({\PWM6/n0_lutinv ,\PWM6/n0_lutinv }),
    .sr(\PWM6/n11 ),
    .q({\PWM6/FreCnt [0],\PWM6/FreCnt [8]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM6/reg0_b10|PWM6/reg0_b7  (
    .b({\PWM6/n12 [10],\PWM6/n12 [7]}),
    .c({freq6[10],freq6[7]}),
    .clk(clk100m),
    .d({\PWM6/n0_lutinv ,\PWM6/n0_lutinv }),
    .sr(\PWM6/n11 ),
    .q({\PWM6/FreCnt [10],\PWM6/FreCnt [7]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM6/reg0_b11|PWM6/reg0_b5  (
    .b({\PWM6/n12 [11],\PWM6/n12 [5]}),
    .c({freq6[11],freq6[5]}),
    .clk(clk100m),
    .d({\PWM6/n0_lutinv ,\PWM6/n0_lutinv }),
    .sr(\PWM6/n11 ),
    .q({\PWM6/FreCnt [11],\PWM6/FreCnt [5]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM6/reg0_b12|PWM6/reg0_b3  (
    .b({\PWM6/n12 [12],\PWM6/n12 [3]}),
    .c({freq6[12],freq6[3]}),
    .clk(clk100m),
    .d({\PWM6/n0_lutinv ,\PWM6/n0_lutinv }),
    .sr(\PWM6/n11 ),
    .q({\PWM6/FreCnt [12],\PWM6/FreCnt [3]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM6/reg0_b13|PWM6/reg0_b25  (
    .b({\PWM6/n12 [13],\PWM6/n12 [25]}),
    .c({freq6[13],freq6[25]}),
    .clk(clk100m),
    .d({\PWM6/n0_lutinv ,\PWM6/n0_lutinv }),
    .sr(\PWM6/n11 ),
    .q({\PWM6/FreCnt [13],\PWM6/FreCnt [25]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM6/reg0_b14|PWM6/reg0_b22  (
    .b({\PWM6/n12 [14],\PWM6/n12 [22]}),
    .c({freq6[14],freq6[22]}),
    .clk(clk100m),
    .d({\PWM6/n0_lutinv ,\PWM6/n0_lutinv }),
    .sr(\PWM6/n11 ),
    .q({\PWM6/FreCnt [14],\PWM6/FreCnt [22]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM6/reg0_b15|PWM6/reg0_b21  (
    .b({\PWM6/n12 [15],\PWM6/n12 [21]}),
    .c({freq6[15],freq6[21]}),
    .clk(clk100m),
    .d({\PWM6/n0_lutinv ,\PWM6/n0_lutinv }),
    .sr(\PWM6/n11 ),
    .q({\PWM6/FreCnt [15],\PWM6/FreCnt [21]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM6/reg0_b16|PWM6/reg0_b19  (
    .b({\PWM6/n12 [16],\PWM6/n12 [19]}),
    .c({freq6[16],freq6[19]}),
    .clk(clk100m),
    .d({\PWM6/n0_lutinv ,\PWM6/n0_lutinv }),
    .sr(\PWM6/n11 ),
    .q({\PWM6/FreCnt [16],\PWM6/FreCnt [19]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM6/reg0_b18|PWM6/reg0_b17  (
    .b(\PWM6/n12 [18:17]),
    .c(freq6[18:17]),
    .clk(clk100m),
    .d({\PWM6/n0_lutinv ,\PWM6/n0_lutinv }),
    .sr(\PWM6/n11 ),
    .q(\PWM6/FreCnt [18:17]));  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM6/reg0_b2  (
    .b({open_n10307,\PWM6/n12 [2]}),
    .c({open_n10308,freq6[2]}),
    .clk(clk100m),
    .d({open_n10310,\PWM6/n0_lutinv }),
    .sr(\PWM6/n11 ),
    .q({open_n10328,\PWM6/FreCnt [2]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM6/reg0_b20|PWM6/reg0_b1  (
    .b({\PWM6/n12 [20],\PWM6/n12 [1]}),
    .c({freq6[20],freq6[1]}),
    .clk(clk100m),
    .d({\PWM6/n0_lutinv ,\PWM6/n0_lutinv }),
    .sr(\PWM6/n11 ),
    .q({\PWM6/FreCnt [20],\PWM6/FreCnt [1]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM6/reg0_b23|PWM6/reg0_b9  (
    .b({\PWM6/n12 [23],\PWM6/n12 [9]}),
    .c({freq6[23],freq6[9]}),
    .clk(clk100m),
    .d({\PWM6/n0_lutinv ,\PWM6/n0_lutinv }),
    .sr(\PWM6/n11 ),
    .q({\PWM6/FreCnt [23],\PWM6/FreCnt [9]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM6/reg0_b24|PWM6/reg0_b6  (
    .b({\PWM6/n12 [24],\PWM6/n12 [6]}),
    .c({freq6[24],freq6[6]}),
    .clk(clk100m),
    .d({\PWM6/n0_lutinv ,\PWM6/n0_lutinv }),
    .sr(\PWM6/n11 ),
    .q({\PWM6/FreCnt [24],\PWM6/FreCnt [6]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM6/reg0_b26|PWM6/reg0_b4  (
    .b({\PWM6/n12 [26],\PWM6/n12 [4]}),
    .c({freq6[26],freq6[4]}),
    .clk(clk100m),
    .d({\PWM6/n0_lutinv ,\PWM6/n0_lutinv }),
    .sr(\PWM6/n11 ),
    .q({\PWM6/FreCnt [26],\PWM6/FreCnt [4]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*~C)*~(D*~B))"),
    //.LUTF1("(A*~(~0*C)*~(D*~B))"),
    //.LUTG0("(A*~(1*~C)*~(D*~B))"),
    //.LUTG1("(A*~(~1*C)*~(D*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000100010101010),
    .INIT_LUTF1(16'b0000100000001010),
    .INIT_LUTG0(16'b1000000010100000),
    .INIT_LUTG1(16'b1000100010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg1_b11|PWM6/reg1_b26  (
    .a({_al_u2235_o,_al_u2231_o}),
    .b({\PWM6/FreCnt [10],\PWM6/FreCnt [17]}),
    .c({\PWM6/FreCnt [25],\PWM6/FreCnt [25]}),
    .ce(\PWM6/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM6/FreCntr [11],\PWM6/FreCntr [18]}),
    .e({\PWM6/FreCntr [26],\PWM6/FreCntr [26]}),
    .mi({freq6[11],freq6[26]}),
    .f({_al_u2236_o,_al_u2232_o}),
    .q({\PWM6/FreCntr [11],\PWM6/FreCntr [26]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(D*~B)*~(C*~A))"),
    //.LUT1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000110010101111),
    .INIT_LUT1(16'b1000010000100001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg1_b14|PWM6/reg1_b8  (
    .a({\PWM6/FreCnt [13],\PWM6/FreCnt [7]}),
    .b({\PWM6/FreCnt [14],\PWM6/FreCnt [8]}),
    .c({\PWM6/FreCntr [14],\PWM6/FreCntr [8]}),
    .ce(\PWM6/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM6/FreCntr [15],\PWM6/FreCntr [9]}),
    .mi({freq6[14],freq6[8]}),
    .f({_al_u2248_o,_al_u2243_o}),
    .q({\PWM6/FreCntr [14],\PWM6/FreCntr [8]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~A*~(0*~C)*~(D@B))"),
    //.LUTF1("(A*~(0@C)*~(D@B))"),
    //.LUTG0("(~A*~(1*~C)*~(D@B))"),
    //.LUTG1("(A*~(1@C)*~(D@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100010000010001),
    .INIT_LUTF1(16'b0000100000000010),
    .INIT_LUTG0(16'b0100000000010000),
    .INIT_LUTG1(16'b1000000000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg1_b15|PWM6/reg1_b12  (
    .a({_al_u1470_o,_al_u2245_o}),
    .b(\PWM6/FreCnt [12:11]),
    .c({\PWM6/FreCnt [15],\PWM6/FreCnt [22]}),
    .ce(\PWM6/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM6/FreCntr [12],\PWM6/FreCntr [12]}),
    .e({\PWM6/FreCntr [15],\PWM6/FreCntr [23]}),
    .mi({freq6[15],freq6[12]}),
    .f({_al_u1471_o,_al_u2246_o}),
    .q({\PWM6/FreCntr [15],\PWM6/FreCntr [12]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*B*A*~(0@D))"),
    //.LUTF1("(~(D*~B)*~(~C*A))"),
    //.LUTG0("(C*B*A*~(1@D))"),
    //.LUTG1("(~(D*~B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b1100010011110101),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b1100010011110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg1_b16|PWM6/reg1_b13  (
    .a({\PWM6/FreCnt [15],_al_u2249_o}),
    .b({\PWM6/FreCnt [21],_al_u2251_o}),
    .c({\PWM6/FreCntr [16],_al_u2252_o}),
    .ce(\PWM6/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM6/FreCntr [22],\PWM6/FreCnt [12]}),
    .e({open_n10467,\PWM6/FreCntr [13]}),
    .mi({freq6[16],freq6[13]}),
    .f({_al_u2252_o,_al_u2253_o}),
    .q({\PWM6/FreCntr [16],\PWM6/FreCntr [13]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg1_b1|PWM6/reg1_b19  (
    .a({\PWM6/FreCnt [0],_al_u1472_o}),
    .b({\PWM6/FreCnt [18],\PWM6/FreCnt [13]}),
    .c({\PWM6/FreCntr [1],\PWM6/FreCnt [19]}),
    .ce(\PWM6/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM6/FreCntr [19],\PWM6/FreCntr [13]}),
    .e({open_n10484,\PWM6/FreCntr [19]}),
    .mi({freq6[1],freq6[19]}),
    .f({_al_u2241_o,_al_u1473_o}),
    .q({\PWM6/FreCntr [1],\PWM6/FreCntr [19]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(D*~B)*~(~C*A))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~(D*~B)*~(~C*A))"),
    //.LUTG1("(~C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100010011110101),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1100010011110101),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg1_b20|PWM6/reg1_b22  (
    .a({open_n10501,\PWM6/FreCnt [21]}),
    .b({open_n10502,\PWM6/FreCnt [5]}),
    .c({\PWM6/FreCntr [20],\PWM6/FreCntr [22]}),
    .ce(\PWM6/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM6/FreCnt [19],\PWM6/FreCntr [6]}),
    .mi({freq6[20],freq6[22]}),
    .f({_al_u2245_o,_al_u2233_o}),
    .q({\PWM6/FreCntr [20],\PWM6/FreCntr [22]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D@C)*~(0@B))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(A*~(D@C)*~(1@B))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010000000000010),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000000000001000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg1_b21|PWM6/reg1_b10  (
    .a({\PWM6/FreCnt [1],_al_u2248_o}),
    .b(\PWM6/FreCnt [21:20]),
    .c({\PWM6/FreCntr [1],\PWM6/FreCnt [9]}),
    .ce(\PWM6/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM6/FreCntr [21],\PWM6/FreCntr [10]}),
    .e({open_n10521,\PWM6/FreCntr [21]}),
    .mi({freq6[21],freq6[10]}),
    .f({_al_u1470_o,_al_u2249_o}),
    .q({\PWM6/FreCntr [21],\PWM6/FreCntr [10]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(A*~(0@C)*~(D@B))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(A*~(1@C)*~(D@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b0000100000000010),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000000000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg1_b25|PWM6/reg1_b24  (
    .a({_al_u2239_o,_al_u1466_o}),
    .b({\PWM6/FreCnt [24],\PWM6/FreCnt [24]}),
    .c({\PWM6/FreCnt [6],\PWM6/FreCnt [7]}),
    .ce(\PWM6/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d(\PWM6/FreCntr [25:24]),
    .e({\PWM6/FreCntr [7],\PWM6/FreCntr [7]}),
    .mi(freq6[25:24]),
    .f({_al_u2240_o,_al_u1467_o}),
    .q(\PWM6/FreCntr [25:24]));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~C*~(~D*B)*~(0@A))"),
    //.LUTF1("(A*~(0@C)*~(D@B))"),
    //.LUTG0("(~C*~(~D*B)*~(1@A))"),
    //.LUTG1("(A*~(1@C)*~(D@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010100000001),
    .INIT_LUTF1(16'b0000100000000010),
    .INIT_LUTG0(16'b0000101000000010),
    .INIT_LUTG1(16'b1000000000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg1_b3|PWM6/reg1_b23  (
    .a({_al_u1476_o,\PWM6/FreCnt [2]}),
    .b({\PWM6/FreCnt [2],\PWM6/FreCnt [22]}),
    .c({\PWM6/FreCnt [3],\PWM6/FreCnt [26]}),
    .ce(\PWM6/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM6/FreCntr [2],\PWM6/FreCntr [23]}),
    .e({\PWM6/FreCntr [3],\PWM6/FreCntr [3]}),
    .mi({freq6[3],freq6[23]}),
    .f({_al_u1477_o,_al_u2239_o}),
    .q({\PWM6/FreCntr [3],\PWM6/FreCntr [23]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(~0*C)*~(~D*B))"),
    //.LUTF1("(~(~D*B)*~(C*~A))"),
    //.LUTG0("(A*~(~1*C)*~(~D*B))"),
    //.LUTG1("(~(~D*B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101000000010),
    .INIT_LUTF1(16'b1010111100100011),
    .INIT_LUTG0(16'b1010101000100010),
    .INIT_LUTG1(16'b1010111100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg1_b4|PWM6/reg1_b18  (
    .a({\PWM6/FreCnt [3],_al_u2243_o}),
    .b({\PWM6/FreCnt [7],\PWM6/FreCnt [17]}),
    .c({\PWM6/FreCntr [4],\PWM6/FreCnt [3]}),
    .ce(\PWM6/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM6/FreCntr [8],\PWM6/FreCntr [18]}),
    .e({open_n10570,\PWM6/FreCntr [4]}),
    .mi({freq6[4],freq6[18]}),
    .f({_al_u2235_o,_al_u2244_o}),
    .q({\PWM6/FreCntr [4],\PWM6/FreCntr [18]}));  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(D*~(C@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100001100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg1_b5  (
    .b({open_n10589,\PWM6/FreCnt [4]}),
    .c({open_n10590,\PWM6/FreCntr [5]}),
    .ce(\PWM6/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({open_n10591,_al_u2241_o}),
    .mi({open_n10602,freq6[5]}),
    .f({open_n10604,_al_u2242_o}),
    .q({open_n10608,\PWM6/FreCntr [5]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~A*~(0@C)*~(~D*B))"),
    //.LUTF1("(~(~D*B)*~(C*~A))"),
    //.LUTG0("(~A*~(1@C)*~(~D*B))"),
    //.LUTG1("(~(~D*B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010100000001),
    .INIT_LUTF1(16'b1010111100100011),
    .INIT_LUTG0(16'b0101000000010000),
    .INIT_LUTG1(16'b1010111100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg1_b6|PWM6/reg1_b2  (
    .a({\PWM6/FreCnt [1],_al_u2250_o}),
    .b({\PWM6/FreCnt [5],\PWM6/FreCnt [1]}),
    .c({\PWM6/FreCntr [2],\PWM6/FreCnt [23]}),
    .ce(\PWM6/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM6/FreCntr [6],\PWM6/FreCntr [2]}),
    .e({open_n10609,\PWM6/FreCntr [24]}),
    .mi({freq6[6],freq6[2]}),
    .f({_al_u2237_o,_al_u2251_o}),
    .q({\PWM6/FreCntr [6],\PWM6/FreCntr [2]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg1_b7|PWM6/reg1_b0  (
    .b({_al_u960_o,open_n10628}),
    .c({_al_u962_o,\PWM6/n11 }),
    .ce(\PWM6/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({_al_u958_o,\PWM6/n0_lutinv }),
    .mi({freq6[7],freq6[0]}),
    .f({\PWM6/n0_lutinv ,\PWM6/mux3_b0_sel_is_3_o }),
    .q({\PWM6/FreCntr [7],\PWM6/FreCntr [0]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*B*A*~(0@D))"),
    //.LUTF1("(B*A*~(~D*C))"),
    //.LUTG0("(C*B*A*~(1@D))"),
    //.LUTG1("(B*A*~(~D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b1000100000001000),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b1000100000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg1_b9|PWM6/reg1_b17  (
    .a({_al_u2232_o,_al_u2234_o}),
    .b({_al_u2233_o,_al_u2236_o}),
    .c({\PWM6/FreCnt [8],_al_u2237_o}),
    .ce(\PWM6/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM6/FreCntr [9],\PWM6/FreCnt [16]}),
    .e({open_n10647,\PWM6/FreCntr [17]}),
    .mi({freq6[9],freq6[17]}),
    .f({_al_u2234_o,_al_u2238_o}),
    .q({\PWM6/FreCntr [9],\PWM6/FreCntr [17]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011100010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg2_b0|PWM6/reg2_b7  (
    .a({\PWM6/pnumr [0],\PWM6/pnumr [7]}),
    .b({pnum6[0],pnum6[32]}),
    .c({pnum6[32],pnum6[7]}),
    .clk(clk100m),
    .d({pwm_start_stop[22],pwm_start_stop[22]}),
    .q({\PWM6/pnumr[0]_keep ,\PWM6/pnumr[7]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg2_b10|PWM6/reg3_b10  (
    .a({\PWM6/pnumr [10],_al_u2225_o}),
    .b({pnum6[10],\PWM6/n24 }),
    .c({pnum6[32],pnumcnt6[10]}),
    .clk(clk100m),
    .d({pwm_start_stop[22],\PWM6/pnumr [10]}),
    .e({open_n10684,pwm_start_stop[22]}),
    .q({\PWM6/pnumr[10]_keep ,\PWM6/RemaTxNum[10]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg2_b11|PWM6/reg3_b11  (
    .a({\PWM6/pnumr [11],_al_u2223_o}),
    .b({pnum6[11],\PWM6/n24 }),
    .c({pnum6[32],pnumcnt6[11]}),
    .clk(clk100m),
    .d({pwm_start_stop[22],\PWM6/pnumr [11]}),
    .e({open_n10706,pwm_start_stop[22]}),
    .q({\PWM6/pnumr[11]_keep ,\PWM6/RemaTxNum[11]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011100010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011100010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg2_b12|PWM6/reg2_b6  (
    .a({\PWM6/pnumr [12],\PWM6/pnumr [6]}),
    .b({pnum6[12],pnum6[32]}),
    .c({pnum6[32],pnum6[6]}),
    .clk(clk100m),
    .d({pwm_start_stop[22],pwm_start_stop[22]}),
    .q({\PWM6/pnumr[12]_keep ,\PWM6/pnumr[6]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg2_b13|PWM6/reg2_b3  (
    .a({\PWM6/pnumr [13],\PWM6/pnumr [3]}),
    .b({pnum6[13],pnum6[3]}),
    .c({pnum6[32],pnum6[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[22],pwm_start_stop[22]}),
    .q({\PWM6/pnumr[13]_keep ,\PWM6/pnumr[3]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg2_b14|PWM6/reg3_b14  (
    .a({\PWM6/pnumr [14],_al_u2217_o}),
    .b({pnum6[14],\PWM6/n24 }),
    .c({pnum6[32],pnumcnt6[14]}),
    .clk(clk100m),
    .d({pwm_start_stop[22],\PWM6/pnumr [14]}),
    .e({open_n10774,pwm_start_stop[22]}),
    .q({\PWM6/pnumr[14]_keep ,\PWM6/RemaTxNum[14]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg2_b15|PWM6/reg3_b15  (
    .a({\PWM6/pnumr [15],_al_u2215_o}),
    .b({pnum6[15],\PWM6/n24 }),
    .c({pnum6[32],pnumcnt6[15]}),
    .clk(clk100m),
    .d({pwm_start_stop[22],\PWM6/pnumr [15]}),
    .e({open_n10796,pwm_start_stop[22]}),
    .q({\PWM6/pnumr[15]_keep ,\PWM6/RemaTxNum[15]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg2_b16|PWM6/reg2_b23  (
    .a({\PWM6/pnumr [16],\PWM6/pnumr [23]}),
    .b({pnum6[16],pnum6[23]}),
    .c({pnum6[32],pnum6[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[22],pwm_start_stop[22]}),
    .q({\PWM6/pnumr[16]_keep ,\PWM6/pnumr[23]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg2_b17|PWM6/reg2_b20  (
    .a({\PWM6/pnumr [17],\PWM6/pnumr [20]}),
    .b({pnum6[17],pnum6[20]}),
    .c({pnum6[32],pnum6[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[22],pwm_start_stop[22]}),
    .q({\PWM6/pnumr[17]_keep ,\PWM6/pnumr[20]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg2_b18|PWM6/reg3_b18  (
    .a({\PWM6/pnumr [18],_al_u2209_o}),
    .b({pnum6[18],\PWM6/n24 }),
    .c({pnum6[32],pnumcnt6[18]}),
    .clk(clk100m),
    .d({pwm_start_stop[22],\PWM6/pnumr [18]}),
    .e({open_n10856,pwm_start_stop[22]}),
    .q({\PWM6/pnumr[18]_keep ,\PWM6/RemaTxNum[18]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg2_b19|PWM6/reg3_b19  (
    .a({\PWM6/pnumr [19],_al_u2207_o}),
    .b({pnum6[19],\PWM6/n24 }),
    .c({pnum6[32],pnumcnt6[19]}),
    .clk(clk100m),
    .d({pwm_start_stop[22],\PWM6/pnumr [19]}),
    .e({open_n10878,pwm_start_stop[22]}),
    .q({\PWM6/pnumr[19]_keep ,\PWM6/RemaTxNum[19]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg2_b1|PWM6/reg2_b2  (
    .a({\PWM6/pnumr [1],\PWM6/pnumr [2]}),
    .b({pnum6[1],pnum6[2]}),
    .c({pnum6[32],pnum6[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[22],pwm_start_stop[22]}),
    .q({\PWM6/pnumr[1]_keep ,\PWM6/pnumr[2]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg2_b21|PWM6/reg3_b21  (
    .a({\PWM6/pnumr [21],_al_u2201_o}),
    .b({pnum6[21],\PWM6/n24 }),
    .c({pnum6[32],pnumcnt6[21]}),
    .clk(clk100m),
    .d({pwm_start_stop[22],\PWM6/pnumr [21]}),
    .e({open_n10923,pwm_start_stop[22]}),
    .q({\PWM6/pnumr[21]_keep ,\PWM6/RemaTxNum[21]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg2_b22|PWM6/reg3_b22  (
    .a({\PWM6/pnumr [22],_al_u2199_o}),
    .b({pnum6[22],\PWM6/n24 }),
    .c({pnum6[32],pnumcnt6[22]}),
    .clk(clk100m),
    .d({pwm_start_stop[22],\PWM6/pnumr [22]}),
    .e({open_n10945,pwm_start_stop[22]}),
    .q({\PWM6/pnumr[22]_keep ,\PWM6/RemaTxNum[22]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg2_b24|PWM6/reg2_b30  (
    .a({\PWM6/pnumr [24],\PWM6/pnumr [30]}),
    .b({pnum6[24],pnum6[30]}),
    .c({pnum6[32],pnum6[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[22],pwm_start_stop[22]}),
    .q({\PWM6/pnumr[24]_keep ,\PWM6/pnumr[30]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg2_b25|PWM6/reg2_b29  (
    .a({\PWM6/pnumr [25],\PWM6/pnumr [29]}),
    .b({pnum6[25],pnum6[29]}),
    .c({pnum6[32],pnum6[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[22],pwm_start_stop[22]}),
    .q({\PWM6/pnumr[25]_keep ,\PWM6/pnumr[29]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg2_b26|PWM6/reg2_b28  (
    .a({\PWM6/pnumr [26],\PWM6/pnumr [28]}),
    .b({pnum6[26],pnum6[28]}),
    .c({pnum6[32],pnum6[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[22],pwm_start_stop[22]}),
    .q({\PWM6/pnumr[26]_keep ,\PWM6/pnumr[28]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~((~0*~(B*A)))+D*C*~((~0*~(B*A)))+~(D)*C*(~0*~(B*A))+D*C*(~0*~(B*A)))"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(D*~(C)*~((~1*~(B*A)))+D*C*~((~1*~(B*A)))+~(D)*C*(~1*~(B*A))+D*C*(~1*~(B*A)))"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111100001110000),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg2_b31|PWM6/dir_reg  (
    .a({\PWM6/pnumr [31],\PWM6/n24 }),
    .b({pnum6[31],\PWM6/n25_neg_lutinv }),
    .c({pnum6[32],dir_pad[6]}),
    .clk(clk100m),
    .d({pwm_start_stop[22],\PWM6/pnumr [31]}),
    .e({open_n11028,pwm_start_stop[22]}),
    .q({\PWM6/pnumr[31]_keep ,\PWM6/dir_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg2_b4|PWM6/reg3_b4  (
    .a({\PWM6/pnumr [4],_al_u2193_o}),
    .b({pnum6[32],\PWM6/n24 }),
    .c({pnum6[4],pnumcnt6[4]}),
    .clk(clk100m),
    .d({pwm_start_stop[22],\PWM6/pnumr [4]}),
    .e({open_n11050,pwm_start_stop[22]}),
    .q({\PWM6/pnumr[4]_keep ,\PWM6/RemaTxNum[4]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg2_b5|PWM6/reg3_b5  (
    .a({\PWM6/pnumr [5],_al_u2191_o}),
    .b({pnum6[32],\PWM6/n24 }),
    .c({pnum6[5],pnumcnt6[5]}),
    .clk(clk100m),
    .d({pwm_start_stop[22],\PWM6/pnumr [5]}),
    .e({open_n11072,pwm_start_stop[22]}),
    .q({\PWM6/pnumr[5]_keep ,\PWM6/RemaTxNum[5]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg2_b8|PWM6/reg3_b8  (
    .a({\PWM6/pnumr [8],_al_u2185_o}),
    .b({pnum6[32],\PWM6/n24 }),
    .c({pnum6[8],pnumcnt6[8]}),
    .clk(clk100m),
    .d({pwm_start_stop[22],\PWM6/pnumr [8]}),
    .e({open_n11094,pwm_start_stop[22]}),
    .q({\PWM6/pnumr[8]_keep ,\PWM6/RemaTxNum[8]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg2_b9|PWM6/reg3_b9  (
    .a({\PWM6/pnumr [9],_al_u2183_o}),
    .b({pnum6[32],\PWM6/n24 }),
    .c({pnum6[9],pnumcnt6[9]}),
    .clk(clk100m),
    .d({pwm_start_stop[22],\PWM6/pnumr [9]}),
    .e({open_n11116,pwm_start_stop[22]}),
    .q({\PWM6/pnumr[9]_keep ,\PWM6/RemaTxNum[9]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg3_b0  (
    .a({_al_u2229_o,_al_u2229_o}),
    .b({\PWM6/n24 ,\PWM6/n24 }),
    .c({pnumcnt6[0],pnumcnt6[0]}),
    .clk(clk100m),
    .d({\PWM6/pnumr [0],\PWM6/pnumr [0]}),
    .mi({open_n11148,pwm_start_stop[22]}),
    .q({open_n11155,\PWM6/RemaTxNum[0]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg3_b1  (
    .a({_al_u2227_o,_al_u2227_o}),
    .b({\PWM6/n24 ,\PWM6/n24 }),
    .c({pnumcnt6[1],pnumcnt6[1]}),
    .clk(clk100m),
    .d({\PWM6/pnumr [1],\PWM6/pnumr [1]}),
    .mi({open_n11167,pwm_start_stop[22]}),
    .q({open_n11174,\PWM6/RemaTxNum[1]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg3_b12  (
    .a({_al_u2221_o,_al_u2221_o}),
    .b({\PWM6/n24 ,\PWM6/n24 }),
    .c({pnumcnt6[12],pnumcnt6[12]}),
    .clk(clk100m),
    .d({\PWM6/pnumr [12],\PWM6/pnumr [12]}),
    .mi({open_n11186,pwm_start_stop[22]}),
    .q({open_n11193,\PWM6/RemaTxNum[12]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg3_b13  (
    .a({_al_u2219_o,_al_u2219_o}),
    .b({\PWM6/n24 ,\PWM6/n24 }),
    .c({pnumcnt6[13],pnumcnt6[13]}),
    .clk(clk100m),
    .d({\PWM6/pnumr [13],\PWM6/pnumr [13]}),
    .mi({open_n11205,pwm_start_stop[22]}),
    .q({open_n11212,\PWM6/RemaTxNum[13]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg3_b16  (
    .a({_al_u2213_o,_al_u2213_o}),
    .b({\PWM6/n24 ,\PWM6/n24 }),
    .c({pnumcnt6[16],pnumcnt6[16]}),
    .clk(clk100m),
    .d({\PWM6/pnumr [16],\PWM6/pnumr [16]}),
    .mi({open_n11224,pwm_start_stop[22]}),
    .q({open_n11231,\PWM6/RemaTxNum[16]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg3_b17  (
    .a({_al_u2211_o,_al_u2211_o}),
    .b({\PWM6/n24 ,\PWM6/n24 }),
    .c({pnumcnt6[17],pnumcnt6[17]}),
    .clk(clk100m),
    .d({\PWM6/pnumr [17],\PWM6/pnumr [17]}),
    .mi({open_n11243,pwm_start_stop[22]}),
    .q({open_n11250,\PWM6/RemaTxNum[17]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg3_b2  (
    .a({_al_u2205_o,_al_u2205_o}),
    .b({\PWM6/n24 ,\PWM6/n24 }),
    .c({pnumcnt6[2],pnumcnt6[2]}),
    .clk(clk100m),
    .d({\PWM6/pnumr [2],\PWM6/pnumr [2]}),
    .mi({open_n11262,pwm_start_stop[22]}),
    .q({open_n11269,\PWM6/RemaTxNum[2]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg3_b20  (
    .a({_al_u2203_o,_al_u2203_o}),
    .b({\PWM6/n24 ,\PWM6/n24 }),
    .c({pnumcnt6[20],pnumcnt6[20]}),
    .clk(clk100m),
    .d({\PWM6/pnumr [20],\PWM6/pnumr [20]}),
    .mi({open_n11281,pwm_start_stop[22]}),
    .q({open_n11288,\PWM6/RemaTxNum[20]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg3_b23  (
    .a({_al_u2197_o,_al_u2197_o}),
    .b({\PWM6/n24 ,\PWM6/n24 }),
    .c({pnumcnt6[23],pnumcnt6[23]}),
    .clk(clk100m),
    .d({\PWM6/pnumr [23],\PWM6/pnumr [23]}),
    .mi({open_n11300,pwm_start_stop[22]}),
    .q({open_n11307,\PWM6/RemaTxNum[23]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg3_b3  (
    .a({_al_u2195_o,_al_u2195_o}),
    .b({\PWM6/n24 ,\PWM6/n24 }),
    .c({pnumcnt6[3],pnumcnt6[3]}),
    .clk(clk100m),
    .d({\PWM6/pnumr [3],\PWM6/pnumr [3]}),
    .mi({open_n11319,pwm_start_stop[22]}),
    .q({open_n11326,\PWM6/RemaTxNum[3]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg3_b6  (
    .a({_al_u2189_o,_al_u2189_o}),
    .b({\PWM6/n24 ,\PWM6/n24 }),
    .c({pnumcnt6[6],pnumcnt6[6]}),
    .clk(clk100m),
    .d({\PWM6/pnumr [6],\PWM6/pnumr [6]}),
    .mi({open_n11338,pwm_start_stop[22]}),
    .q({open_n11345,\PWM6/RemaTxNum[6]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/reg3_b7  (
    .a({_al_u2187_o,_al_u2187_o}),
    .b({\PWM6/n24 ,\PWM6/n24 }),
    .c({pnumcnt6[7],pnumcnt6[7]}),
    .clk(clk100m),
    .d({\PWM6/pnumr [7],\PWM6/pnumr [7]}),
    .mi({open_n11357,pwm_start_stop[22]}),
    .q({open_n11364,\PWM6/RemaTxNum[7]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_LSLICE #(
    //.MACRO("PWM6/sub0/ucin_al_u3405"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM6/sub0/u11_al_u3408  (
    .a({\PWM6/FreCnt [13],\PWM6/FreCnt [11]}),
    .b({\PWM6/FreCnt [14],\PWM6/FreCnt [12]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM6/sub0/c11 ),
    .f({\PWM6/n12 [13],\PWM6/n12 [11]}),
    .fco(\PWM6/sub0/c15 ),
    .fx({\PWM6/n12 [14],\PWM6/n12 [12]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM6/sub0/ucin_al_u3405"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM6/sub0/u15_al_u3409  (
    .a({\PWM6/FreCnt [17],\PWM6/FreCnt [15]}),
    .b({\PWM6/FreCnt [18],\PWM6/FreCnt [16]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM6/sub0/c15 ),
    .f({\PWM6/n12 [17],\PWM6/n12 [15]}),
    .fco(\PWM6/sub0/c19 ),
    .fx({\PWM6/n12 [18],\PWM6/n12 [16]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM6/sub0/ucin_al_u3405"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM6/sub0/u19_al_u3410  (
    .a({\PWM6/FreCnt [21],\PWM6/FreCnt [19]}),
    .b({\PWM6/FreCnt [22],\PWM6/FreCnt [20]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM6/sub0/c19 ),
    .f({\PWM6/n12 [21],\PWM6/n12 [19]}),
    .fco(\PWM6/sub0/c23 ),
    .fx({\PWM6/n12 [22],\PWM6/n12 [20]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM6/sub0/ucin_al_u3405"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM6/sub0/u23_al_u3411  (
    .a({\PWM6/FreCnt [25],\PWM6/FreCnt [23]}),
    .b({\PWM6/FreCnt [26],\PWM6/FreCnt [24]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM6/sub0/c23 ),
    .f({\PWM6/n12 [25],\PWM6/n12 [23]}),
    .fx({\PWM6/n12 [26],\PWM6/n12 [24]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM6/sub0/ucin_al_u3405"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM6/sub0/u3_al_u3406  (
    .a({\PWM6/FreCnt [5],\PWM6/FreCnt [3]}),
    .b({\PWM6/FreCnt [6],\PWM6/FreCnt [4]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM6/sub0/c3 ),
    .f({\PWM6/n12 [5],\PWM6/n12 [3]}),
    .fco(\PWM6/sub0/c7 ),
    .fx({\PWM6/n12 [6],\PWM6/n12 [4]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM6/sub0/ucin_al_u3405"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM6/sub0/u7_al_u3407  (
    .a({\PWM6/FreCnt [9],\PWM6/FreCnt [7]}),
    .b({\PWM6/FreCnt [10],\PWM6/FreCnt [8]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM6/sub0/c7 ),
    .f({\PWM6/n12 [9],\PWM6/n12 [7]}),
    .fco(\PWM6/sub0/c11 ),
    .fx({\PWM6/n12 [10],\PWM6/n12 [8]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM6/sub0/ucin_al_u3405"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'h0005),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM6/sub0/ucin_al_u3405  (
    .a({\PWM6/FreCnt [1],1'b0}),
    .b({\PWM6/FreCnt [2],\PWM6/FreCnt [0]}),
    .c(2'b11),
    .ce(\U_AHB/n16 ),
    .clk(clk100m),
    .d(2'b01),
    .e(2'b01),
    .mi(\U_AHB/h2h_hwdata [2:1]),
    .f({\PWM6/n12 [1],open_n11487}),
    .fco(\PWM6/sub0/c3 ),
    .fx({\PWM6/n12 [2],\PWM6/n12 [0]}),
    .q(freq6[2:1]));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM6/sub1/u0|PWM6/sub1/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("SUB_CARRY"),
    .INIT_LUT0(16'b0000000000000101),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM6/sub1/u0|PWM6/sub1/ucin  (
    .a({pnumcnt6[0],1'b0}),
    .b({1'b1,open_n11488}),
    .f({\PWM6/n26 [0],open_n11508}),
    .fco(\PWM6/sub1/c1 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM6/sub1/u0|PWM6/sub1/ucin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM6/sub1/u10|PWM6/sub1/u9  (
    .a(pnumcnt6[10:9]),
    .b(2'b00),
    .fci(\PWM6/sub1/c9 ),
    .f(\PWM6/n26 [10:9]),
    .fco(\PWM6/sub1/c11 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM6/sub1/u0|PWM6/sub1/ucin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM6/sub1/u12|PWM6/sub1/u11  (
    .a(pnumcnt6[12:11]),
    .b(2'b00),
    .fci(\PWM6/sub1/c11 ),
    .f(\PWM6/n26 [12:11]),
    .fco(\PWM6/sub1/c13 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM6/sub1/u0|PWM6/sub1/ucin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM6/sub1/u14|PWM6/sub1/u13  (
    .a(pnumcnt6[14:13]),
    .b(2'b00),
    .fci(\PWM6/sub1/c13 ),
    .f(\PWM6/n26 [14:13]),
    .fco(\PWM6/sub1/c15 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM6/sub1/u0|PWM6/sub1/ucin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM6/sub1/u16|PWM6/sub1/u15  (
    .a(pnumcnt6[16:15]),
    .b(2'b00),
    .fci(\PWM6/sub1/c15 ),
    .f(\PWM6/n26 [16:15]),
    .fco(\PWM6/sub1/c17 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM6/sub1/u0|PWM6/sub1/ucin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM6/sub1/u18|PWM6/sub1/u17  (
    .a(pnumcnt6[18:17]),
    .b(2'b00),
    .fci(\PWM6/sub1/c17 ),
    .f(\PWM6/n26 [18:17]),
    .fco(\PWM6/sub1/c19 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM6/sub1/u0|PWM6/sub1/ucin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM6/sub1/u20|PWM6/sub1/u19  (
    .a(pnumcnt6[20:19]),
    .b(2'b00),
    .fci(\PWM6/sub1/c19 ),
    .f(\PWM6/n26 [20:19]),
    .fco(\PWM6/sub1/c21 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM6/sub1/u0|PWM6/sub1/ucin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM6/sub1/u22|PWM6/sub1/u21  (
    .a(pnumcnt6[22:21]),
    .b(2'b00),
    .fci(\PWM6/sub1/c21 ),
    .f(\PWM6/n26 [22:21]),
    .fco(\PWM6/sub1/c23 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM6/sub1/u0|PWM6/sub1/ucin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM6/sub1/u23_al_u3474  (
    .a({open_n11667,pnumcnt6[23]}),
    .b({open_n11668,1'b0}),
    .fci(\PWM6/sub1/c23 ),
    .f({open_n11687,\PWM6/n26 [23]}));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM6/sub1/u0|PWM6/sub1/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM6/sub1/u2|PWM6/sub1/u1  (
    .a(pnumcnt6[2:1]),
    .b(2'b00),
    .fci(\PWM6/sub1/c1 ),
    .f(\PWM6/n26 [2:1]),
    .fco(\PWM6/sub1/c3 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM6/sub1/u0|PWM6/sub1/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM6/sub1/u4|PWM6/sub1/u3  (
    .a(pnumcnt6[4:3]),
    .b(2'b00),
    .fci(\PWM6/sub1/c3 ),
    .f(\PWM6/n26 [4:3]),
    .fco(\PWM6/sub1/c5 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM6/sub1/u0|PWM6/sub1/ucin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM6/sub1/u6|PWM6/sub1/u5  (
    .a(pnumcnt6[6:5]),
    .b(2'b00),
    .fci(\PWM6/sub1/c5 ),
    .f(\PWM6/n26 [6:5]),
    .fco(\PWM6/sub1/c7 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM6/sub1/u0|PWM6/sub1/ucin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM6/sub1/u8|PWM6/sub1/u7  (
    .a(pnumcnt6[8:7]),
    .b(2'b00),
    .fci(\PWM6/sub1/c7 ),
    .f(\PWM6/n26 [8:7]),
    .fco(\PWM6/sub1/c9 ));
  // src/OnePWM.v(26)
  // src/OnePWM.v(26)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*~(~D*B*~A))"),
    //.LUT1("(C*~(~D*B*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000010110000),
    .INIT_LUT1(16'b1111000010110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \PWM7/State_reg|PWM8/State_reg  (
    .a({_al_u3028_o,_al_u3031_o}),
    .b({\PWM7/n0_lutinv ,\PWM8/n0_lutinv }),
    .c({_al_u3029_o,_al_u3032_o}),
    .clk(clk100m),
    .d({pwm_start_stop[23],pwm_start_stop[24]}),
    .sr(rstn),
    .q({pwm_state_read[7],pwm_state_read[8]}));  // src/OnePWM.v(26)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[0]  (
    .i(\PWM7/RemaTxNum[0]_keep ),
    .o(pnumcnt7[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[10]  (
    .i(\PWM7/RemaTxNum[10]_keep ),
    .o(pnumcnt7[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[11]  (
    .i(\PWM7/RemaTxNum[11]_keep ),
    .o(pnumcnt7[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[12]  (
    .i(\PWM7/RemaTxNum[12]_keep ),
    .o(pnumcnt7[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[13]  (
    .i(\PWM7/RemaTxNum[13]_keep ),
    .o(pnumcnt7[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[14]  (
    .i(\PWM7/RemaTxNum[14]_keep ),
    .o(pnumcnt7[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[15]  (
    .i(\PWM7/RemaTxNum[15]_keep ),
    .o(pnumcnt7[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[16]  (
    .i(\PWM7/RemaTxNum[16]_keep ),
    .o(pnumcnt7[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[17]  (
    .i(\PWM7/RemaTxNum[17]_keep ),
    .o(pnumcnt7[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[18]  (
    .i(\PWM7/RemaTxNum[18]_keep ),
    .o(pnumcnt7[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[19]  (
    .i(\PWM7/RemaTxNum[19]_keep ),
    .o(pnumcnt7[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[1]  (
    .i(\PWM7/RemaTxNum[1]_keep ),
    .o(pnumcnt7[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[20]  (
    .i(\PWM7/RemaTxNum[20]_keep ),
    .o(pnumcnt7[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[21]  (
    .i(\PWM7/RemaTxNum[21]_keep ),
    .o(pnumcnt7[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[22]  (
    .i(\PWM7/RemaTxNum[22]_keep ),
    .o(pnumcnt7[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[23]  (
    .i(\PWM7/RemaTxNum[23]_keep ),
    .o(pnumcnt7[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[2]  (
    .i(\PWM7/RemaTxNum[2]_keep ),
    .o(pnumcnt7[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[3]  (
    .i(\PWM7/RemaTxNum[3]_keep ),
    .o(pnumcnt7[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[4]  (
    .i(\PWM7/RemaTxNum[4]_keep ),
    .o(pnumcnt7[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[5]  (
    .i(\PWM7/RemaTxNum[5]_keep ),
    .o(pnumcnt7[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[6]  (
    .i(\PWM7/RemaTxNum[6]_keep ),
    .o(pnumcnt7[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[7]  (
    .i(\PWM7/RemaTxNum[7]_keep ),
    .o(pnumcnt7[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[8]  (
    .i(\PWM7/RemaTxNum[8]_keep ),
    .o(pnumcnt7[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[9]  (
    .i(\PWM7/RemaTxNum[9]_keep ),
    .o(pnumcnt7[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_dir  (
    .i(\PWM7/dir_keep ),
    .o(dir_pad[7]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[0]  (
    .i(\PWM7/pnumr[0]_keep ),
    .o(\PWM7/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[10]  (
    .i(\PWM7/pnumr[10]_keep ),
    .o(\PWM7/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[11]  (
    .i(\PWM7/pnumr[11]_keep ),
    .o(\PWM7/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[12]  (
    .i(\PWM7/pnumr[12]_keep ),
    .o(\PWM7/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[13]  (
    .i(\PWM7/pnumr[13]_keep ),
    .o(\PWM7/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[14]  (
    .i(\PWM7/pnumr[14]_keep ),
    .o(\PWM7/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[15]  (
    .i(\PWM7/pnumr[15]_keep ),
    .o(\PWM7/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[16]  (
    .i(\PWM7/pnumr[16]_keep ),
    .o(\PWM7/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[17]  (
    .i(\PWM7/pnumr[17]_keep ),
    .o(\PWM7/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[18]  (
    .i(\PWM7/pnumr[18]_keep ),
    .o(\PWM7/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[19]  (
    .i(\PWM7/pnumr[19]_keep ),
    .o(\PWM7/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[1]  (
    .i(\PWM7/pnumr[1]_keep ),
    .o(\PWM7/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[20]  (
    .i(\PWM7/pnumr[20]_keep ),
    .o(\PWM7/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[21]  (
    .i(\PWM7/pnumr[21]_keep ),
    .o(\PWM7/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[22]  (
    .i(\PWM7/pnumr[22]_keep ),
    .o(\PWM7/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[23]  (
    .i(\PWM7/pnumr[23]_keep ),
    .o(\PWM7/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[24]  (
    .i(\PWM7/pnumr[24]_keep ),
    .o(\PWM7/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[25]  (
    .i(\PWM7/pnumr[25]_keep ),
    .o(\PWM7/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[26]  (
    .i(\PWM7/pnumr[26]_keep ),
    .o(\PWM7/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[27]  (
    .i(\PWM7/pnumr[27]_keep ),
    .o(\PWM7/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[28]  (
    .i(\PWM7/pnumr[28]_keep ),
    .o(\PWM7/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[29]  (
    .i(\PWM7/pnumr[29]_keep ),
    .o(\PWM7/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[2]  (
    .i(\PWM7/pnumr[2]_keep ),
    .o(\PWM7/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[30]  (
    .i(\PWM7/pnumr[30]_keep ),
    .o(\PWM7/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[31]  (
    .i(\PWM7/pnumr[31]_keep ),
    .o(\PWM7/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[3]  (
    .i(\PWM7/pnumr[3]_keep ),
    .o(\PWM7/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[4]  (
    .i(\PWM7/pnumr[4]_keep ),
    .o(\PWM7/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[5]  (
    .i(\PWM7/pnumr[5]_keep ),
    .o(\PWM7/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[6]  (
    .i(\PWM7/pnumr[6]_keep ),
    .o(\PWM7/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[7]  (
    .i(\PWM7/pnumr[7]_keep ),
    .o(\PWM7/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[8]  (
    .i(\PWM7/pnumr[8]_keep ),
    .o(\PWM7/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[9]  (
    .i(\PWM7/pnumr[9]_keep ),
    .o(\PWM7/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pwm  (
    .i(\PWM7/pwm_keep ),
    .o(pwm_pad[7]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_stopreq  (
    .i(\PWM7/stopreq_keep ),
    .o(\PWM7/stopreq ));  // src/OnePWM.v(14)
  EF2_PHY_MSLICE #(
    //.LUT0("~(~0*~(D*C*B*A))"),
    //.LUT1("~(~1*~(D*C*B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b1111111111111111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM7/pwm_reg  (
    .a({_al_u1485_o,_al_u1485_o}),
    .b({_al_u1492_o,_al_u1492_o}),
    .c({_al_u1494_o,_al_u1494_o}),
    .clk(clk100m),
    .d({_al_u1496_o,_al_u1496_o}),
    .mi({open_n11810,pwm_pad[7]}),
    .sr(\PWM7/u14_sel_is_1_o ),
    .q({open_n11816,\PWM7/pwm_keep }));  // src/OnePWM.v(45)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM7/reg0_b0|PWM7/reg0_b15  (
    .b({\PWM7/n12 [0],\PWM7/n12 [15]}),
    .c({freq7[0],freq7[15]}),
    .clk(clk100m),
    .d({\PWM7/n0_lutinv ,\PWM7/n0_lutinv }),
    .sr(\PWM7/n11 ),
    .q({\PWM7/FreCnt [0],\PWM7/FreCnt [15]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM7/reg0_b10|PWM7/reg0_b12  (
    .b({\PWM7/n12 [10],\PWM7/n12 [12]}),
    .c({freq7[10],freq7[12]}),
    .clk(clk100m),
    .d({\PWM7/n0_lutinv ,\PWM7/n0_lutinv }),
    .sr(\PWM7/n11 ),
    .q({\PWM7/FreCnt [10],\PWM7/FreCnt [12]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM7/reg0_b11|PWM7/reg0_b1  (
    .b({\PWM7/n12 [11],\PWM7/n12 [1]}),
    .c({freq7[11],freq7[1]}),
    .clk(clk100m),
    .d({\PWM7/n0_lutinv ,\PWM7/n0_lutinv }),
    .sr(\PWM7/n11 ),
    .q({\PWM7/FreCnt [11],\PWM7/FreCnt [1]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM7/reg0_b13|PWM7/reg0_b7  (
    .b({\PWM7/n12 [13],\PWM7/n12 [7]}),
    .c({freq7[13],freq7[7]}),
    .clk(clk100m),
    .d({\PWM7/n0_lutinv ,\PWM7/n0_lutinv }),
    .sr(\PWM7/n11 ),
    .q({\PWM7/FreCnt [13],\PWM7/FreCnt [7]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM7/reg0_b14|PWM7/reg0_b5  (
    .b({\PWM7/n12 [14],\PWM7/n12 [5]}),
    .c({freq7[14],freq7[5]}),
    .clk(clk100m),
    .d({\PWM7/n0_lutinv ,\PWM7/n0_lutinv }),
    .sr(\PWM7/n11 ),
    .q({\PWM7/FreCnt [14],\PWM7/FreCnt [5]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM7/reg0_b16|PWM7/reg0_b3  (
    .b({\PWM7/n12 [16],\PWM7/n12 [3]}),
    .c({freq7[16],freq7[3]}),
    .clk(clk100m),
    .d({\PWM7/n0_lutinv ,\PWM7/n0_lutinv }),
    .sr(\PWM7/n11 ),
    .q({\PWM7/FreCnt [16],\PWM7/FreCnt [3]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM7/reg0_b17|PWM7/reg0_b23  (
    .b({\PWM7/n12 [17],\PWM7/n12 [23]}),
    .c({freq7[17],freq7[23]}),
    .clk(clk100m),
    .d({\PWM7/n0_lutinv ,\PWM7/n0_lutinv }),
    .sr(\PWM7/n11 ),
    .q({\PWM7/FreCnt [17],\PWM7/FreCnt [23]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM7/reg0_b18|PWM7/reg0_b21  (
    .b({\PWM7/n12 [18],\PWM7/n12 [21]}),
    .c({freq7[18],freq7[21]}),
    .clk(clk100m),
    .d({\PWM7/n0_lutinv ,\PWM7/n0_lutinv }),
    .sr(\PWM7/n11 ),
    .q({\PWM7/FreCnt [18],\PWM7/FreCnt [21]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM7/reg0_b19|PWM7/reg0_b2  (
    .b({\PWM7/n12 [19],\PWM7/n12 [2]}),
    .c({freq7[19],freq7[2]}),
    .clk(clk100m),
    .d({\PWM7/n0_lutinv ,\PWM7/n0_lutinv }),
    .sr(\PWM7/n11 ),
    .q({\PWM7/FreCnt [19],\PWM7/FreCnt [2]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM7/reg0_b20|PWM7/reg0_b9  (
    .b({\PWM7/n12 [20],\PWM7/n12 [9]}),
    .c({freq7[20],freq7[9]}),
    .clk(clk100m),
    .d({\PWM7/n0_lutinv ,\PWM7/n0_lutinv }),
    .sr(\PWM7/n11 ),
    .q({\PWM7/FreCnt [20],\PWM7/FreCnt [9]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM7/reg0_b22|PWM7/reg0_b8  (
    .b({\PWM7/n12 [22],\PWM7/n12 [8]}),
    .c({freq7[22],freq7[8]}),
    .clk(clk100m),
    .d({\PWM7/n0_lutinv ,\PWM7/n0_lutinv }),
    .sr(\PWM7/n11 ),
    .q({\PWM7/FreCnt [22],\PWM7/FreCnt [8]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM7/reg0_b24|PWM7/reg0_b6  (
    .b({\PWM7/n12 [24],\PWM7/n12 [6]}),
    .c({freq7[24],freq7[6]}),
    .clk(clk100m),
    .d({\PWM7/n0_lutinv ,\PWM7/n0_lutinv }),
    .sr(\PWM7/n11 ),
    .q({\PWM7/FreCnt [24],\PWM7/FreCnt [6]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM7/reg0_b25|PWM7/reg0_b4  (
    .b({\PWM7/n12 [25],\PWM7/n12 [4]}),
    .c({freq7[25],freq7[4]}),
    .clk(clk100m),
    .d({\PWM7/n0_lutinv ,\PWM7/n0_lutinv }),
    .sr(\PWM7/n11 ),
    .q({\PWM7/FreCnt [25],\PWM7/FreCnt [4]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~(C@B)*~(D@A))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~(C@B)*~(D@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1000001001000001),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1000001001000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg1_b10|PWM7/reg1_b0  (
    .a({\PWM7/FreCnt [24],open_n12097}),
    .b({\PWM7/FreCnt [9],open_n12098}),
    .c({\PWM7/FreCntr [10],\PWM7/n11 }),
    .ce(\PWM7/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM7/FreCntr [25],\PWM7/n0_lutinv }),
    .mi({freq7[10],freq7[0]}),
    .f({_al_u2320_o,\PWM7/mux3_b0_sel_is_3_o }),
    .q({\PWM7/FreCntr [10],\PWM7/FreCntr [0]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~B*~(0@C)*~(~D*A))"),
    //.LUTF1("(A*~(0*~C)*~(D*~B))"),
    //.LUTG0("(~B*~(1@C)*~(~D*A))"),
    //.LUTG1("(A*~(1*~C)*~(D*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001100000001),
    .INIT_LUTF1(16'b1000100010101010),
    .INIT_LUTG0(16'b0011000000010000),
    .INIT_LUTG1(16'b1000000010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg1_b11|PWM7/reg1_b14  (
    .a({_al_u2331_o,\PWM7/FreCnt [13]}),
    .b({\PWM7/FreCnt [10],\PWM7/FreCnt [26]}),
    .c({\PWM7/FreCnt [13],\PWM7/FreCnt [8]}),
    .ce(\PWM7/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM7/FreCntr [11],\PWM7/FreCntr [14]}),
    .e({\PWM7/FreCntr [14],\PWM7/FreCntr [9]}),
    .mi({freq7[11],freq7[14]}),
    .f({_al_u2332_o,_al_u2326_o}),
    .q({\PWM7/FreCntr [11],\PWM7/FreCntr [14]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(~0*C)*~(D*~B))"),
    //.LUTF1("(~(~D*B)*~(~C*A))"),
    //.LUTG0("(A*~(~1*C)*~(D*~B))"),
    //.LUTG1("(~(~D*B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000001010),
    .INIT_LUTF1(16'b1111010100110001),
    .INIT_LUTG0(16'b1000100010101010),
    .INIT_LUTG1(16'b1111010100110001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg1_b12|PWM7/reg1_b22  (
    .a({\PWM7/FreCnt [11],_al_u2317_o}),
    .b({\PWM7/FreCnt [21],\PWM7/FreCnt [21]}),
    .c({\PWM7/FreCntr [12],\PWM7/FreCnt [23]}),
    .ce(\PWM7/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM7/FreCntr [22],\PWM7/FreCntr [22]}),
    .e({open_n12133,\PWM7/FreCntr [24]}),
    .mi({freq7[12],freq7[22]}),
    .f({_al_u2331_o,_al_u2318_o}),
    .q({\PWM7/FreCntr [12],\PWM7/FreCntr [22]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(D*~B)*~(C*~A))"),
    //.LUTF1("(B*A*~(D@C))"),
    //.LUTG0("(~(D*~B)*~(C*~A))"),
    //.LUTG1("(B*A*~(D@C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000110010101111),
    .INIT_LUTF1(16'b1000000000001000),
    .INIT_LUTG0(16'b1000110010101111),
    .INIT_LUTG1(16'b1000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg1_b15|PWM7/reg1_b13  (
    .a({_al_u2312_o,\PWM7/FreCnt [12]}),
    .b({_al_u2313_o,\PWM7/FreCnt [17]}),
    .c({\PWM7/FreCnt [14],\PWM7/FreCntr [13]}),
    .ce(\PWM7/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM7/FreCntr [15],\PWM7/FreCntr [18]}),
    .mi({freq7[15],freq7[13]}),
    .f({_al_u2314_o,_al_u2317_o}),
    .q({\PWM7/FreCntr [15],\PWM7/FreCntr [13]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*~C)*~(D*~B))"),
    //.LUTF1("(~(~D*B)*~(~C*A))"),
    //.LUTG0("(A*~(1*~C)*~(D*~B))"),
    //.LUTG1("(~(~D*B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000100010101010),
    .INIT_LUTF1(16'b1111010100110001),
    .INIT_LUTG0(16'b1000000010100000),
    .INIT_LUTG1(16'b1111010100110001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg1_b16|PWM7/reg1_b4  (
    .a({\PWM7/FreCnt [15],_al_u2328_o}),
    .b({\PWM7/FreCnt [3],\PWM7/FreCnt [3]}),
    .c({\PWM7/FreCntr [16],\PWM7/FreCnt [7]}),
    .ce(\PWM7/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM7/FreCntr [4],\PWM7/FreCntr [4]}),
    .e({open_n12168,\PWM7/FreCntr [8]}),
    .mi({freq7[16],freq7[4]}),
    .f({_al_u2313_o,_al_u2329_o}),
    .q({\PWM7/FreCntr [16],\PWM7/FreCntr [4]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~A*~(0@C)*~(~D*B))"),
    //.LUTF1("(~(D*~B)*~(~C*A))"),
    //.LUTG0("(~A*~(1@C)*~(~D*B))"),
    //.LUTG1("(~(D*~B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010100000001),
    .INIT_LUTF1(16'b1100010011110101),
    .INIT_LUTG0(16'b0101000000010000),
    .INIT_LUTG1(16'b1100010011110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg1_b18|PWM7/reg1_b24  (
    .a({\PWM7/FreCnt [17],_al_u1489_o}),
    .b({\PWM7/FreCnt [23],\PWM7/FreCnt [12]}),
    .c({\PWM7/FreCntr [18],\PWM7/FreCnt [24]}),
    .ce(\PWM7/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM7/FreCntr [24],\PWM7/FreCntr [12]}),
    .e({open_n12185,\PWM7/FreCntr [24]}),
    .mi({freq7[18],freq7[24]}),
    .f({_al_u2324_o,_al_u1490_o}),
    .q({\PWM7/FreCntr [18],\PWM7/FreCntr [24]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*~C)*~(~D*B))"),
    //.LUTF1("(~(~D*B)*~(~C*A))"),
    //.LUTG0("(A*~(1*~C)*~(~D*B))"),
    //.LUTG1("(~(~D*B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101000100010),
    .INIT_LUTF1(16'b1111010100110001),
    .INIT_LUTG0(16'b1010000000100000),
    .INIT_LUTG1(16'b1111010100110001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg1_b20|PWM7/reg1_b2  (
    .a({\PWM7/FreCnt [10],_al_u2324_o}),
    .b({\PWM7/FreCnt [19],\PWM7/FreCnt [1]}),
    .c({\PWM7/FreCntr [11],\PWM7/FreCnt [19]}),
    .ce(\PWM7/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM7/FreCntr [20],\PWM7/FreCntr [2]}),
    .e({open_n12202,\PWM7/FreCntr [20]}),
    .mi({freq7[20],freq7[2]}),
    .f({_al_u2315_o,_al_u2325_o}),
    .q({\PWM7/FreCntr [20],\PWM7/FreCntr [2]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(D@B)*~(C@A))"),
    //.LUT1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000010000100001),
    .INIT_LUT1(16'b1000010000100001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg1_b21|PWM7/reg1_b25  (
    .a({\PWM7/FreCnt [20],\PWM7/FreCnt [11]}),
    .b({\PWM7/FreCnt [6],\PWM7/FreCnt [25]}),
    .c({\PWM7/FreCntr [21],\PWM7/FreCntr [11]}),
    .ce(\PWM7/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM7/FreCntr [7],\PWM7/FreCntr [25]}),
    .mi({freq7[21],freq7[25]}),
    .f({_al_u2322_o,_al_u1493_o}),
    .q({\PWM7/FreCntr [21],\PWM7/FreCntr [25]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(D*~(C@B))"),
    //.LUTF1("(D*~(C@B))"),
    //.LUTG0("(D*~(C@B))"),
    //.LUTG1("(D*~(C@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100001100000000),
    .INIT_LUTF1(16'b1100001100000000),
    .INIT_LUTG0(16'b1100001100000000),
    .INIT_LUTG1(16'b1100001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg1_b23|PWM7/reg1_b5  (
    .b({\PWM7/FreCnt [22],\PWM7/FreCnt [4]}),
    .c({\PWM7/FreCntr [23],\PWM7/FreCntr [5]}),
    .ce(\PWM7/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({_al_u2320_o,_al_u2311_o}),
    .mi({freq7[23],freq7[5]}),
    .f({_al_u2321_o,_al_u2312_o}),
    .q({\PWM7/FreCntr [23],\PWM7/FreCntr [5]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg1_b26|PWM7/reg1_b19  (
    .a({\PWM7/FreCnt [16],_al_u2322_o}),
    .b({\PWM7/FreCnt [26],\PWM7/FreCnt [18]}),
    .c({\PWM7/FreCntr [16],\PWM7/FreCnt [25]}),
    .ce(\PWM7/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM7/FreCntr [26],\PWM7/FreCntr [19]}),
    .e({open_n12253,\PWM7/FreCntr [26]}),
    .mi({freq7[26],freq7[19]}),
    .f({_al_u1495_o,_al_u2323_o}),
    .q({\PWM7/FreCntr [26],\PWM7/FreCntr [19]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*~C)*~(~D*B))"),
    //.LUTF1("(~(~D*B)*~(~C*A))"),
    //.LUTG0("(A*~(1*~C)*~(~D*B))"),
    //.LUTG1("(~(~D*B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101000100010),
    .INIT_LUTF1(16'b1111010100110001),
    .INIT_LUTG0(16'b1010000000100000),
    .INIT_LUTG1(16'b1111010100110001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg1_b3|PWM7/reg1_b6  (
    .a({\PWM7/FreCnt [2],_al_u2315_o}),
    .b({\PWM7/FreCnt [5],\PWM7/FreCnt [12]}),
    .c({\PWM7/FreCntr [3],\PWM7/FreCnt [5]}),
    .ce(\PWM7/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM7/FreCntr [6],\PWM7/FreCntr [13]}),
    .e({open_n12270,\PWM7/FreCntr [6]}),
    .mi({freq7[3],freq7[6]}),
    .f({_al_u2328_o,_al_u2316_o}),
    .q({\PWM7/FreCntr [3],\PWM7/FreCntr [6]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg1_b7|PWM7/reg1_b9  (
    .a({\PWM7/FreCnt [6],_al_u1482_o}),
    .b({\PWM7/FreCnt [7],\PWM7/FreCnt [4]}),
    .c({\PWM7/FreCntr [6],\PWM7/FreCnt [9]}),
    .ce(\PWM7/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM7/FreCntr [7],\PWM7/FreCntr [4]}),
    .e({open_n12287,\PWM7/FreCntr [9]}),
    .mi({freq7[7],freq7[9]}),
    .f({_al_u1482_o,_al_u1483_o}),
    .q({\PWM7/FreCntr [7],\PWM7/FreCntr [9]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~A*~(0*~C)*~(D@B))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~A*~(1*~C)*~(D@B))"),
    //.LUTG1("(~C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100010000010001),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0100000000010000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg1_b8|PWM7/reg1_b1  (
    .a({open_n12304,_al_u2333_o}),
    .b({open_n12305,\PWM7/FreCnt [0]}),
    .c({\PWM7/FreCntr [8],\PWM7/FreCnt [11]}),
    .ce(\PWM7/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM7/FreCnt [7],\PWM7/FreCntr [1]}),
    .e({open_n12306,\PWM7/FreCntr [12]}),
    .mi({freq7[8],freq7[1]}),
    .f({_al_u2333_o,_al_u2334_o}),
    .q({\PWM7/FreCntr [8],\PWM7/FreCntr [1]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011100010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011100010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg2_b0|PWM7/reg2_b8  (
    .a({\PWM7/pnumr [0],\PWM7/pnumr [8]}),
    .b({pnum7[0],pnum7[32]}),
    .c({pnum7[32],pnum7[8]}),
    .clk(clk100m),
    .d({pwm_start_stop[23],pwm_start_stop[23]}),
    .q({\PWM7/pnumr[0]_keep ,\PWM7/pnumr[8]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011100010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011100010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg2_b10|PWM7/reg2_b7  (
    .a({\PWM7/pnumr [10],\PWM7/pnumr [7]}),
    .b({pnum7[10],pnum7[32]}),
    .c({pnum7[32],pnum7[7]}),
    .clk(clk100m),
    .d({pwm_start_stop[23],pwm_start_stop[23]}),
    .q({\PWM7/pnumr[10]_keep ,\PWM7/pnumr[7]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg2_b11|PWM7/reg3_b11  (
    .a({\PWM7/pnumr [11],_al_u2303_o}),
    .b({pnum7[11],\PWM7/n24 }),
    .c({pnum7[32],pnumcnt7[11]}),
    .clk(clk100m),
    .d({pwm_start_stop[23],\PWM7/pnumr [11]}),
    .e({open_n12370,pwm_start_stop[23]}),
    .q({\PWM7/pnumr[11]_keep ,\PWM7/RemaTxNum[11]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg2_b12|PWM7/reg3_b12  (
    .a({\PWM7/pnumr [12],_al_u2301_o}),
    .b({pnum7[12],\PWM7/n24 }),
    .c({pnum7[32],pnumcnt7[12]}),
    .clk(clk100m),
    .d({pwm_start_stop[23],\PWM7/pnumr [12]}),
    .e({open_n12392,pwm_start_stop[23]}),
    .q({\PWM7/pnumr[12]_keep ,\PWM7/RemaTxNum[12]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011100010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg2_b13|PWM7/reg2_b4  (
    .a({\PWM7/pnumr [13],\PWM7/pnumr [4]}),
    .b({pnum7[13],pnum7[32]}),
    .c({pnum7[32],pnum7[4]}),
    .clk(clk100m),
    .d({pwm_start_stop[23],pwm_start_stop[23]}),
    .q({\PWM7/pnumr[13]_keep ,\PWM7/pnumr[4]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg2_b14|PWM7/reg2_b3  (
    .a({\PWM7/pnumr [14],\PWM7/pnumr [3]}),
    .b({pnum7[14],pnum7[3]}),
    .c({pnum7[32],pnum7[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[23],pwm_start_stop[23]}),
    .q({\PWM7/pnumr[14]_keep ,\PWM7/pnumr[3]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg2_b15|PWM7/reg3_b15  (
    .a({\PWM7/pnumr [15],_al_u2295_o}),
    .b({pnum7[15],\PWM7/n24 }),
    .c({pnum7[32],pnumcnt7[15]}),
    .clk(clk100m),
    .d({pwm_start_stop[23],\PWM7/pnumr [15]}),
    .e({open_n12452,pwm_start_stop[23]}),
    .q({\PWM7/pnumr[15]_keep ,\PWM7/RemaTxNum[15]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg2_b16|PWM7/reg3_b16  (
    .a({\PWM7/pnumr [16],_al_u2293_o}),
    .b({pnum7[16],\PWM7/n24 }),
    .c({pnum7[32],pnumcnt7[16]}),
    .clk(clk100m),
    .d({pwm_start_stop[23],\PWM7/pnumr [16]}),
    .e({open_n12474,pwm_start_stop[23]}),
    .q({\PWM7/pnumr[16]_keep ,\PWM7/RemaTxNum[16]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg2_b17|PWM7/reg2_b21  (
    .a({\PWM7/pnumr [17],\PWM7/pnumr [21]}),
    .b({pnum7[17],pnum7[21]}),
    .c({pnum7[32],pnum7[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[23],pwm_start_stop[23]}),
    .q({\PWM7/pnumr[17]_keep ,\PWM7/pnumr[21]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg2_b18|PWM7/reg2_b20  (
    .a({\PWM7/pnumr [18],\PWM7/pnumr [20]}),
    .b({pnum7[18],pnum7[20]}),
    .c({pnum7[32],pnum7[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[23],pwm_start_stop[23]}),
    .q({\PWM7/pnumr[18]_keep ,\PWM7/pnumr[20]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg2_b19|PWM7/reg3_b19  (
    .a({\PWM7/pnumr [19],_al_u2287_o}),
    .b({pnum7[19],\PWM7/n24 }),
    .c({pnum7[32],pnumcnt7[19]}),
    .clk(clk100m),
    .d({pwm_start_stop[23],\PWM7/pnumr [19]}),
    .e({open_n12542,pwm_start_stop[23]}),
    .q({\PWM7/pnumr[19]_keep ,\PWM7/RemaTxNum[19]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg2_b22|PWM7/reg3_b22  (
    .a({\PWM7/pnumr [22],_al_u2279_o}),
    .b({pnum7[22],\PWM7/n24 }),
    .c({pnum7[32],pnumcnt7[22]}),
    .clk(clk100m),
    .d({pwm_start_stop[23],\PWM7/pnumr [22]}),
    .e({open_n12564,pwm_start_stop[23]}),
    .q({\PWM7/pnumr[22]_keep ,\PWM7/RemaTxNum[22]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg2_b23|PWM7/reg3_b23  (
    .a({\PWM7/pnumr [23],_al_u2277_o}),
    .b({pnum7[23],\PWM7/n24 }),
    .c({pnum7[32],pnumcnt7[23]}),
    .clk(clk100m),
    .d({pwm_start_stop[23],\PWM7/pnumr [23]}),
    .e({open_n12586,pwm_start_stop[23]}),
    .q({\PWM7/pnumr[23]_keep ,\PWM7/RemaTxNum[23]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg2_b24|PWM7/reg2_b30  (
    .a({\PWM7/pnumr [24],\PWM7/pnumr [30]}),
    .b({pnum7[24],pnum7[30]}),
    .c({pnum7[32],pnum7[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[23],pwm_start_stop[23]}),
    .q({\PWM7/pnumr[24]_keep ,\PWM7/pnumr[30]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg2_b25|PWM7/reg2_b29  (
    .a({\PWM7/pnumr [25],\PWM7/pnumr [29]}),
    .b({pnum7[25],pnum7[29]}),
    .c({pnum7[32],pnum7[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[23],pwm_start_stop[23]}),
    .q({\PWM7/pnumr[25]_keep ,\PWM7/pnumr[29]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg2_b26|PWM7/reg2_b28  (
    .a({\PWM7/pnumr [26],\PWM7/pnumr [28]}),
    .b({pnum7[26],pnum7[28]}),
    .c({pnum7[32],pnum7[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[23],pwm_start_stop[23]}),
    .q({\PWM7/pnumr[26]_keep ,\PWM7/pnumr[28]_keep }));  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg2_b27  (
    .a({open_n12668,\PWM7/pnumr [27]}),
    .b({open_n12669,pnum7[27]}),
    .c({open_n12670,pnum7[32]}),
    .clk(clk100m),
    .d({open_n12672,pwm_start_stop[23]}),
    .q({open_n12695,\PWM7/pnumr[27]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg2_b2|PWM7/reg3_b2  (
    .a({\PWM7/pnumr [2],_al_u2285_o}),
    .b({pnum7[2],\PWM7/n24 }),
    .c({pnum7[32],pnumcnt7[2]}),
    .clk(clk100m),
    .d({pwm_start_stop[23],\PWM7/pnumr [2]}),
    .e({open_n12697,pwm_start_stop[23]}),
    .q({\PWM7/pnumr[2]_keep ,\PWM7/RemaTxNum[2]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(D*~(C)*~((~0*~(B*A)))+D*C*~((~0*~(B*A)))+~(D)*C*(~0*~(B*A))+D*C*(~0*~(B*A)))"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(D*~(C)*~((~1*~(B*A)))+D*C*~((~1*~(B*A)))+~(D)*C*(~1*~(B*A))+D*C*(~1*~(B*A)))"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111100001110000),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg2_b31|PWM7/dir_reg  (
    .a({\PWM7/pnumr [31],\PWM7/n24 }),
    .b({pnum7[31],\PWM7/n25_neg_lutinv }),
    .c({pnum7[32],dir_pad[7]}),
    .clk(clk100m),
    .d({pwm_start_stop[23],\PWM7/pnumr [31]}),
    .e({open_n12719,pwm_start_stop[23]}),
    .q({\PWM7/pnumr[31]_keep ,\PWM7/dir_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg2_b5|PWM7/reg3_b5  (
    .a({\PWM7/pnumr [5],_al_u2271_o}),
    .b({pnum7[32],\PWM7/n24 }),
    .c({pnum7[5],pnumcnt7[5]}),
    .clk(clk100m),
    .d({pwm_start_stop[23],\PWM7/pnumr [5]}),
    .e({open_n12741,pwm_start_stop[23]}),
    .q({\PWM7/pnumr[5]_keep ,\PWM7/RemaTxNum[5]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg2_b6|PWM7/reg3_b6  (
    .a({\PWM7/pnumr [6],_al_u2269_o}),
    .b({pnum7[32],\PWM7/n24 }),
    .c({pnum7[6],pnumcnt7[6]}),
    .clk(clk100m),
    .d({pwm_start_stop[23],\PWM7/pnumr [6]}),
    .e({open_n12763,pwm_start_stop[23]}),
    .q({\PWM7/pnumr[6]_keep ,\PWM7/RemaTxNum[6]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg2_b9|PWM7/reg3_b9  (
    .a({\PWM7/pnumr [9],_al_u2263_o}),
    .b({pnum7[32],\PWM7/n24 }),
    .c({pnum7[9],pnumcnt7[9]}),
    .clk(clk100m),
    .d({pwm_start_stop[23],\PWM7/pnumr [9]}),
    .e({open_n12785,pwm_start_stop[23]}),
    .q({\PWM7/pnumr[9]_keep ,\PWM7/RemaTxNum[9]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg3_b1  (
    .a({_al_u2307_o,_al_u2307_o}),
    .b({\PWM7/n24 ,\PWM7/n24 }),
    .c({pnumcnt7[1],pnumcnt7[1]}),
    .clk(clk100m),
    .d({\PWM7/pnumr [1],\PWM7/pnumr [1]}),
    .mi({open_n12817,pwm_start_stop[23]}),
    .q({open_n12824,\PWM7/RemaTxNum[1]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg3_b10  (
    .a({_al_u2305_o,_al_u2305_o}),
    .b({\PWM7/n24 ,\PWM7/n24 }),
    .c({pnumcnt7[10],pnumcnt7[10]}),
    .clk(clk100m),
    .d({\PWM7/pnumr [10],\PWM7/pnumr [10]}),
    .mi({open_n12836,pwm_start_stop[23]}),
    .q({open_n12843,\PWM7/RemaTxNum[10]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg3_b13  (
    .a({_al_u2299_o,_al_u2299_o}),
    .b({\PWM7/n24 ,\PWM7/n24 }),
    .c({pnumcnt7[13],pnumcnt7[13]}),
    .clk(clk100m),
    .d({\PWM7/pnumr [13],\PWM7/pnumr [13]}),
    .mi({open_n12855,pwm_start_stop[23]}),
    .q({open_n12862,\PWM7/RemaTxNum[13]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg3_b14  (
    .a({_al_u2297_o,_al_u2297_o}),
    .b({\PWM7/n24 ,\PWM7/n24 }),
    .c({pnumcnt7[14],pnumcnt7[14]}),
    .clk(clk100m),
    .d({\PWM7/pnumr [14],\PWM7/pnumr [14]}),
    .mi({open_n12874,pwm_start_stop[23]}),
    .q({open_n12881,\PWM7/RemaTxNum[14]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg3_b17  (
    .a({_al_u2291_o,_al_u2291_o}),
    .b({\PWM7/n24 ,\PWM7/n24 }),
    .c({pnumcnt7[17],pnumcnt7[17]}),
    .clk(clk100m),
    .d({\PWM7/pnumr [17],\PWM7/pnumr [17]}),
    .mi({open_n12893,pwm_start_stop[23]}),
    .q({open_n12900,\PWM7/RemaTxNum[17]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg3_b18  (
    .a({_al_u2289_o,_al_u2289_o}),
    .b({\PWM7/n24 ,\PWM7/n24 }),
    .c({pnumcnt7[18],pnumcnt7[18]}),
    .clk(clk100m),
    .d({\PWM7/pnumr [18],\PWM7/pnumr [18]}),
    .mi({open_n12912,pwm_start_stop[23]}),
    .q({open_n12919,\PWM7/RemaTxNum[18]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg3_b20  (
    .a({_al_u2283_o,_al_u2283_o}),
    .b({\PWM7/n24 ,\PWM7/n24 }),
    .c({pnumcnt7[20],pnumcnt7[20]}),
    .clk(clk100m),
    .d({\PWM7/pnumr [20],\PWM7/pnumr [20]}),
    .mi({open_n12931,pwm_start_stop[23]}),
    .q({open_n12938,\PWM7/RemaTxNum[20]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg3_b21  (
    .a({_al_u2281_o,_al_u2281_o}),
    .b({\PWM7/n24 ,\PWM7/n24 }),
    .c({pnumcnt7[21],pnumcnt7[21]}),
    .clk(clk100m),
    .d({\PWM7/pnumr [21],\PWM7/pnumr [21]}),
    .mi({open_n12950,pwm_start_stop[23]}),
    .q({open_n12957,\PWM7/RemaTxNum[21]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg3_b3  (
    .a({_al_u2275_o,_al_u2275_o}),
    .b({\PWM7/n24 ,\PWM7/n24 }),
    .c({pnumcnt7[3],pnumcnt7[3]}),
    .clk(clk100m),
    .d({\PWM7/pnumr [3],\PWM7/pnumr [3]}),
    .mi({open_n12969,pwm_start_stop[23]}),
    .q({open_n12976,\PWM7/RemaTxNum[3]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg3_b4  (
    .a({_al_u2273_o,_al_u2273_o}),
    .b({\PWM7/n24 ,\PWM7/n24 }),
    .c({pnumcnt7[4],pnumcnt7[4]}),
    .clk(clk100m),
    .d({\PWM7/pnumr [4],\PWM7/pnumr [4]}),
    .mi({open_n12988,pwm_start_stop[23]}),
    .q({open_n12995,\PWM7/RemaTxNum[4]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg3_b7  (
    .a({_al_u2267_o,_al_u2267_o}),
    .b({\PWM7/n24 ,\PWM7/n24 }),
    .c({pnumcnt7[7],pnumcnt7[7]}),
    .clk(clk100m),
    .d({\PWM7/pnumr [7],\PWM7/pnumr [7]}),
    .mi({open_n13007,pwm_start_stop[23]}),
    .q({open_n13014,\PWM7/RemaTxNum[7]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/reg3_b8  (
    .a({_al_u2265_o,_al_u2265_o}),
    .b({\PWM7/n24 ,\PWM7/n24 }),
    .c({pnumcnt7[8],pnumcnt7[8]}),
    .clk(clk100m),
    .d({\PWM7/pnumr [8],\PWM7/pnumr [8]}),
    .mi({open_n13026,pwm_start_stop[23]}),
    .q({open_n13033,\PWM7/RemaTxNum[8]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_LSLICE #(
    //.MACRO("PWM7/sub0/ucin_al_u3412"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM7/sub0/u11_al_u3415  (
    .a({\PWM7/FreCnt [13],\PWM7/FreCnt [11]}),
    .b({\PWM7/FreCnt [14],\PWM7/FreCnt [12]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM7/sub0/c11 ),
    .f({\PWM7/n12 [13],\PWM7/n12 [11]}),
    .fco(\PWM7/sub0/c15 ),
    .fx({\PWM7/n12 [14],\PWM7/n12 [12]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM7/sub0/ucin_al_u3412"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM7/sub0/u15_al_u3416  (
    .a({\PWM7/FreCnt [17],\PWM7/FreCnt [15]}),
    .b({\PWM7/FreCnt [18],\PWM7/FreCnt [16]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM7/sub0/c15 ),
    .f({\PWM7/n12 [17],\PWM7/n12 [15]}),
    .fco(\PWM7/sub0/c19 ),
    .fx({\PWM7/n12 [18],\PWM7/n12 [16]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM7/sub0/ucin_al_u3412"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM7/sub0/u19_al_u3417  (
    .a({\PWM7/FreCnt [21],\PWM7/FreCnt [19]}),
    .b({\PWM7/FreCnt [22],\PWM7/FreCnt [20]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM7/sub0/c19 ),
    .f({\PWM7/n12 [21],\PWM7/n12 [19]}),
    .fco(\PWM7/sub0/c23 ),
    .fx({\PWM7/n12 [22],\PWM7/n12 [20]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM7/sub0/ucin_al_u3412"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM7/sub0/u23_al_u3418  (
    .a({\PWM7/FreCnt [25],\PWM7/FreCnt [23]}),
    .b({\PWM7/FreCnt [26],\PWM7/FreCnt [24]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM7/sub0/c23 ),
    .f({\PWM7/n12 [25],\PWM7/n12 [23]}),
    .fx({\PWM7/n12 [26],\PWM7/n12 [24]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM7/sub0/ucin_al_u3412"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM7/sub0/u3_al_u3413  (
    .a({\PWM7/FreCnt [5],\PWM7/FreCnt [3]}),
    .b({\PWM7/FreCnt [6],\PWM7/FreCnt [4]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM7/sub0/c3 ),
    .f({\PWM7/n12 [5],\PWM7/n12 [3]}),
    .fco(\PWM7/sub0/c7 ),
    .fx({\PWM7/n12 [6],\PWM7/n12 [4]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM7/sub0/ucin_al_u3412"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM7/sub0/u7_al_u3414  (
    .a({\PWM7/FreCnt [9],\PWM7/FreCnt [7]}),
    .b({\PWM7/FreCnt [10],\PWM7/FreCnt [8]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM7/sub0/c7 ),
    .f({\PWM7/n12 [9],\PWM7/n12 [7]}),
    .fco(\PWM7/sub0/c11 ),
    .fx({\PWM7/n12 [10],\PWM7/n12 [8]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM7/sub0/ucin_al_u3412"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'h0005),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM7/sub0/ucin_al_u3412  (
    .a({\PWM7/FreCnt [1],1'b0}),
    .b({\PWM7/FreCnt [2],\PWM7/FreCnt [0]}),
    .c(2'b11),
    .ce(\U_AHB/n18 ),
    .clk(clk100m),
    .d(2'b01),
    .e(2'b01),
    .mi({\U_AHB/h2h_hwdata [24],\U_AHB/h2h_hwdata [2]}),
    .f({\PWM7/n12 [1],open_n13156}),
    .fco(\PWM7/sub0/c3 ),
    .fx({\PWM7/n12 [2],\PWM7/n12 [0]}),
    .q({freq7[24],freq7[2]}));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM7/sub1/u0|PWM7/sub1/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("SUB_CARRY"),
    .INIT_LUT0(16'b0000000000000101),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM7/sub1/u0|PWM7/sub1/ucin  (
    .a({pnumcnt7[0],1'b0}),
    .b({1'b1,open_n13157}),
    .f({\PWM7/n26 [0],open_n13177}),
    .fco(\PWM7/sub1/c1 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM7/sub1/u0|PWM7/sub1/ucin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM7/sub1/u10|PWM7/sub1/u9  (
    .a(pnumcnt7[10:9]),
    .b(2'b00),
    .fci(\PWM7/sub1/c9 ),
    .f(\PWM7/n26 [10:9]),
    .fco(\PWM7/sub1/c11 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM7/sub1/u0|PWM7/sub1/ucin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM7/sub1/u12|PWM7/sub1/u11  (
    .a(pnumcnt7[12:11]),
    .b(2'b00),
    .fci(\PWM7/sub1/c11 ),
    .f(\PWM7/n26 [12:11]),
    .fco(\PWM7/sub1/c13 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM7/sub1/u0|PWM7/sub1/ucin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM7/sub1/u14|PWM7/sub1/u13  (
    .a(pnumcnt7[14:13]),
    .b(2'b00),
    .fci(\PWM7/sub1/c13 ),
    .f(\PWM7/n26 [14:13]),
    .fco(\PWM7/sub1/c15 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM7/sub1/u0|PWM7/sub1/ucin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM7/sub1/u16|PWM7/sub1/u15  (
    .a(pnumcnt7[16:15]),
    .b(2'b00),
    .fci(\PWM7/sub1/c15 ),
    .f(\PWM7/n26 [16:15]),
    .fco(\PWM7/sub1/c17 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM7/sub1/u0|PWM7/sub1/ucin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM7/sub1/u18|PWM7/sub1/u17  (
    .a(pnumcnt7[18:17]),
    .b(2'b00),
    .fci(\PWM7/sub1/c17 ),
    .f(\PWM7/n26 [18:17]),
    .fco(\PWM7/sub1/c19 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM7/sub1/u0|PWM7/sub1/ucin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM7/sub1/u20|PWM7/sub1/u19  (
    .a(pnumcnt7[20:19]),
    .b(2'b00),
    .fci(\PWM7/sub1/c19 ),
    .f(\PWM7/n26 [20:19]),
    .fco(\PWM7/sub1/c21 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM7/sub1/u0|PWM7/sub1/ucin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM7/sub1/u22|PWM7/sub1/u21  (
    .a(pnumcnt7[22:21]),
    .b(2'b00),
    .fci(\PWM7/sub1/c21 ),
    .f(\PWM7/n26 [22:21]),
    .fco(\PWM7/sub1/c23 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM7/sub1/u0|PWM7/sub1/ucin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM7/sub1/u23_al_u3475  (
    .a({open_n13336,pnumcnt7[23]}),
    .b({open_n13337,1'b0}),
    .fci(\PWM7/sub1/c23 ),
    .f({open_n13356,\PWM7/n26 [23]}));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM7/sub1/u0|PWM7/sub1/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM7/sub1/u2|PWM7/sub1/u1  (
    .a(pnumcnt7[2:1]),
    .b(2'b00),
    .fci(\PWM7/sub1/c1 ),
    .f(\PWM7/n26 [2:1]),
    .fco(\PWM7/sub1/c3 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM7/sub1/u0|PWM7/sub1/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM7/sub1/u4|PWM7/sub1/u3  (
    .a(pnumcnt7[4:3]),
    .b(2'b00),
    .fci(\PWM7/sub1/c3 ),
    .f(\PWM7/n26 [4:3]),
    .fco(\PWM7/sub1/c5 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM7/sub1/u0|PWM7/sub1/ucin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM7/sub1/u6|PWM7/sub1/u5  (
    .a(pnumcnt7[6:5]),
    .b(2'b00),
    .fci(\PWM7/sub1/c5 ),
    .f(\PWM7/n26 [6:5]),
    .fco(\PWM7/sub1/c7 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM7/sub1/u0|PWM7/sub1/ucin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM7/sub1/u8|PWM7/sub1/u7  (
    .a(pnumcnt7[8:7]),
    .b(2'b00),
    .fci(\PWM7/sub1/c7 ),
    .f(\PWM7/n26 [8:7]),
    .fco(\PWM7/sub1/c9 ));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[0]  (
    .i(\PWM8/RemaTxNum[0]_keep ),
    .o(pnumcnt8[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[10]  (
    .i(\PWM8/RemaTxNum[10]_keep ),
    .o(pnumcnt8[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[11]  (
    .i(\PWM8/RemaTxNum[11]_keep ),
    .o(pnumcnt8[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[12]  (
    .i(\PWM8/RemaTxNum[12]_keep ),
    .o(pnumcnt8[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[13]  (
    .i(\PWM8/RemaTxNum[13]_keep ),
    .o(pnumcnt8[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[14]  (
    .i(\PWM8/RemaTxNum[14]_keep ),
    .o(pnumcnt8[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[15]  (
    .i(\PWM8/RemaTxNum[15]_keep ),
    .o(pnumcnt8[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[16]  (
    .i(\PWM8/RemaTxNum[16]_keep ),
    .o(pnumcnt8[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[17]  (
    .i(\PWM8/RemaTxNum[17]_keep ),
    .o(pnumcnt8[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[18]  (
    .i(\PWM8/RemaTxNum[18]_keep ),
    .o(pnumcnt8[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[19]  (
    .i(\PWM8/RemaTxNum[19]_keep ),
    .o(pnumcnt8[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[1]  (
    .i(\PWM8/RemaTxNum[1]_keep ),
    .o(pnumcnt8[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[20]  (
    .i(\PWM8/RemaTxNum[20]_keep ),
    .o(pnumcnt8[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[21]  (
    .i(\PWM8/RemaTxNum[21]_keep ),
    .o(pnumcnt8[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[22]  (
    .i(\PWM8/RemaTxNum[22]_keep ),
    .o(pnumcnt8[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[23]  (
    .i(\PWM8/RemaTxNum[23]_keep ),
    .o(pnumcnt8[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[2]  (
    .i(\PWM8/RemaTxNum[2]_keep ),
    .o(pnumcnt8[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[3]  (
    .i(\PWM8/RemaTxNum[3]_keep ),
    .o(pnumcnt8[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[4]  (
    .i(\PWM8/RemaTxNum[4]_keep ),
    .o(pnumcnt8[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[5]  (
    .i(\PWM8/RemaTxNum[5]_keep ),
    .o(pnumcnt8[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[6]  (
    .i(\PWM8/RemaTxNum[6]_keep ),
    .o(pnumcnt8[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[7]  (
    .i(\PWM8/RemaTxNum[7]_keep ),
    .o(pnumcnt8[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[8]  (
    .i(\PWM8/RemaTxNum[8]_keep ),
    .o(pnumcnt8[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[9]  (
    .i(\PWM8/RemaTxNum[9]_keep ),
    .o(pnumcnt8[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_dir  (
    .i(\PWM8/dir_keep ),
    .o(dir_pad[8]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[0]  (
    .i(\PWM8/pnumr[0]_keep ),
    .o(\PWM8/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[10]  (
    .i(\PWM8/pnumr[10]_keep ),
    .o(\PWM8/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[11]  (
    .i(\PWM8/pnumr[11]_keep ),
    .o(\PWM8/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[12]  (
    .i(\PWM8/pnumr[12]_keep ),
    .o(\PWM8/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[13]  (
    .i(\PWM8/pnumr[13]_keep ),
    .o(\PWM8/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[14]  (
    .i(\PWM8/pnumr[14]_keep ),
    .o(\PWM8/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[15]  (
    .i(\PWM8/pnumr[15]_keep ),
    .o(\PWM8/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[16]  (
    .i(\PWM8/pnumr[16]_keep ),
    .o(\PWM8/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[17]  (
    .i(\PWM8/pnumr[17]_keep ),
    .o(\PWM8/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[18]  (
    .i(\PWM8/pnumr[18]_keep ),
    .o(\PWM8/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[19]  (
    .i(\PWM8/pnumr[19]_keep ),
    .o(\PWM8/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[1]  (
    .i(\PWM8/pnumr[1]_keep ),
    .o(\PWM8/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[20]  (
    .i(\PWM8/pnumr[20]_keep ),
    .o(\PWM8/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[21]  (
    .i(\PWM8/pnumr[21]_keep ),
    .o(\PWM8/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[22]  (
    .i(\PWM8/pnumr[22]_keep ),
    .o(\PWM8/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[23]  (
    .i(\PWM8/pnumr[23]_keep ),
    .o(\PWM8/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[24]  (
    .i(\PWM8/pnumr[24]_keep ),
    .o(\PWM8/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[25]  (
    .i(\PWM8/pnumr[25]_keep ),
    .o(\PWM8/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[26]  (
    .i(\PWM8/pnumr[26]_keep ),
    .o(\PWM8/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[27]  (
    .i(\PWM8/pnumr[27]_keep ),
    .o(\PWM8/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[28]  (
    .i(\PWM8/pnumr[28]_keep ),
    .o(\PWM8/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[29]  (
    .i(\PWM8/pnumr[29]_keep ),
    .o(\PWM8/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[2]  (
    .i(\PWM8/pnumr[2]_keep ),
    .o(\PWM8/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[30]  (
    .i(\PWM8/pnumr[30]_keep ),
    .o(\PWM8/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[31]  (
    .i(\PWM8/pnumr[31]_keep ),
    .o(\PWM8/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[3]  (
    .i(\PWM8/pnumr[3]_keep ),
    .o(\PWM8/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[4]  (
    .i(\PWM8/pnumr[4]_keep ),
    .o(\PWM8/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[5]  (
    .i(\PWM8/pnumr[5]_keep ),
    .o(\PWM8/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[6]  (
    .i(\PWM8/pnumr[6]_keep ),
    .o(\PWM8/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[7]  (
    .i(\PWM8/pnumr[7]_keep ),
    .o(\PWM8/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[8]  (
    .i(\PWM8/pnumr[8]_keep ),
    .o(\PWM8/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[9]  (
    .i(\PWM8/pnumr[9]_keep ),
    .o(\PWM8/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pwm  (
    .i(\PWM8/pwm_keep ),
    .o(pwm_pad[8]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_stopreq  (
    .i(\PWM8/stopreq_keep ),
    .o(\PWM8/stopreq ));  // src/OnePWM.v(14)
  EF2_PHY_MSLICE #(
    //.LUT0("(D*~(C)*~((~0*~(B*A)))+D*C*~((~0*~(B*A)))+~(D)*C*(~0*~(B*A))+D*C*(~0*~(B*A)))"),
    //.LUT1("(D*~(C)*~((~1*~(B*A)))+D*C*~((~1*~(B*A)))+~(D)*C*(~1*~(B*A))+D*C*(~1*~(B*A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111100001110000),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/dir_reg  (
    .a({\PWM8/n24 ,\PWM8/n24 }),
    .b({\PWM8/n25_neg_lutinv ,\PWM8/n25_neg_lutinv }),
    .c({dir_pad[8],dir_pad[8]}),
    .clk(clk100m),
    .d({\PWM8/pnumr [31],\PWM8/pnumr [31]}),
    .mi({open_n13461,pwm_start_stop[24]}),
    .q({open_n13468,\PWM8/dir_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("~(~0*~(D*C*B*A))"),
    //.LUT1("~(~1*~(D*C*B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b1111111111111111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM8/pwm_reg  (
    .a({_al_u1503_o,_al_u1503_o}),
    .b({_al_u1510_o,_al_u1510_o}),
    .c({_al_u1512_o,_al_u1512_o}),
    .clk(clk100m),
    .d({_al_u1514_o,_al_u1514_o}),
    .mi({open_n13480,pwm_pad[8]}),
    .sr(\PWM8/u14_sel_is_1_o ),
    .q({open_n13486,\PWM8/pwm_keep }));  // src/OnePWM.v(45)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM8/reg0_b0|PWM8/reg0_b15  (
    .b({\PWM8/n12 [0],\PWM8/n12 [15]}),
    .c({freq8[0],freq8[15]}),
    .clk(clk100m),
    .d({\PWM8/n0_lutinv ,\PWM8/n0_lutinv }),
    .sr(\PWM8/n11 ),
    .q({\PWM8/FreCnt [0],\PWM8/FreCnt [15]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM8/reg0_b10|PWM8/reg0_b1  (
    .b({\PWM8/n12 [10],\PWM8/n12 [1]}),
    .c({freq8[10],freq8[1]}),
    .clk(clk100m),
    .d({\PWM8/n0_lutinv ,\PWM8/n0_lutinv }),
    .sr(\PWM8/n11 ),
    .q({\PWM8/FreCnt [10],\PWM8/FreCnt [1]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM8/reg0_b11|PWM8/reg0_b8  (
    .b({\PWM8/n12 [11],\PWM8/n12 [8]}),
    .c({freq8[11],freq8[8]}),
    .clk(clk100m),
    .d({\PWM8/n0_lutinv ,\PWM8/n0_lutinv }),
    .sr(\PWM8/n11 ),
    .q({\PWM8/FreCnt [11],\PWM8/FreCnt [8]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM8/reg0_b12|PWM8/reg0_b7  (
    .b({\PWM8/n12 [12],\PWM8/n12 [7]}),
    .c({freq8[12],freq8[7]}),
    .clk(clk100m),
    .d({\PWM8/n0_lutinv ,\PWM8/n0_lutinv }),
    .sr(\PWM8/n11 ),
    .q({\PWM8/FreCnt [12],\PWM8/FreCnt [7]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM8/reg0_b13|PWM8/reg0_b5  (
    .b({\PWM8/n12 [13],\PWM8/n12 [5]}),
    .c({freq8[13],freq8[5]}),
    .clk(clk100m),
    .d({\PWM8/n0_lutinv ,\PWM8/n0_lutinv }),
    .sr(\PWM8/n11 ),
    .q({\PWM8/FreCnt [13],\PWM8/FreCnt [5]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM8/reg0_b14|PWM8/reg0_b3  (
    .b({\PWM8/n12 [14],\PWM8/n12 [3]}),
    .c({freq8[14],freq8[3]}),
    .clk(clk100m),
    .d({\PWM8/n0_lutinv ,\PWM8/n0_lutinv }),
    .sr(\PWM8/n11 ),
    .q({\PWM8/FreCnt [14],\PWM8/FreCnt [3]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM8/reg0_b16|PWM8/reg0_b25  (
    .b({\PWM8/n12 [16],\PWM8/n12 [25]}),
    .c({freq8[16],freq8[25]}),
    .clk(clk100m),
    .d({\PWM8/n0_lutinv ,\PWM8/n0_lutinv }),
    .sr(\PWM8/n11 ),
    .q({\PWM8/FreCnt [16],\PWM8/FreCnt [25]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM8/reg0_b17|PWM8/reg0_b23  (
    .b({\PWM8/n12 [17],\PWM8/n12 [23]}),
    .c({freq8[17],freq8[23]}),
    .clk(clk100m),
    .d({\PWM8/n0_lutinv ,\PWM8/n0_lutinv }),
    .sr(\PWM8/n11 ),
    .q({\PWM8/FreCnt [17],\PWM8/FreCnt [23]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM8/reg0_b18|PWM8/reg0_b22  (
    .b({\PWM8/n12 [18],\PWM8/n12 [22]}),
    .c({freq8[18],freq8[22]}),
    .clk(clk100m),
    .d({\PWM8/n0_lutinv ,\PWM8/n0_lutinv }),
    .sr(\PWM8/n11 ),
    .q({\PWM8/FreCnt [18],\PWM8/FreCnt [22]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM8/reg0_b19|PWM8/reg0_b21  (
    .b({\PWM8/n12 [19],\PWM8/n12 [21]}),
    .c({freq8[19],freq8[21]}),
    .clk(clk100m),
    .d({\PWM8/n0_lutinv ,\PWM8/n0_lutinv }),
    .sr(\PWM8/n11 ),
    .q({\PWM8/FreCnt [19],\PWM8/FreCnt [21]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM8/reg0_b20|PWM8/reg0_b9  (
    .b({\PWM8/n12 [20],\PWM8/n12 [9]}),
    .c({freq8[20],freq8[9]}),
    .clk(clk100m),
    .d({\PWM8/n0_lutinv ,\PWM8/n0_lutinv }),
    .sr(\PWM8/n11 ),
    .q({\PWM8/FreCnt [20],\PWM8/FreCnt [9]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM8/reg0_b24|PWM8/reg0_b6  (
    .b({\PWM8/n12 [24],\PWM8/n12 [6]}),
    .c({freq8[24],freq8[6]}),
    .clk(clk100m),
    .d({\PWM8/n0_lutinv ,\PWM8/n0_lutinv }),
    .sr(\PWM8/n11 ),
    .q({\PWM8/FreCnt [24],\PWM8/FreCnt [6]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM8/reg0_b26|PWM8/reg0_b4  (
    .b({\PWM8/n12 [26],\PWM8/n12 [4]}),
    .c({freq8[26],freq8[4]}),
    .clk(clk100m),
    .d({\PWM8/n0_lutinv ,\PWM8/n0_lutinv }),
    .sr(\PWM8/n11 ),
    .q({\PWM8/FreCnt [26],\PWM8/FreCnt [4]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(~(C@B)*~(D@A))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(~(C@B)*~(D@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b1000001001000001),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000001001000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg1_b10|PWM8/reg1_b17  (
    .a({\PWM8/FreCnt [16],_al_u1498_o}),
    .b({\PWM8/FreCnt [9],\PWM8/FreCnt [17]}),
    .c({\PWM8/FreCntr [10],\PWM8/FreCnt [8]}),
    .ce(\PWM8/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM8/FreCntr [17],\PWM8/FreCntr [17]}),
    .e({open_n13771,\PWM8/FreCntr [8]}),
    .mi({freq8[10],freq8[17]}),
    .f({_al_u2397_o,_al_u1499_o}),
    .q({\PWM8/FreCntr [10],\PWM8/FreCntr [17]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(D*~B)*~(~C*A))"),
    //.LUT1("(B*A*~(D@C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100010011110101),
    .INIT_LUT1(16'b1000000000001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg1_b14|PWM8/reg1_b11  (
    .a({_al_u2408_o,\PWM8/FreCnt [10]}),
    .b({_al_u2409_o,\PWM8/FreCnt [5]}),
    .c({\PWM8/FreCnt [13],\PWM8/FreCntr [11]}),
    .ce(\PWM8/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM8/FreCntr [14],\PWM8/FreCntr [6]}),
    .mi({freq8[14],freq8[11]}),
    .f({_al_u2410_o,_al_u2411_o}),
    .q({\PWM8/FreCntr [14],\PWM8/FreCntr [11]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(D@B)*~(C@A))"),
    //.LUTF1("(D*~(C@B))"),
    //.LUTG0("(~(D@B)*~(C@A))"),
    //.LUTG1("(D*~(C@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000010000100001),
    .INIT_LUTF1(16'b1100001100000000),
    .INIT_LUTG0(16'b1000010000100001),
    .INIT_LUTG1(16'b1100001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg1_b1|PWM8/reg1_b19  (
    .a({open_n13802,\PWM8/FreCnt [18]}),
    .b({\PWM8/FreCnt [0],\PWM8/FreCnt [6]}),
    .c({\PWM8/FreCntr [1],\PWM8/FreCntr [19]}),
    .ce(\PWM8/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({_al_u2401_o,\PWM8/FreCntr [7]}),
    .mi({freq8[1],freq8[19]}),
    .f({_al_u2402_o,_al_u2401_o}),
    .q({\PWM8/FreCntr [1],\PWM8/FreCntr [19]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~A*~(0@C)*~(D*~B))"),
    //.LUTF1("(A*~(0@C)*~(D@B))"),
    //.LUTG0("(~A*~(1@C)*~(D*~B))"),
    //.LUTG1("(A*~(1@C)*~(D@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010000000101),
    .INIT_LUTF1(16'b0000100000000010),
    .INIT_LUTG0(16'b0100000001010000),
    .INIT_LUTG1(16'b1000000000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg1_b20|PWM8/reg1_b18  (
    .a({_al_u1511_o,_al_u2413_o}),
    .b({\PWM8/FreCnt [14],\PWM8/FreCnt [17]}),
    .c(\PWM8/FreCnt [20:19]),
    .ce(\PWM8/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM8/FreCntr [14],\PWM8/FreCntr [18]}),
    .e({\PWM8/FreCntr [20],\PWM8/FreCntr [20]}),
    .mi({freq8[20],freq8[18]}),
    .f({_al_u1512_o,_al_u2414_o}),
    .q({\PWM8/FreCntr [20],\PWM8/FreCntr [18]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(D@B)*~(C@A))"),
    //.LUTF1("(B*A*~(D@C))"),
    //.LUTG0("(~(D@B)*~(C@A))"),
    //.LUTG1("(B*A*~(D@C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000010000100001),
    .INIT_LUTF1(16'b1000000000001000),
    .INIT_LUTG0(16'b1000010000100001),
    .INIT_LUTG1(16'b1000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg1_b21|PWM8/reg1_b15  (
    .a({_al_u1504_o,\PWM8/FreCnt [14]}),
    .b({_al_u1505_o,\PWM8/FreCnt [20]}),
    .c({\PWM8/FreCnt [21],\PWM8/FreCntr [15]}),
    .ce(\PWM8/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM8/FreCntr [21],\PWM8/FreCntr [21]}),
    .mi({freq8[21],freq8[15]}),
    .f({_al_u1506_o,_al_u2408_o}),
    .q({\PWM8/FreCntr [21],\PWM8/FreCntr [15]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*~C)*~(D@B))"),
    //.LUTF1("(~(~D*B)*~(~C*A))"),
    //.LUTG0("(A*~(1*~C)*~(D@B))"),
    //.LUTG1("(~(~D*B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000100000100010),
    .INIT_LUTF1(16'b1111010100110001),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1111010100110001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg1_b23|PWM8/reg1_b12  (
    .a({\PWM8/FreCnt [22],_al_u2394_o}),
    .b({\PWM8/FreCnt [8],\PWM8/FreCnt [11]}),
    .c({\PWM8/FreCntr [23],\PWM8/FreCnt [22]}),
    .ce(\PWM8/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM8/FreCntr [9],\PWM8/FreCntr [12]}),
    .e({open_n13855,\PWM8/FreCntr [23]}),
    .mi({freq8[23],freq8[12]}),
    .f({_al_u2393_o,_al_u2395_o}),
    .q({\PWM8/FreCntr [23],\PWM8/FreCntr [12]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~B*~(0@C)*~(~D*A))"),
    //.LUTF1("(~(D*~B)*~(~C*A))"),
    //.LUTG0("(~B*~(1@C)*~(~D*A))"),
    //.LUTG1("(~(D*~B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001100000001),
    .INIT_LUTF1(16'b1100010011110101),
    .INIT_LUTG0(16'b0011000000010000),
    .INIT_LUTG1(16'b1100010011110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg1_b24|PWM8/reg1_b5  (
    .a({\PWM8/FreCnt [15],\PWM8/FreCnt [23]}),
    .b({\PWM8/FreCnt [23],\PWM8/FreCnt [26]}),
    .c({\PWM8/FreCntr [16],\PWM8/FreCnt [4]}),
    .ce(\PWM8/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM8/FreCntr [24],\PWM8/FreCntr [24]}),
    .e({open_n13872,\PWM8/FreCntr [5]}),
    .mi({freq8[24],freq8[5]}),
    .f({_al_u2409_o,_al_u2399_o}),
    .q({\PWM8/FreCntr [24],\PWM8/FreCntr [5]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*~C)*~(D*~B))"),
    //.LUTF1("(A*~(0*~C)*~(~D*B))"),
    //.LUTG0("(A*~(1*~C)*~(D*~B))"),
    //.LUTG1("(A*~(1*~C)*~(~D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000100010101010),
    .INIT_LUTF1(16'b1010101000100010),
    .INIT_LUTG0(16'b1000000010100000),
    .INIT_LUTG1(16'b1010000000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg1_b26|PWM8/reg1_b16  (
    .a({_al_u2403_o,_al_u2411_o}),
    .b({\PWM8/FreCnt [25],\PWM8/FreCnt [15]}),
    .c({\PWM8/FreCnt [3],\PWM8/FreCnt [25]}),
    .ce(\PWM8/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM8/FreCntr [26],\PWM8/FreCntr [16]}),
    .e({\PWM8/FreCntr [4],\PWM8/FreCntr [26]}),
    .mi({freq8[26],freq8[16]}),
    .f({_al_u2404_o,_al_u2412_o}),
    .q({\PWM8/FreCntr [26],\PWM8/FreCntr [16]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D@C)*~(0@B))"),
    //.LUTF1("(C*B*A*~(0@D))"),
    //.LUTG0("(A*~(D@C)*~(1@B))"),
    //.LUTG1("(C*B*A*~(1@D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010000000000010),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b1000000000001000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg1_b3|PWM8/reg1_b25  (
    .a({_al_u1499_o,_al_u2399_o}),
    .b({_al_u1501_o,\PWM8/FreCnt [2]}),
    .c({_al_u1502_o,\PWM8/FreCnt [24]}),
    .ce(\PWM8/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM8/FreCnt [3],\PWM8/FreCntr [25]}),
    .e({\PWM8/FreCntr [3],\PWM8/FreCntr [3]}),
    .mi({freq8[3],freq8[25]}),
    .f({_al_u1503_o,_al_u2400_o}),
    .q({\PWM8/FreCntr [3],\PWM8/FreCntr [25]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(~0*C)*~(~D*B))"),
    //.LUTF1("(A*~(0@C)*~(D@B))"),
    //.LUTG0("(A*~(~1*C)*~(~D*B))"),
    //.LUTG1("(A*~(1@C)*~(D@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101000000010),
    .INIT_LUTF1(16'b0000100000000010),
    .INIT_LUTG0(16'b1010101000100010),
    .INIT_LUTG1(16'b1000000000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg1_b4|PWM8/reg1_b22  (
    .a({_al_u1500_o,_al_u2405_o}),
    .b({\PWM8/FreCnt [4],\PWM8/FreCnt [21]}),
    .c({\PWM8/FreCnt [9],\PWM8/FreCnt [3]}),
    .ce(\PWM8/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM8/FreCntr [4],\PWM8/FreCntr [22]}),
    .e({\PWM8/FreCntr [9],\PWM8/FreCntr [4]}),
    .mi({freq8[4],freq8[22]}),
    .f({_al_u1501_o,_al_u2406_o}),
    .q({\PWM8/FreCntr [4],\PWM8/FreCntr [22]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*B*A*~(0@D))"),
    //.LUTF1("(~(~D*B)*~(C*~A))"),
    //.LUTG0("(C*B*A*~(1@D))"),
    //.LUTG1("(~(~D*B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b1010111100100011),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b1010111100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg1_b6|PWM8/reg1_b13  (
    .a({\PWM8/FreCnt [1],_al_u2395_o}),
    .b({\PWM8/FreCnt [5],_al_u2396_o}),
    .c({\PWM8/FreCntr [2],_al_u2397_o}),
    .ce(\PWM8/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM8/FreCntr [6],\PWM8/FreCnt [12]}),
    .e({open_n13937,\PWM8/FreCntr [13]}),
    .mi({freq8[6],freq8[13]}),
    .f({_al_u2396_o,_al_u2398_o}),
    .q({\PWM8/FreCntr [6],\PWM8/FreCntr [13]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(D*~B)*~(C*~A))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(~(D*~B)*~(C*~A))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000110010101111),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000110010101111),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg1_b7|PWM8/reg1_b8  (
    .a({\PWM8/FreCnt [6],\PWM8/FreCnt [7]}),
    .b({\PWM8/FreCnt [7],\PWM8/FreCnt [8]}),
    .c({\PWM8/FreCntr [6],\PWM8/FreCntr [8]}),
    .ce(\PWM8/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM8/FreCntr [7],\PWM8/FreCntr [9]}),
    .mi({freq8[7],freq8[8]}),
    .f({_al_u1500_o,_al_u2405_o}),
    .q({\PWM8/FreCntr [7],\PWM8/FreCntr [8]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg1_b9|PWM8/reg1_b0  (
    .b({_al_u1034_o,open_n13974}),
    .c({_al_u1036_o,\PWM8/n11 }),
    .ce(\PWM8/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({_al_u1032_o,\PWM8/n0_lutinv }),
    .mi({freq8[9],freq8[0]}),
    .f({\PWM8/n0_lutinv ,\PWM8/mux3_b0_sel_is_3_o }),
    .q({\PWM8/FreCntr [9],\PWM8/FreCntr [0]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg2_b0|PWM8/reg3_b0  (
    .a({\PWM8/pnumr [0],_al_u2391_o}),
    .b({pnum8[0],\PWM8/n24 }),
    .c({pnum8[32],pnumcnt8[0]}),
    .clk(clk100m),
    .d({pwm_start_stop[24],\PWM8/pnumr [0]}),
    .e({open_n13990,pwm_start_stop[24]}),
    .q({\PWM8/pnumr[0]_keep ,\PWM8/RemaTxNum[0]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011100010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg2_b10|PWM8/reg2_b9  (
    .a(\PWM8/pnumr [10:9]),
    .b({pnum8[10],pnum8[32]}),
    .c({pnum8[32],pnum8[9]}),
    .clk(clk100m),
    .d({pwm_start_stop[24],pwm_start_stop[24]}),
    .q({\PWM8/pnumr[10]_keep ,\PWM8/pnumr[9]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011100010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg2_b11|PWM8/reg2_b8  (
    .a({\PWM8/pnumr [11],\PWM8/pnumr [8]}),
    .b({pnum8[11],pnum8[32]}),
    .c({pnum8[32],pnum8[8]}),
    .clk(clk100m),
    .d({pwm_start_stop[24],pwm_start_stop[24]}),
    .q({\PWM8/pnumr[11]_keep ,\PWM8/pnumr[8]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg2_b12|PWM8/reg3_b12  (
    .a({\PWM8/pnumr [12],_al_u2383_o}),
    .b({pnum8[12],\PWM8/n24 }),
    .c({pnum8[32],pnumcnt8[12]}),
    .clk(clk100m),
    .d({pwm_start_stop[24],\PWM8/pnumr [12]}),
    .e({open_n14050,pwm_start_stop[24]}),
    .q({\PWM8/pnumr[12]_keep ,\PWM8/RemaTxNum[12]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg2_b13|PWM8/reg3_b13  (
    .a({\PWM8/pnumr [13],_al_u2381_o}),
    .b({pnum8[13],\PWM8/n24 }),
    .c({pnum8[32],pnumcnt8[13]}),
    .clk(clk100m),
    .d({pwm_start_stop[24],\PWM8/pnumr [13]}),
    .e({open_n14072,pwm_start_stop[24]}),
    .q({\PWM8/pnumr[13]_keep ,\PWM8/RemaTxNum[13]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011100010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011100010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg2_b14|PWM8/reg2_b5  (
    .a({\PWM8/pnumr [14],\PWM8/pnumr [5]}),
    .b({pnum8[14],pnum8[32]}),
    .c({pnum8[32],pnum8[5]}),
    .clk(clk100m),
    .d({pwm_start_stop[24],pwm_start_stop[24]}),
    .q({\PWM8/pnumr[14]_keep ,\PWM8/pnumr[5]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011100010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011100010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg2_b15|PWM8/reg2_b4  (
    .a({\PWM8/pnumr [15],\PWM8/pnumr [4]}),
    .b({pnum8[15],pnum8[32]}),
    .c({pnum8[32],pnum8[4]}),
    .clk(clk100m),
    .d({pwm_start_stop[24],pwm_start_stop[24]}),
    .q({\PWM8/pnumr[15]_keep ,\PWM8/pnumr[4]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg2_b16|PWM8/reg3_b16  (
    .a({\PWM8/pnumr [16],_al_u2375_o}),
    .b({pnum8[16],\PWM8/n24 }),
    .c({pnum8[32],pnumcnt8[16]}),
    .clk(clk100m),
    .d({pwm_start_stop[24],\PWM8/pnumr [16]}),
    .e({open_n14140,pwm_start_stop[24]}),
    .q({\PWM8/pnumr[16]_keep ,\PWM8/RemaTxNum[16]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg2_b17|PWM8/reg3_b17  (
    .a({\PWM8/pnumr [17],_al_u2373_o}),
    .b({pnum8[17],\PWM8/n24 }),
    .c({pnum8[32],pnumcnt8[17]}),
    .clk(clk100m),
    .d({pwm_start_stop[24],\PWM8/pnumr [17]}),
    .e({open_n14162,pwm_start_stop[24]}),
    .q({\PWM8/pnumr[17]_keep ,\PWM8/RemaTxNum[17]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg2_b18|PWM8/reg2_b22  (
    .a({\PWM8/pnumr [18],\PWM8/pnumr [22]}),
    .b({pnum8[18],pnum8[22]}),
    .c({pnum8[32],pnum8[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[24],pwm_start_stop[24]}),
    .q({\PWM8/pnumr[18]_keep ,\PWM8/pnumr[22]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg2_b19|PWM8/reg2_b21  (
    .a({\PWM8/pnumr [19],\PWM8/pnumr [21]}),
    .b({pnum8[19],pnum8[21]}),
    .c({pnum8[32],pnum8[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[24],pwm_start_stop[24]}),
    .q({\PWM8/pnumr[19]_keep ,\PWM8/pnumr[21]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg2_b1|PWM8/reg3_b1  (
    .a({\PWM8/pnumr [1],_al_u2389_o}),
    .b({pnum8[1],\PWM8/n24 }),
    .c({pnum8[32],pnumcnt8[1]}),
    .clk(clk100m),
    .d({pwm_start_stop[24],\PWM8/pnumr [1]}),
    .e({open_n14222,pwm_start_stop[24]}),
    .q({\PWM8/pnumr[1]_keep ,\PWM8/RemaTxNum[1]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg2_b20|PWM8/reg3_b20  (
    .a({\PWM8/pnumr [20],_al_u2365_o}),
    .b({pnum8[20],\PWM8/n24 }),
    .c({pnum8[32],pnumcnt8[20]}),
    .clk(clk100m),
    .d({pwm_start_stop[24],\PWM8/pnumr [20]}),
    .e({open_n14244,pwm_start_stop[24]}),
    .q({\PWM8/pnumr[20]_keep ,\PWM8/RemaTxNum[20]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg2_b23|PWM8/reg3_b23  (
    .a({\PWM8/pnumr [23],_al_u2359_o}),
    .b({pnum8[23],\PWM8/n24 }),
    .c({pnum8[32],pnumcnt8[23]}),
    .clk(clk100m),
    .d({pwm_start_stop[24],\PWM8/pnumr [23]}),
    .e({open_n14266,pwm_start_stop[24]}),
    .q({\PWM8/pnumr[23]_keep ,\PWM8/RemaTxNum[23]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg2_b24|PWM8/reg2_b31  (
    .a({\PWM8/pnumr [24],\PWM8/pnumr [31]}),
    .b({pnum8[24],pnum8[31]}),
    .c({pnum8[32],pnum8[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[24],pwm_start_stop[24]}),
    .q({\PWM8/pnumr[24]_keep ,\PWM8/pnumr[31]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg2_b25|PWM8/reg2_b30  (
    .a({\PWM8/pnumr [25],\PWM8/pnumr [30]}),
    .b({pnum8[25],pnum8[30]}),
    .c({pnum8[32],pnum8[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[24],pwm_start_stop[24]}),
    .q({\PWM8/pnumr[25]_keep ,\PWM8/pnumr[30]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg2_b26|PWM8/reg2_b29  (
    .a({\PWM8/pnumr [26],\PWM8/pnumr [29]}),
    .b({pnum8[26],pnum8[29]}),
    .c({pnum8[32],pnum8[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[24],pwm_start_stop[24]}),
    .q({\PWM8/pnumr[26]_keep ,\PWM8/pnumr[29]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg2_b27|PWM8/reg2_b28  (
    .a({\PWM8/pnumr [27],\PWM8/pnumr [28]}),
    .b({pnum8[27],pnum8[28]}),
    .c({pnum8[32],pnum8[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[24],pwm_start_stop[24]}),
    .q({\PWM8/pnumr[27]_keep ,\PWM8/pnumr[28]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg2_b2|PWM8/reg3_b2  (
    .a({\PWM8/pnumr [2],_al_u2367_o}),
    .b({pnum8[2],\PWM8/n24 }),
    .c({pnum8[32],pnumcnt8[2]}),
    .clk(clk100m),
    .d({pwm_start_stop[24],\PWM8/pnumr [2]}),
    .e({open_n14376,pwm_start_stop[24]}),
    .q({\PWM8/pnumr[2]_keep ,\PWM8/RemaTxNum[2]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg2_b3|PWM8/reg3_b3  (
    .a({\PWM8/pnumr [3],_al_u2357_o}),
    .b({pnum8[3],\PWM8/n24 }),
    .c({pnum8[32],pnumcnt8[3]}),
    .clk(clk100m),
    .d({pwm_start_stop[24],\PWM8/pnumr [3]}),
    .e({open_n14398,pwm_start_stop[24]}),
    .q({\PWM8/pnumr[3]_keep ,\PWM8/RemaTxNum[3]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg2_b6|PWM8/reg3_b6  (
    .a({\PWM8/pnumr [6],_al_u2351_o}),
    .b({pnum8[32],\PWM8/n24 }),
    .c({pnum8[6],pnumcnt8[6]}),
    .clk(clk100m),
    .d({pwm_start_stop[24],\PWM8/pnumr [6]}),
    .e({open_n14420,pwm_start_stop[24]}),
    .q({\PWM8/pnumr[6]_keep ,\PWM8/RemaTxNum[6]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg2_b7|PWM8/reg3_b7  (
    .a({\PWM8/pnumr [7],_al_u2349_o}),
    .b({pnum8[32],\PWM8/n24 }),
    .c({pnum8[7],pnumcnt8[7]}),
    .clk(clk100m),
    .d({pwm_start_stop[24],\PWM8/pnumr [7]}),
    .e({open_n14442,pwm_start_stop[24]}),
    .q({\PWM8/pnumr[7]_keep ,\PWM8/RemaTxNum[7]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg3_b10  (
    .a({_al_u2387_o,_al_u2387_o}),
    .b({\PWM8/n24 ,\PWM8/n24 }),
    .c({pnumcnt8[10],pnumcnt8[10]}),
    .clk(clk100m),
    .d({\PWM8/pnumr [10],\PWM8/pnumr [10]}),
    .mi({open_n14474,pwm_start_stop[24]}),
    .q({open_n14481,\PWM8/RemaTxNum[10]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg3_b11  (
    .a({_al_u2385_o,_al_u2385_o}),
    .b({\PWM8/n24 ,\PWM8/n24 }),
    .c({pnumcnt8[11],pnumcnt8[11]}),
    .clk(clk100m),
    .d({\PWM8/pnumr [11],\PWM8/pnumr [11]}),
    .mi({open_n14493,pwm_start_stop[24]}),
    .q({open_n14500,\PWM8/RemaTxNum[11]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg3_b14  (
    .a({_al_u2379_o,_al_u2379_o}),
    .b({\PWM8/n24 ,\PWM8/n24 }),
    .c({pnumcnt8[14],pnumcnt8[14]}),
    .clk(clk100m),
    .d({\PWM8/pnumr [14],\PWM8/pnumr [14]}),
    .mi({open_n14512,pwm_start_stop[24]}),
    .q({open_n14519,\PWM8/RemaTxNum[14]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg3_b15  (
    .a({_al_u2377_o,_al_u2377_o}),
    .b({\PWM8/n24 ,\PWM8/n24 }),
    .c({pnumcnt8[15],pnumcnt8[15]}),
    .clk(clk100m),
    .d({\PWM8/pnumr [15],\PWM8/pnumr [15]}),
    .mi({open_n14531,pwm_start_stop[24]}),
    .q({open_n14538,\PWM8/RemaTxNum[15]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg3_b18  (
    .a({_al_u2371_o,_al_u2371_o}),
    .b({\PWM8/n24 ,\PWM8/n24 }),
    .c({pnumcnt8[18],pnumcnt8[18]}),
    .clk(clk100m),
    .d({\PWM8/pnumr [18],\PWM8/pnumr [18]}),
    .mi({open_n14550,pwm_start_stop[24]}),
    .q({open_n14557,\PWM8/RemaTxNum[18]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg3_b19  (
    .a({_al_u2369_o,_al_u2369_o}),
    .b({\PWM8/n24 ,\PWM8/n24 }),
    .c({pnumcnt8[19],pnumcnt8[19]}),
    .clk(clk100m),
    .d({\PWM8/pnumr [19],\PWM8/pnumr [19]}),
    .mi({open_n14569,pwm_start_stop[24]}),
    .q({open_n14576,\PWM8/RemaTxNum[19]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg3_b21  (
    .a({_al_u2363_o,_al_u2363_o}),
    .b({\PWM8/n24 ,\PWM8/n24 }),
    .c({pnumcnt8[21],pnumcnt8[21]}),
    .clk(clk100m),
    .d({\PWM8/pnumr [21],\PWM8/pnumr [21]}),
    .mi({open_n14588,pwm_start_stop[24]}),
    .q({open_n14595,\PWM8/RemaTxNum[21]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg3_b22  (
    .a({_al_u2361_o,_al_u2361_o}),
    .b({\PWM8/n24 ,\PWM8/n24 }),
    .c({pnumcnt8[22],pnumcnt8[22]}),
    .clk(clk100m),
    .d({\PWM8/pnumr [22],\PWM8/pnumr [22]}),
    .mi({open_n14607,pwm_start_stop[24]}),
    .q({open_n14614,\PWM8/RemaTxNum[22]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg3_b4  (
    .a({_al_u2355_o,_al_u2355_o}),
    .b({\PWM8/n24 ,\PWM8/n24 }),
    .c({pnumcnt8[4],pnumcnt8[4]}),
    .clk(clk100m),
    .d({\PWM8/pnumr [4],\PWM8/pnumr [4]}),
    .mi({open_n14626,pwm_start_stop[24]}),
    .q({open_n14633,\PWM8/RemaTxNum[4]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg3_b5  (
    .a({_al_u2353_o,_al_u2353_o}),
    .b({\PWM8/n24 ,\PWM8/n24 }),
    .c({pnumcnt8[5],pnumcnt8[5]}),
    .clk(clk100m),
    .d({\PWM8/pnumr [5],\PWM8/pnumr [5]}),
    .mi({open_n14645,pwm_start_stop[24]}),
    .q({open_n14652,\PWM8/RemaTxNum[5]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg3_b8  (
    .a({_al_u2347_o,_al_u2347_o}),
    .b({\PWM8/n24 ,\PWM8/n24 }),
    .c({pnumcnt8[8],pnumcnt8[8]}),
    .clk(clk100m),
    .d({\PWM8/pnumr [8],\PWM8/pnumr [8]}),
    .mi({open_n14664,pwm_start_stop[24]}),
    .q({open_n14671,\PWM8/RemaTxNum[8]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/reg3_b9  (
    .a({_al_u2345_o,_al_u2345_o}),
    .b({\PWM8/n24 ,\PWM8/n24 }),
    .c({pnumcnt8[9],pnumcnt8[9]}),
    .clk(clk100m),
    .d({\PWM8/pnumr [9],\PWM8/pnumr [9]}),
    .mi({open_n14683,pwm_start_stop[24]}),
    .q({open_n14690,\PWM8/RemaTxNum[9]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_LSLICE #(
    //.MACRO("PWM8/sub0/ucin_al_u3419"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM8/sub0/u11_al_u3422  (
    .a({\PWM8/FreCnt [13],\PWM8/FreCnt [11]}),
    .b({\PWM8/FreCnt [14],\PWM8/FreCnt [12]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM8/sub0/c11 ),
    .f({\PWM8/n12 [13],\PWM8/n12 [11]}),
    .fco(\PWM8/sub0/c15 ),
    .fx({\PWM8/n12 [14],\PWM8/n12 [12]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM8/sub0/ucin_al_u3419"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM8/sub0/u15_al_u3423  (
    .a({\PWM8/FreCnt [17],\PWM8/FreCnt [15]}),
    .b({\PWM8/FreCnt [18],\PWM8/FreCnt [16]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM8/sub0/c15 ),
    .f({\PWM8/n12 [17],\PWM8/n12 [15]}),
    .fco(\PWM8/sub0/c19 ),
    .fx({\PWM8/n12 [18],\PWM8/n12 [16]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM8/sub0/ucin_al_u3419"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM8/sub0/u19_al_u3424  (
    .a({\PWM8/FreCnt [21],\PWM8/FreCnt [19]}),
    .b({\PWM8/FreCnt [22],\PWM8/FreCnt [20]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM8/sub0/c19 ),
    .f({\PWM8/n12 [21],\PWM8/n12 [19]}),
    .fco(\PWM8/sub0/c23 ),
    .fx({\PWM8/n12 [22],\PWM8/n12 [20]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM8/sub0/ucin_al_u3419"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM8/sub0/u23_al_u3425  (
    .a({\PWM8/FreCnt [25],\PWM8/FreCnt [23]}),
    .b({\PWM8/FreCnt [26],\PWM8/FreCnt [24]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM8/sub0/c23 ),
    .f({\PWM8/n12 [25],\PWM8/n12 [23]}),
    .fx({\PWM8/n12 [26],\PWM8/n12 [24]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM8/sub0/ucin_al_u3419"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM8/sub0/u3_al_u3420  (
    .a({\PWM8/FreCnt [5],\PWM8/FreCnt [3]}),
    .b({\PWM8/FreCnt [6],\PWM8/FreCnt [4]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM8/sub0/c3 ),
    .f({\PWM8/n12 [5],\PWM8/n12 [3]}),
    .fco(\PWM8/sub0/c7 ),
    .fx({\PWM8/n12 [6],\PWM8/n12 [4]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM8/sub0/ucin_al_u3419"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM8/sub0/u7_al_u3421  (
    .a({\PWM8/FreCnt [9],\PWM8/FreCnt [7]}),
    .b({\PWM8/FreCnt [10],\PWM8/FreCnt [8]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM8/sub0/c7 ),
    .f({\PWM8/n12 [9],\PWM8/n12 [7]}),
    .fco(\PWM8/sub0/c11 ),
    .fx({\PWM8/n12 [10],\PWM8/n12 [8]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM8/sub0/ucin_al_u3419"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'h0005),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM8/sub0/ucin_al_u3419  (
    .a({\PWM8/FreCnt [1],1'b0}),
    .b({\PWM8/FreCnt [2],\PWM8/FreCnt [0]}),
    .c(2'b11),
    .ce(\U_AHB/n20 ),
    .clk(clk100m),
    .d(2'b01),
    .e(2'b01),
    .mi({\U_AHB/h2h_hwdata [19],\U_AHB/h2h_hwdata [2]}),
    .f({\PWM8/n12 [1],open_n14813}),
    .fco(\PWM8/sub0/c3 ),
    .fx({\PWM8/n12 [2],\PWM8/n12 [0]}),
    .q({freq8[19],freq8[2]}));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM8/sub1/u0|PWM8/sub1/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("SUB_CARRY"),
    .INIT_LUT0(16'b0000000000000101),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM8/sub1/u0|PWM8/sub1/ucin  (
    .a({pnumcnt8[0],1'b0}),
    .b({1'b1,open_n14814}),
    .f({\PWM8/n26 [0],open_n14834}),
    .fco(\PWM8/sub1/c1 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM8/sub1/u0|PWM8/sub1/ucin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM8/sub1/u10|PWM8/sub1/u9  (
    .a(pnumcnt8[10:9]),
    .b(2'b00),
    .fci(\PWM8/sub1/c9 ),
    .f(\PWM8/n26 [10:9]),
    .fco(\PWM8/sub1/c11 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM8/sub1/u0|PWM8/sub1/ucin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM8/sub1/u12|PWM8/sub1/u11  (
    .a(pnumcnt8[12:11]),
    .b(2'b00),
    .fci(\PWM8/sub1/c11 ),
    .f(\PWM8/n26 [12:11]),
    .fco(\PWM8/sub1/c13 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM8/sub1/u0|PWM8/sub1/ucin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM8/sub1/u14|PWM8/sub1/u13  (
    .a(pnumcnt8[14:13]),
    .b(2'b00),
    .fci(\PWM8/sub1/c13 ),
    .f(\PWM8/n26 [14:13]),
    .fco(\PWM8/sub1/c15 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM8/sub1/u0|PWM8/sub1/ucin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM8/sub1/u16|PWM8/sub1/u15  (
    .a(pnumcnt8[16:15]),
    .b(2'b00),
    .fci(\PWM8/sub1/c15 ),
    .f(\PWM8/n26 [16:15]),
    .fco(\PWM8/sub1/c17 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM8/sub1/u0|PWM8/sub1/ucin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM8/sub1/u18|PWM8/sub1/u17  (
    .a(pnumcnt8[18:17]),
    .b(2'b00),
    .fci(\PWM8/sub1/c17 ),
    .f(\PWM8/n26 [18:17]),
    .fco(\PWM8/sub1/c19 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM8/sub1/u0|PWM8/sub1/ucin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM8/sub1/u20|PWM8/sub1/u19  (
    .a(pnumcnt8[20:19]),
    .b(2'b00),
    .fci(\PWM8/sub1/c19 ),
    .f(\PWM8/n26 [20:19]),
    .fco(\PWM8/sub1/c21 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM8/sub1/u0|PWM8/sub1/ucin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM8/sub1/u22|PWM8/sub1/u21  (
    .a(pnumcnt8[22:21]),
    .b(2'b00),
    .fci(\PWM8/sub1/c21 ),
    .f(\PWM8/n26 [22:21]),
    .fco(\PWM8/sub1/c23 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM8/sub1/u0|PWM8/sub1/ucin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM8/sub1/u23_al_u3476  (
    .a({open_n14993,pnumcnt8[23]}),
    .b({open_n14994,1'b0}),
    .fci(\PWM8/sub1/c23 ),
    .f({open_n15013,\PWM8/n26 [23]}));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM8/sub1/u0|PWM8/sub1/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM8/sub1/u2|PWM8/sub1/u1  (
    .a(pnumcnt8[2:1]),
    .b(2'b00),
    .fci(\PWM8/sub1/c1 ),
    .f(\PWM8/n26 [2:1]),
    .fco(\PWM8/sub1/c3 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM8/sub1/u0|PWM8/sub1/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM8/sub1/u4|PWM8/sub1/u3  (
    .a(pnumcnt8[4:3]),
    .b(2'b00),
    .fci(\PWM8/sub1/c3 ),
    .f(\PWM8/n26 [4:3]),
    .fco(\PWM8/sub1/c5 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM8/sub1/u0|PWM8/sub1/ucin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM8/sub1/u6|PWM8/sub1/u5  (
    .a(pnumcnt8[6:5]),
    .b(2'b00),
    .fci(\PWM8/sub1/c5 ),
    .f(\PWM8/n26 [6:5]),
    .fco(\PWM8/sub1/c7 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM8/sub1/u0|PWM8/sub1/ucin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM8/sub1/u8|PWM8/sub1/u7  (
    .a(pnumcnt8[8:7]),
    .b(2'b00),
    .fci(\PWM8/sub1/c7 ),
    .f(\PWM8/n26 [8:7]),
    .fco(\PWM8/sub1/c9 ));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[0]  (
    .i(\PWM9/RemaTxNum[0]_keep ),
    .o(pnumcnt9[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[10]  (
    .i(\PWM9/RemaTxNum[10]_keep ),
    .o(pnumcnt9[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[11]  (
    .i(\PWM9/RemaTxNum[11]_keep ),
    .o(pnumcnt9[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[12]  (
    .i(\PWM9/RemaTxNum[12]_keep ),
    .o(pnumcnt9[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[13]  (
    .i(\PWM9/RemaTxNum[13]_keep ),
    .o(pnumcnt9[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[14]  (
    .i(\PWM9/RemaTxNum[14]_keep ),
    .o(pnumcnt9[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[15]  (
    .i(\PWM9/RemaTxNum[15]_keep ),
    .o(pnumcnt9[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[16]  (
    .i(\PWM9/RemaTxNum[16]_keep ),
    .o(pnumcnt9[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[17]  (
    .i(\PWM9/RemaTxNum[17]_keep ),
    .o(pnumcnt9[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[18]  (
    .i(\PWM9/RemaTxNum[18]_keep ),
    .o(pnumcnt9[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[19]  (
    .i(\PWM9/RemaTxNum[19]_keep ),
    .o(pnumcnt9[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[1]  (
    .i(\PWM9/RemaTxNum[1]_keep ),
    .o(pnumcnt9[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[20]  (
    .i(\PWM9/RemaTxNum[20]_keep ),
    .o(pnumcnt9[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[21]  (
    .i(\PWM9/RemaTxNum[21]_keep ),
    .o(pnumcnt9[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[22]  (
    .i(\PWM9/RemaTxNum[22]_keep ),
    .o(pnumcnt9[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[23]  (
    .i(\PWM9/RemaTxNum[23]_keep ),
    .o(pnumcnt9[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[2]  (
    .i(\PWM9/RemaTxNum[2]_keep ),
    .o(pnumcnt9[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[3]  (
    .i(\PWM9/RemaTxNum[3]_keep ),
    .o(pnumcnt9[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[4]  (
    .i(\PWM9/RemaTxNum[4]_keep ),
    .o(pnumcnt9[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[5]  (
    .i(\PWM9/RemaTxNum[5]_keep ),
    .o(pnumcnt9[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[6]  (
    .i(\PWM9/RemaTxNum[6]_keep ),
    .o(pnumcnt9[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[7]  (
    .i(\PWM9/RemaTxNum[7]_keep ),
    .o(pnumcnt9[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[8]  (
    .i(\PWM9/RemaTxNum[8]_keep ),
    .o(pnumcnt9[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[9]  (
    .i(\PWM9/RemaTxNum[9]_keep ),
    .o(pnumcnt9[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_dir  (
    .i(\PWM9/dir_keep ),
    .o(dir_pad[9]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[0]  (
    .i(\PWM9/pnumr[0]_keep ),
    .o(\PWM9/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[10]  (
    .i(\PWM9/pnumr[10]_keep ),
    .o(\PWM9/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[11]  (
    .i(\PWM9/pnumr[11]_keep ),
    .o(\PWM9/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[12]  (
    .i(\PWM9/pnumr[12]_keep ),
    .o(\PWM9/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[13]  (
    .i(\PWM9/pnumr[13]_keep ),
    .o(\PWM9/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[14]  (
    .i(\PWM9/pnumr[14]_keep ),
    .o(\PWM9/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[15]  (
    .i(\PWM9/pnumr[15]_keep ),
    .o(\PWM9/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[16]  (
    .i(\PWM9/pnumr[16]_keep ),
    .o(\PWM9/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[17]  (
    .i(\PWM9/pnumr[17]_keep ),
    .o(\PWM9/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[18]  (
    .i(\PWM9/pnumr[18]_keep ),
    .o(\PWM9/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[19]  (
    .i(\PWM9/pnumr[19]_keep ),
    .o(\PWM9/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[1]  (
    .i(\PWM9/pnumr[1]_keep ),
    .o(\PWM9/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[20]  (
    .i(\PWM9/pnumr[20]_keep ),
    .o(\PWM9/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[21]  (
    .i(\PWM9/pnumr[21]_keep ),
    .o(\PWM9/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[22]  (
    .i(\PWM9/pnumr[22]_keep ),
    .o(\PWM9/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[23]  (
    .i(\PWM9/pnumr[23]_keep ),
    .o(\PWM9/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[24]  (
    .i(\PWM9/pnumr[24]_keep ),
    .o(\PWM9/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[25]  (
    .i(\PWM9/pnumr[25]_keep ),
    .o(\PWM9/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[26]  (
    .i(\PWM9/pnumr[26]_keep ),
    .o(\PWM9/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[27]  (
    .i(\PWM9/pnumr[27]_keep ),
    .o(\PWM9/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[28]  (
    .i(\PWM9/pnumr[28]_keep ),
    .o(\PWM9/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[29]  (
    .i(\PWM9/pnumr[29]_keep ),
    .o(\PWM9/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[2]  (
    .i(\PWM9/pnumr[2]_keep ),
    .o(\PWM9/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[30]  (
    .i(\PWM9/pnumr[30]_keep ),
    .o(\PWM9/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[31]  (
    .i(\PWM9/pnumr[31]_keep ),
    .o(\PWM9/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[3]  (
    .i(\PWM9/pnumr[3]_keep ),
    .o(\PWM9/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[4]  (
    .i(\PWM9/pnumr[4]_keep ),
    .o(\PWM9/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[5]  (
    .i(\PWM9/pnumr[5]_keep ),
    .o(\PWM9/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[6]  (
    .i(\PWM9/pnumr[6]_keep ),
    .o(\PWM9/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[7]  (
    .i(\PWM9/pnumr[7]_keep ),
    .o(\PWM9/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[8]  (
    .i(\PWM9/pnumr[8]_keep ),
    .o(\PWM9/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[9]  (
    .i(\PWM9/pnumr[9]_keep ),
    .o(\PWM9/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pwm  (
    .i(\PWM9/pwm_keep ),
    .o(pwm_pad[9]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_stopreq  (
    .i(\PWM9/stopreq_keep ),
    .o(\PWM9/stopreq ));  // src/OnePWM.v(14)
  EF2_PHY_MSLICE #(
    //.LUT0("(D*~(C)*~((~0*~(B*A)))+D*C*~((~0*~(B*A)))+~(D)*C*(~0*~(B*A))+D*C*(~0*~(B*A)))"),
    //.LUT1("(D*~(C)*~((~1*~(B*A)))+D*C*~((~1*~(B*A)))+~(D)*C*(~1*~(B*A))+D*C*(~1*~(B*A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111100001110000),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/dir_reg  (
    .a({\PWM9/n24 ,\PWM9/n24 }),
    .b({\PWM9/n25_neg_lutinv ,\PWM9/n25_neg_lutinv }),
    .c({dir_pad[9],dir_pad[9]}),
    .clk(clk100m),
    .d({\PWM9/pnumr [31],\PWM9/pnumr [31]}),
    .mi({open_n15118,pwm_start_stop[25]}),
    .q({open_n15125,\PWM9/dir_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("~(~0*~(D*C*B*A))"),
    //.LUT1("~(~1*~(D*C*B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b1111111111111111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM9/pwm_reg  (
    .a({_al_u1521_o,_al_u1521_o}),
    .b({_al_u1527_o,_al_u1527_o}),
    .c({_al_u1529_o,_al_u1529_o}),
    .clk(clk100m),
    .d({_al_u1531_o,_al_u1531_o}),
    .mi({open_n15137,pwm_pad[9]}),
    .sr(\PWM9/u14_sel_is_1_o ),
    .q({open_n15143,\PWM9/pwm_keep }));  // src/OnePWM.v(45)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM9/reg0_b0|PWM9/reg0_b8  (
    .b({\PWM9/n12 [0],\PWM9/n12 [8]}),
    .c({freq9[0],freq9[8]}),
    .clk(clk100m),
    .d({\PWM9/n0_lutinv ,\PWM9/n0_lutinv }),
    .sr(\PWM9/n11 ),
    .q({\PWM9/FreCnt [0],\PWM9/FreCnt [8]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM9/reg0_b10|PWM9/reg0_b7  (
    .b({\PWM9/n12 [10],\PWM9/n12 [7]}),
    .c({freq9[10],freq9[7]}),
    .clk(clk100m),
    .d({\PWM9/n0_lutinv ,\PWM9/n0_lutinv }),
    .sr(\PWM9/n11 ),
    .q({\PWM9/FreCnt [10],\PWM9/FreCnt [7]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM9/reg0_b11|PWM9/reg0_b18  (
    .b({\PWM9/n12 [11],\PWM9/n12 [18]}),
    .c({freq9[11],freq9[18]}),
    .clk(clk100m),
    .d({\PWM9/n0_lutinv ,\PWM9/n0_lutinv }),
    .sr(\PWM9/n11 ),
    .q({\PWM9/FreCnt [11],\PWM9/FreCnt [18]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM9/reg0_b14|PWM9/reg0_b9  (
    .b({\PWM9/n12 [14],\PWM9/n12 [9]}),
    .c({freq9[14],freq9[9]}),
    .clk(clk100m),
    .d({\PWM9/n0_lutinv ,\PWM9/n0_lutinv }),
    .sr(\PWM9/n11 ),
    .q({\PWM9/FreCnt [14],\PWM9/FreCnt [9]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM9/reg0_b16|PWM9/reg0_b26  (
    .b({\PWM9/n12 [16],\PWM9/n12 [26]}),
    .c({freq9[16],freq9[26]}),
    .clk(clk100m),
    .d({\PWM9/n0_lutinv ,\PWM9/n0_lutinv }),
    .sr(\PWM9/n11 ),
    .q({\PWM9/FreCnt [16],\PWM9/FreCnt [26]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM9/reg0_b20|PWM9/reg0_b25  (
    .b({\PWM9/n12 [20],\PWM9/n12 [25]}),
    .c({freq9[20],freq9[25]}),
    .clk(clk100m),
    .d({\PWM9/n0_lutinv ,\PWM9/n0_lutinv }),
    .sr(\PWM9/n11 ),
    .q({\PWM9/FreCnt [20],\PWM9/FreCnt [25]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWM9/reg0_b22|PWM9/reg0_b24  (
    .b({\PWM9/n12 [22],\PWM9/n12 [24]}),
    .c({freq9[22],freq9[24]}),
    .clk(clk100m),
    .d({\PWM9/n0_lutinv ,\PWM9/n0_lutinv }),
    .sr(\PWM9/n11 ),
    .q({\PWM9/FreCnt [22],\PWM9/FreCnt [24]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(~0*C)*~(D@B))"),
    //.LUTF1("(C*B*A*~(0@D))"),
    //.LUTG0("(A*~(~1*C)*~(D@B))"),
    //.LUTG1("(C*B*A*~(1@D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b1000100000100010),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg1_b10|PWM9/reg1_b15  (
    .a({_al_u2475_o,_al_u2474_o}),
    .b({_al_u2477_o,\PWM9/FreCnt [14]}),
    .c({_al_u2478_o,\PWM9/FreCnt [8]}),
    .ce(\PWM9/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM9/FreCnt [9],\PWM9/FreCntr [15]}),
    .e(\PWM9/FreCntr [10:9]),
    .mi({freq9[10],freq9[15]}),
    .f({_al_u2479_o,_al_u2475_o}),
    .q({\PWM9/FreCntr [10],\PWM9/FreCntr [15]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~D*B)*~(~C*A))"),
    //.LUT1("(C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111010100110001),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg1_b11|PWM9/reg1_b4  (
    .a({open_n15308,\PWM9/FreCnt [10]}),
    .b({open_n15309,\PWM9/FreCnt [3]}),
    .c({\PWM9/FreCntr [11],\PWM9/FreCntr [11]}),
    .ce(\PWM9/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM9/FreCnt [10],\PWM9/FreCntr [4]}),
    .mi({freq9[11],freq9[4]}),
    .f({_al_u2484_o,_al_u2473_o}),
    .q({\PWM9/FreCntr [11],\PWM9/FreCntr [4]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(D*~B)*~(~C*A))"),
    //.LUTF1("(~(~D*B)*~(~C*A))"),
    //.LUTG0("(~(D*~B)*~(~C*A))"),
    //.LUTG1("(~(~D*B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100010011110101),
    .INIT_LUTF1(16'b1111010100110001),
    .INIT_LUTG0(16'b1100010011110101),
    .INIT_LUTG1(16'b1111010100110001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg1_b14|PWM9/reg1_b2  (
    .a({\PWM9/FreCnt [13],\PWM9/FreCnt [1]}),
    .b({\PWM9/FreCnt [7],\PWM9/FreCnt [23]}),
    .c({\PWM9/FreCntr [14],\PWM9/FreCntr [2]}),
    .ce(\PWM9/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM9/FreCntr [8],\PWM9/FreCntr [24]}),
    .mi({freq9[14],freq9[2]}),
    .f({_al_u2482_o,_al_u2480_o}),
    .q({\PWM9/FreCntr [14],\PWM9/FreCntr [2]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~A*~(0@C)*~(~D*B))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(~A*~(1@C)*~(~D*B))"),
    //.LUTG1("(C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010100000001),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0101000000010000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg1_b16|PWM9/reg1_b21  (
    .a({open_n15342,_al_u2486_o}),
    .b({open_n15343,\PWM9/FreCnt [15]}),
    .c({\PWM9/FreCntr [16],\PWM9/FreCnt [20]}),
    .ce(\PWM9/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM9/FreCnt [15],\PWM9/FreCntr [16]}),
    .e({open_n15344,\PWM9/FreCntr [21]}),
    .mi({freq9[16],freq9[21]}),
    .f({_al_u2495_o,_al_u2487_o}),
    .q({\PWM9/FreCntr [16],\PWM9/FreCntr [21]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(D@B)*~(C@A))"),
    //.LUT1("(D*~(C@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000010000100001),
    .INIT_LUT1(16'b1100001100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg1_b17|PWM9/reg1_b26  (
    .a({open_n15361,\PWM9/FreCnt [20]}),
    .b({\PWM9/FreCnt [16],\PWM9/FreCnt [26]}),
    .c({\PWM9/FreCntr [17],\PWM9/FreCntr [20]}),
    .ce(\PWM9/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({_al_u2476_o,\PWM9/FreCntr [26]}),
    .mi({freq9[17],freq9[26]}),
    .f({_al_u2477_o,_al_u1520_o}),
    .q({\PWM9/FreCntr [17],\PWM9/FreCntr [26]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(~0*C)*~(D*~B))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(A*~(~1*C)*~(D*~B))"),
    //.LUTG1("(~C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000001010),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b1000100010101010),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg1_b19|PWM9/reg1_b24  (
    .a({open_n15376,_al_u2482_o}),
    .b({open_n15377,\PWM9/FreCnt [18]}),
    .c({\PWM9/FreCntr [19],\PWM9/FreCnt [23]}),
    .ce(\PWM9/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM9/FreCnt [18],\PWM9/FreCntr [19]}),
    .e({open_n15378,\PWM9/FreCntr [24]}),
    .mi({freq9[19],freq9[24]}),
    .f({_al_u2486_o,_al_u2483_o}),
    .q({\PWM9/FreCntr [19],\PWM9/FreCntr [24]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~D*B)*~(~C*A))"),
    //.LUT1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111010100110001),
    .INIT_LUT1(16'b1000010000100001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg1_b1|PWM9/reg1_b12  (
    .a({\PWM9/FreCnt [0],\PWM9/FreCnt [12]}),
    .b({\PWM9/FreCnt [11],\PWM9/FreCnt [15]}),
    .c({\PWM9/FreCntr [1],\PWM9/FreCntr [12]}),
    .ce(\PWM9/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM9/FreCntr [12],\PWM9/FreCntr [15]}),
    .mi({freq9[1],freq9[12]}),
    .f({_al_u2491_o,_al_u1526_o}),
    .q({\PWM9/FreCntr [1],\PWM9/FreCntr [12]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~B*~(0@C)*~(D*~A))"),
    //.LUTF1("(~A*~(0@C)*~(~D*B))"),
    //.LUTG0("(~B*~(1@C)*~(D*~A))"),
    //.LUTG1("(~A*~(1@C)*~(~D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000000011),
    .INIT_LUTF1(16'b0000010100000001),
    .INIT_LUTG0(16'b0010000000110000),
    .INIT_LUTG1(16'b0101000000010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg1_b20|PWM9/reg1_b5  (
    .a({_al_u2495_o,\PWM9/FreCnt [19]}),
    .b({\PWM9/FreCnt [19],\PWM9/FreCnt [26]}),
    .c({\PWM9/FreCnt [25],\PWM9/FreCnt [4]}),
    .ce(\PWM9/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM9/FreCntr [20],\PWM9/FreCntr [20]}),
    .e({\PWM9/FreCntr [26],\PWM9/FreCntr [5]}),
    .mi({freq9[20],freq9[5]}),
    .f({_al_u2496_o,_al_u2489_o}),
    .q({\PWM9/FreCntr [20],\PWM9/FreCntr [5]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(~0*C)*~(~D*B))"),
    //.LUTF1("(~(D*~B)*~(C*~A))"),
    //.LUTG0("(A*~(~1*C)*~(~D*B))"),
    //.LUTG1("(~(D*~B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101000000010),
    .INIT_LUTF1(16'b1000110010101111),
    .INIT_LUTG0(16'b1010101000100010),
    .INIT_LUTG1(16'b1000110010101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg1_b22|PWM9/reg1_b18  (
    .a({\PWM9/FreCnt [12],_al_u2493_o}),
    .b({\PWM9/FreCnt [21],\PWM9/FreCnt [17]}),
    .c({\PWM9/FreCntr [13],\PWM9/FreCnt [21]}),
    .ce(\PWM9/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM9/FreCntr [22],\PWM9/FreCntr [18]}),
    .e({open_n15425,\PWM9/FreCntr [22]}),
    .mi({freq9[22],freq9[18]}),
    .f({_al_u2476_o,_al_u2494_o}),
    .q({\PWM9/FreCntr [22],\PWM9/FreCntr [18]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*~C)*~(~D*B))"),
    //.LUTF1("(A*~(~0*C)*~(D*~B))"),
    //.LUTG0("(A*~(1*~C)*~(~D*B))"),
    //.LUTG1("(A*~(~1*C)*~(D*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101000100010),
    .INIT_LUTF1(16'b0000100000001010),
    .INIT_LUTG0(16'b1010000000100000),
    .INIT_LUTG1(16'b1000100010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg1_b6|PWM9/reg1_b13  (
    .a({_al_u2473_o,_al_u2480_o}),
    .b({\PWM9/FreCnt [1],\PWM9/FreCnt [12]}),
    .c({\PWM9/FreCnt [5],\PWM9/FreCnt [5]}),
    .ce(\PWM9/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM9/FreCntr [2],\PWM9/FreCntr [13]}),
    .e({\PWM9/FreCntr [6],\PWM9/FreCntr [6]}),
    .mi({freq9[6],freq9[13]}),
    .f({_al_u2474_o,_al_u2481_o}),
    .q({\PWM9/FreCntr [6],\PWM9/FreCntr [13]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg1_b7|PWM9/reg1_b25  (
    .a({\PWM9/FreCnt [7],_al_u2489_o}),
    .b({\PWM9/FreCnt [9],\PWM9/FreCnt [24]}),
    .c({\PWM9/FreCntr [7],\PWM9/FreCnt [6]}),
    .ce(\PWM9/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM9/FreCntr [9],\PWM9/FreCntr [25]}),
    .e({open_n15458,\PWM9/FreCntr [7]}),
    .mi({freq9[7],freq9[25]}),
    .f({_al_u1528_o,_al_u2490_o}),
    .q({\PWM9/FreCntr [7],\PWM9/FreCntr [25]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(~(D*~B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b1000110010101111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg1_b8|PWM9/reg1_b9  (
    .a({\PWM9/FreCnt [7],open_n15475}),
    .b({\PWM9/FreCnt [8],_al_u1071_o}),
    .c({\PWM9/FreCntr [8],_al_u1073_o}),
    .ce(\PWM9/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM9/FreCntr [9],_al_u1069_o}),
    .mi({freq9[8],freq9[9]}),
    .f({_al_u2493_o,\PWM9/n0_lutinv }),
    .q({\PWM9/FreCntr [8],\PWM9/FreCntr [9]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011100010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011100010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg2_b0|PWM9/reg2_b9  (
    .a({\PWM9/pnumr [0],\PWM9/pnumr [9]}),
    .b({pnum9[0],pnum9[32]}),
    .c({pnum9[32],pnum9[9]}),
    .clk(clk100m),
    .d({pwm_start_stop[25],pwm_start_stop[25]}),
    .q({\PWM9/pnumr[0]_keep ,\PWM9/pnumr[9]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg2_b10|PWM9/reg3_b10  (
    .a({\PWM9/pnumr [10],_al_u2467_o}),
    .b({pnum9[10],\PWM9/n24 }),
    .c({pnum9[32],pnumcnt9[10]}),
    .clk(clk100m),
    .d({pwm_start_stop[25],\PWM9/pnumr [10]}),
    .e({open_n15514,pwm_start_stop[25]}),
    .q({\PWM9/pnumr[10]_keep ,\PWM9/RemaTxNum[10]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011100010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011100010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg2_b11|PWM9/reg2_b6  (
    .a({\PWM9/pnumr [11],\PWM9/pnumr [6]}),
    .b({pnum9[11],pnum9[32]}),
    .c({pnum9[32],pnum9[6]}),
    .clk(clk100m),
    .d({pwm_start_stop[25],pwm_start_stop[25]}),
    .q({\PWM9/pnumr[11]_keep ,\PWM9/pnumr[6]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011100010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg2_b12|PWM9/reg2_b5  (
    .a({\PWM9/pnumr [12],\PWM9/pnumr [5]}),
    .b({pnum9[12],pnum9[32]}),
    .c({pnum9[32],pnum9[5]}),
    .clk(clk100m),
    .d({pwm_start_stop[25],pwm_start_stop[25]}),
    .q({\PWM9/pnumr[12]_keep ,\PWM9/pnumr[5]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg2_b13|PWM9/reg3_b13  (
    .a({\PWM9/pnumr [13],_al_u2461_o}),
    .b({pnum9[13],\PWM9/n24 }),
    .c({pnum9[32],pnumcnt9[13]}),
    .clk(clk100m),
    .d({pwm_start_stop[25],\PWM9/pnumr [13]}),
    .e({open_n15578,pwm_start_stop[25]}),
    .q({\PWM9/pnumr[13]_keep ,\PWM9/RemaTxNum[13]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg2_b14|PWM9/reg3_b14  (
    .a({\PWM9/pnumr [14],_al_u2459_o}),
    .b({pnum9[14],\PWM9/n24 }),
    .c({pnum9[32],pnumcnt9[14]}),
    .clk(clk100m),
    .d({pwm_start_stop[25],\PWM9/pnumr [14]}),
    .e({open_n15600,pwm_start_stop[25]}),
    .q({\PWM9/pnumr[14]_keep ,\PWM9/RemaTxNum[14]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg2_b15|PWM9/reg2_b23  (
    .a({\PWM9/pnumr [15],\PWM9/pnumr [23]}),
    .b({pnum9[15],pnum9[23]}),
    .c({pnum9[32],pnum9[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[25],pwm_start_stop[25]}),
    .q({\PWM9/pnumr[15]_keep ,\PWM9/pnumr[23]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg2_b16|PWM9/reg2_b22  (
    .a({\PWM9/pnumr [16],\PWM9/pnumr [22]}),
    .b({pnum9[16],pnum9[22]}),
    .c({pnum9[32],pnum9[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[25],pwm_start_stop[25]}),
    .q({\PWM9/pnumr[16]_keep ,\PWM9/pnumr[22]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg2_b17|PWM9/reg3_b17  (
    .a({\PWM9/pnumr [17],_al_u2453_o}),
    .b({pnum9[17],\PWM9/n24 }),
    .c({pnum9[32],pnumcnt9[17]}),
    .clk(clk100m),
    .d({pwm_start_stop[25],\PWM9/pnumr [17]}),
    .e({open_n15664,pwm_start_stop[25]}),
    .q({\PWM9/pnumr[17]_keep ,\PWM9/RemaTxNum[17]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg2_b18|PWM9/reg3_b18  (
    .a({\PWM9/pnumr [18],_al_u2451_o}),
    .b({pnum9[18],\PWM9/n24 }),
    .c({pnum9[32],pnumcnt9[18]}),
    .clk(clk100m),
    .d({pwm_start_stop[25],\PWM9/pnumr [18]}),
    .e({open_n15686,pwm_start_stop[25]}),
    .q({\PWM9/pnumr[18]_keep ,\PWM9/RemaTxNum[18]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg2_b19|PWM9/reg2_b2  (
    .a({\PWM9/pnumr [19],\PWM9/pnumr [2]}),
    .b({pnum9[19],pnum9[2]}),
    .c({pnum9[32],pnum9[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[25],pwm_start_stop[25]}),
    .q({\PWM9/pnumr[19]_keep ,\PWM9/pnumr[2]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg2_b1|PWM9/reg3_b1  (
    .a({\PWM9/pnumr [1],_al_u2469_o}),
    .b({pnum9[1],\PWM9/n24 }),
    .c({pnum9[32],pnumcnt9[1]}),
    .clk(clk100m),
    .d({pwm_start_stop[25],\PWM9/pnumr [1]}),
    .e({open_n15731,pwm_start_stop[25]}),
    .q({\PWM9/pnumr[1]_keep ,\PWM9/RemaTxNum[1]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg2_b20|PWM9/reg3_b20  (
    .a({\PWM9/pnumr [20],_al_u2445_o}),
    .b({pnum9[20],\PWM9/n24 }),
    .c({pnum9[32],pnumcnt9[20]}),
    .clk(clk100m),
    .d({pwm_start_stop[25],\PWM9/pnumr [20]}),
    .e({open_n15753,pwm_start_stop[25]}),
    .q({\PWM9/pnumr[20]_keep ,\PWM9/RemaTxNum[20]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg2_b21|PWM9/reg3_b21  (
    .a({\PWM9/pnumr [21],_al_u2443_o}),
    .b({pnum9[21],\PWM9/n24 }),
    .c({pnum9[32],pnumcnt9[21]}),
    .clk(clk100m),
    .d({pwm_start_stop[25],\PWM9/pnumr [21]}),
    .e({open_n15775,pwm_start_stop[25]}),
    .q({\PWM9/pnumr[21]_keep ,\PWM9/RemaTxNum[21]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg2_b24|PWM9/reg2_b31  (
    .a({\PWM9/pnumr [24],\PWM9/pnumr [31]}),
    .b({pnum9[24],pnum9[31]}),
    .c({pnum9[32],pnum9[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[25],pwm_start_stop[25]}),
    .q({\PWM9/pnumr[24]_keep ,\PWM9/pnumr[31]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg2_b25|PWM9/reg2_b30  (
    .a({\PWM9/pnumr [25],\PWM9/pnumr [30]}),
    .b({pnum9[25],pnum9[30]}),
    .c({pnum9[32],pnum9[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[25],pwm_start_stop[25]}),
    .q({\PWM9/pnumr[25]_keep ,\PWM9/pnumr[30]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg2_b26|PWM9/reg2_b29  (
    .a({\PWM9/pnumr [26],\PWM9/pnumr [29]}),
    .b({pnum9[26],pnum9[29]}),
    .c({pnum9[32],pnum9[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[25],pwm_start_stop[25]}),
    .q({\PWM9/pnumr[26]_keep ,\PWM9/pnumr[29]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg2_b27|PWM9/reg2_b28  (
    .a({\PWM9/pnumr [27],\PWM9/pnumr [28]}),
    .b({pnum9[27],pnum9[28]}),
    .c({pnum9[32],pnum9[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[25],pwm_start_stop[25]}),
    .q({\PWM9/pnumr[27]_keep ,\PWM9/pnumr[28]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg2_b3|PWM9/reg3_b3  (
    .a({\PWM9/pnumr [3],_al_u2437_o}),
    .b({pnum9[3],\PWM9/n24 }),
    .c({pnum9[32],pnumcnt9[3]}),
    .clk(clk100m),
    .d({pwm_start_stop[25],\PWM9/pnumr [3]}),
    .e({open_n15885,pwm_start_stop[25]}),
    .q({\PWM9/pnumr[3]_keep ,\PWM9/RemaTxNum[3]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg2_b4|PWM9/reg3_b4  (
    .a({\PWM9/pnumr [4],_al_u2435_o}),
    .b({pnum9[32],\PWM9/n24 }),
    .c({pnum9[4],pnumcnt9[4]}),
    .clk(clk100m),
    .d({pwm_start_stop[25],\PWM9/pnumr [4]}),
    .e({open_n15907,pwm_start_stop[25]}),
    .q({\PWM9/pnumr[4]_keep ,\PWM9/RemaTxNum[4]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg2_b7|PWM9/reg3_b7  (
    .a({\PWM9/pnumr [7],_al_u2429_o}),
    .b({pnum9[32],\PWM9/n24 }),
    .c({pnum9[7],pnumcnt9[7]}),
    .clk(clk100m),
    .d({pwm_start_stop[25],\PWM9/pnumr [7]}),
    .e({open_n15929,pwm_start_stop[25]}),
    .q({\PWM9/pnumr[7]_keep ,\PWM9/RemaTxNum[7]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg2_b8|PWM9/reg3_b8  (
    .a({\PWM9/pnumr [8],_al_u2427_o}),
    .b({pnum9[32],\PWM9/n24 }),
    .c({pnum9[8],pnumcnt9[8]}),
    .clk(clk100m),
    .d({pwm_start_stop[25],\PWM9/pnumr [8]}),
    .e({open_n15951,pwm_start_stop[25]}),
    .q({\PWM9/pnumr[8]_keep ,\PWM9/RemaTxNum[8]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg3_b0  (
    .a({_al_u2471_o,_al_u2471_o}),
    .b({\PWM9/n24 ,\PWM9/n24 }),
    .c({pnumcnt9[0],pnumcnt9[0]}),
    .clk(clk100m),
    .d({\PWM9/pnumr [0],\PWM9/pnumr [0]}),
    .mi({open_n15983,pwm_start_stop[25]}),
    .q({open_n15990,\PWM9/RemaTxNum[0]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg3_b11  (
    .a({_al_u2465_o,_al_u2465_o}),
    .b({\PWM9/n24 ,\PWM9/n24 }),
    .c({pnumcnt9[11],pnumcnt9[11]}),
    .clk(clk100m),
    .d({\PWM9/pnumr [11],\PWM9/pnumr [11]}),
    .mi({open_n16002,pwm_start_stop[25]}),
    .q({open_n16009,\PWM9/RemaTxNum[11]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg3_b12  (
    .a({_al_u2463_o,_al_u2463_o}),
    .b({\PWM9/n24 ,\PWM9/n24 }),
    .c({pnumcnt9[12],pnumcnt9[12]}),
    .clk(clk100m),
    .d({\PWM9/pnumr [12],\PWM9/pnumr [12]}),
    .mi({open_n16021,pwm_start_stop[25]}),
    .q({open_n16028,\PWM9/RemaTxNum[12]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg3_b15  (
    .a({_al_u2457_o,_al_u2457_o}),
    .b({\PWM9/n24 ,\PWM9/n24 }),
    .c({pnumcnt9[15],pnumcnt9[15]}),
    .clk(clk100m),
    .d({\PWM9/pnumr [15],\PWM9/pnumr [15]}),
    .mi({open_n16040,pwm_start_stop[25]}),
    .q({open_n16047,\PWM9/RemaTxNum[15]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg3_b16  (
    .a({_al_u2455_o,_al_u2455_o}),
    .b({\PWM9/n24 ,\PWM9/n24 }),
    .c({pnumcnt9[16],pnumcnt9[16]}),
    .clk(clk100m),
    .d({\PWM9/pnumr [16],\PWM9/pnumr [16]}),
    .mi({open_n16059,pwm_start_stop[25]}),
    .q({open_n16066,\PWM9/RemaTxNum[16]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg3_b19  (
    .a({_al_u2449_o,_al_u2449_o}),
    .b({\PWM9/n24 ,\PWM9/n24 }),
    .c({pnumcnt9[19],pnumcnt9[19]}),
    .clk(clk100m),
    .d({\PWM9/pnumr [19],\PWM9/pnumr [19]}),
    .mi({open_n16078,pwm_start_stop[25]}),
    .q({open_n16085,\PWM9/RemaTxNum[19]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg3_b2  (
    .a({_al_u2447_o,_al_u2447_o}),
    .b({\PWM9/n24 ,\PWM9/n24 }),
    .c({pnumcnt9[2],pnumcnt9[2]}),
    .clk(clk100m),
    .d({\PWM9/pnumr [2],\PWM9/pnumr [2]}),
    .mi({open_n16097,pwm_start_stop[25]}),
    .q({open_n16104,\PWM9/RemaTxNum[2]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg3_b22  (
    .a({_al_u2441_o,_al_u2441_o}),
    .b({\PWM9/n24 ,\PWM9/n24 }),
    .c({pnumcnt9[22],pnumcnt9[22]}),
    .clk(clk100m),
    .d({\PWM9/pnumr [22],\PWM9/pnumr [22]}),
    .mi({open_n16116,pwm_start_stop[25]}),
    .q({open_n16123,\PWM9/RemaTxNum[22]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg3_b23  (
    .a({_al_u2439_o,_al_u2439_o}),
    .b({\PWM9/n24 ,\PWM9/n24 }),
    .c({pnumcnt9[23],pnumcnt9[23]}),
    .clk(clk100m),
    .d({\PWM9/pnumr [23],\PWM9/pnumr [23]}),
    .mi({open_n16135,pwm_start_stop[25]}),
    .q({open_n16142,\PWM9/RemaTxNum[23]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg3_b5  (
    .a({_al_u2433_o,_al_u2433_o}),
    .b({\PWM9/n24 ,\PWM9/n24 }),
    .c({pnumcnt9[5],pnumcnt9[5]}),
    .clk(clk100m),
    .d({\PWM9/pnumr [5],\PWM9/pnumr [5]}),
    .mi({open_n16154,pwm_start_stop[25]}),
    .q({open_n16161,\PWM9/RemaTxNum[5]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg3_b6  (
    .a({_al_u2431_o,_al_u2431_o}),
    .b({\PWM9/n24 ,\PWM9/n24 }),
    .c({pnumcnt9[6],pnumcnt9[6]}),
    .clk(clk100m),
    .d({\PWM9/pnumr [6],\PWM9/pnumr [6]}),
    .mi({open_n16173,pwm_start_stop[25]}),
    .q({open_n16180,\PWM9/RemaTxNum[6]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWM9/reg3_b9  (
    .a({_al_u2425_o,_al_u2425_o}),
    .b({\PWM9/n24 ,\PWM9/n24 }),
    .c({pnumcnt9[9],pnumcnt9[9]}),
    .clk(clk100m),
    .d({\PWM9/pnumr [9],\PWM9/pnumr [9]}),
    .mi({open_n16192,pwm_start_stop[25]}),
    .q({open_n16199,\PWM9/RemaTxNum[9]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \PWM9/stopreq_reg  (
    .c({open_n16204,\PWM9/stopreq }),
    .clk(clk100m),
    .d({open_n16206,\PWM9/n0_lutinv }),
    .sr(pwm_start_stop[9]),
    .q({open_n16224,\PWM9/stopreq_keep }));  // src/OnePWM.v(15)
  EF2_PHY_LSLICE #(
    //.MACRO("PWM9/sub0/ucin_al_u3426"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM9/sub0/u11_al_u3429  (
    .a({\PWM9/FreCnt [13],\PWM9/FreCnt [11]}),
    .b({\PWM9/FreCnt [14],\PWM9/FreCnt [12]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM9/sub0/c11 ),
    .f({\PWM9/n12 [13],\PWM9/n12 [11]}),
    .fco(\PWM9/sub0/c15 ),
    .fx({\PWM9/n12 [14],\PWM9/n12 [12]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM9/sub0/ucin_al_u3426"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM9/sub0/u15_al_u3430  (
    .a({\PWM9/FreCnt [17],\PWM9/FreCnt [15]}),
    .b({\PWM9/FreCnt [18],\PWM9/FreCnt [16]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM9/sub0/c15 ),
    .f({\PWM9/n12 [17],\PWM9/n12 [15]}),
    .fco(\PWM9/sub0/c19 ),
    .fx({\PWM9/n12 [18],\PWM9/n12 [16]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM9/sub0/ucin_al_u3426"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM9/sub0/u19_al_u3431  (
    .a({\PWM9/FreCnt [21],\PWM9/FreCnt [19]}),
    .b({\PWM9/FreCnt [22],\PWM9/FreCnt [20]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM9/sub0/c19 ),
    .f({\PWM9/n12 [21],\PWM9/n12 [19]}),
    .fco(\PWM9/sub0/c23 ),
    .fx({\PWM9/n12 [22],\PWM9/n12 [20]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM9/sub0/ucin_al_u3426"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM9/sub0/u23_al_u3432  (
    .a({\PWM9/FreCnt [25],\PWM9/FreCnt [23]}),
    .b({\PWM9/FreCnt [26],\PWM9/FreCnt [24]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM9/sub0/c23 ),
    .f({\PWM9/n12 [25],\PWM9/n12 [23]}),
    .fx({\PWM9/n12 [26],\PWM9/n12 [24]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM9/sub0/ucin_al_u3426"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM9/sub0/u3_al_u3427  (
    .a({\PWM9/FreCnt [5],\PWM9/FreCnt [3]}),
    .b({\PWM9/FreCnt [6],\PWM9/FreCnt [4]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM9/sub0/c3 ),
    .f({\PWM9/n12 [5],\PWM9/n12 [3]}),
    .fco(\PWM9/sub0/c7 ),
    .fx({\PWM9/n12 [6],\PWM9/n12 [4]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM9/sub0/ucin_al_u3426"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM9/sub0/u7_al_u3428  (
    .a({\PWM9/FreCnt [9],\PWM9/FreCnt [7]}),
    .b({\PWM9/FreCnt [10],\PWM9/FreCnt [8]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWM9/sub0/c7 ),
    .f({\PWM9/n12 [9],\PWM9/n12 [7]}),
    .fco(\PWM9/sub0/c11 ),
    .fx({\PWM9/n12 [10],\PWM9/n12 [8]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWM9/sub0/ucin_al_u3426"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h0005),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWM9/sub0/ucin_al_u3426  (
    .a({\PWM9/FreCnt [1],1'b0}),
    .b({\PWM9/FreCnt [2],\PWM9/FreCnt [0]}),
    .c(2'b11),
    .d(2'b01),
    .e(2'b01),
    .f({\PWM9/n12 [1],open_n16351}),
    .fco(\PWM9/sub0/c3 ),
    .fx({\PWM9/n12 [2],\PWM9/n12 [0]}));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM9/sub1/u0|PWM9/sub1/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("SUB_CARRY"),
    .INIT_LUT0(16'b0000000000000101),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM9/sub1/u0|PWM9/sub1/ucin  (
    .a({pnumcnt9[0],1'b0}),
    .b({1'b1,open_n16354}),
    .f({\PWM9/n26 [0],open_n16374}),
    .fco(\PWM9/sub1/c1 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM9/sub1/u0|PWM9/sub1/ucin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM9/sub1/u10|PWM9/sub1/u9  (
    .a(pnumcnt9[10:9]),
    .b(2'b00),
    .fci(\PWM9/sub1/c9 ),
    .f(\PWM9/n26 [10:9]),
    .fco(\PWM9/sub1/c11 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM9/sub1/u0|PWM9/sub1/ucin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM9/sub1/u12|PWM9/sub1/u11  (
    .a(pnumcnt9[12:11]),
    .b(2'b00),
    .fci(\PWM9/sub1/c11 ),
    .f(\PWM9/n26 [12:11]),
    .fco(\PWM9/sub1/c13 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM9/sub1/u0|PWM9/sub1/ucin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM9/sub1/u14|PWM9/sub1/u13  (
    .a(pnumcnt9[14:13]),
    .b(2'b00),
    .fci(\PWM9/sub1/c13 ),
    .f(\PWM9/n26 [14:13]),
    .fco(\PWM9/sub1/c15 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM9/sub1/u0|PWM9/sub1/ucin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM9/sub1/u16|PWM9/sub1/u15  (
    .a(pnumcnt9[16:15]),
    .b(2'b00),
    .fci(\PWM9/sub1/c15 ),
    .f(\PWM9/n26 [16:15]),
    .fco(\PWM9/sub1/c17 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM9/sub1/u0|PWM9/sub1/ucin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM9/sub1/u18|PWM9/sub1/u17  (
    .a(pnumcnt9[18:17]),
    .b(2'b00),
    .fci(\PWM9/sub1/c17 ),
    .f(\PWM9/n26 [18:17]),
    .fco(\PWM9/sub1/c19 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM9/sub1/u0|PWM9/sub1/ucin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM9/sub1/u20|PWM9/sub1/u19  (
    .a(pnumcnt9[20:19]),
    .b(2'b00),
    .fci(\PWM9/sub1/c19 ),
    .f(\PWM9/n26 [20:19]),
    .fco(\PWM9/sub1/c21 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM9/sub1/u0|PWM9/sub1/ucin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM9/sub1/u22|PWM9/sub1/u21  (
    .a(pnumcnt9[22:21]),
    .b(2'b00),
    .fci(\PWM9/sub1/c21 ),
    .f(\PWM9/n26 [22:21]),
    .fco(\PWM9/sub1/c23 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM9/sub1/u0|PWM9/sub1/ucin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM9/sub1/u23_al_u3477  (
    .a({open_n16533,pnumcnt9[23]}),
    .b({open_n16534,1'b0}),
    .fci(\PWM9/sub1/c23 ),
    .f({open_n16553,\PWM9/n26 [23]}));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM9/sub1/u0|PWM9/sub1/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM9/sub1/u2|PWM9/sub1/u1  (
    .a(pnumcnt9[2:1]),
    .b(2'b00),
    .fci(\PWM9/sub1/c1 ),
    .f(\PWM9/n26 [2:1]),
    .fco(\PWM9/sub1/c3 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM9/sub1/u0|PWM9/sub1/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM9/sub1/u4|PWM9/sub1/u3  (
    .a(pnumcnt9[4:3]),
    .b(2'b00),
    .fci(\PWM9/sub1/c3 ),
    .f(\PWM9/n26 [4:3]),
    .fco(\PWM9/sub1/c5 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM9/sub1/u0|PWM9/sub1/ucin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM9/sub1/u6|PWM9/sub1/u5  (
    .a(pnumcnt9[6:5]),
    .b(2'b00),
    .fci(\PWM9/sub1/c5 ),
    .f(\PWM9/n26 [6:5]),
    .fco(\PWM9/sub1/c7 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWM9/sub1/u0|PWM9/sub1/ucin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWM9/sub1/u8|PWM9/sub1/u7  (
    .a(pnumcnt9[8:7]),
    .b(2'b00),
    .fci(\PWM9/sub1/c7 ),
    .f(\PWM9/n26 [8:7]),
    .fco(\PWM9/sub1/c9 ));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[0]  (
    .i(\PWMA/RemaTxNum[0]_keep ),
    .o(pnumcntA[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[10]  (
    .i(\PWMA/RemaTxNum[10]_keep ),
    .o(pnumcntA[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[11]  (
    .i(\PWMA/RemaTxNum[11]_keep ),
    .o(pnumcntA[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[12]  (
    .i(\PWMA/RemaTxNum[12]_keep ),
    .o(pnumcntA[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[13]  (
    .i(\PWMA/RemaTxNum[13]_keep ),
    .o(pnumcntA[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[14]  (
    .i(\PWMA/RemaTxNum[14]_keep ),
    .o(pnumcntA[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[15]  (
    .i(\PWMA/RemaTxNum[15]_keep ),
    .o(pnumcntA[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[16]  (
    .i(\PWMA/RemaTxNum[16]_keep ),
    .o(pnumcntA[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[17]  (
    .i(\PWMA/RemaTxNum[17]_keep ),
    .o(pnumcntA[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[18]  (
    .i(\PWMA/RemaTxNum[18]_keep ),
    .o(pnumcntA[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[19]  (
    .i(\PWMA/RemaTxNum[19]_keep ),
    .o(pnumcntA[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[1]  (
    .i(\PWMA/RemaTxNum[1]_keep ),
    .o(pnumcntA[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[20]  (
    .i(\PWMA/RemaTxNum[20]_keep ),
    .o(pnumcntA[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[21]  (
    .i(\PWMA/RemaTxNum[21]_keep ),
    .o(pnumcntA[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[22]  (
    .i(\PWMA/RemaTxNum[22]_keep ),
    .o(pnumcntA[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[23]  (
    .i(\PWMA/RemaTxNum[23]_keep ),
    .o(pnumcntA[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[2]  (
    .i(\PWMA/RemaTxNum[2]_keep ),
    .o(pnumcntA[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[3]  (
    .i(\PWMA/RemaTxNum[3]_keep ),
    .o(pnumcntA[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[4]  (
    .i(\PWMA/RemaTxNum[4]_keep ),
    .o(pnumcntA[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[5]  (
    .i(\PWMA/RemaTxNum[5]_keep ),
    .o(pnumcntA[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[6]  (
    .i(\PWMA/RemaTxNum[6]_keep ),
    .o(pnumcntA[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[7]  (
    .i(\PWMA/RemaTxNum[7]_keep ),
    .o(pnumcntA[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[8]  (
    .i(\PWMA/RemaTxNum[8]_keep ),
    .o(pnumcntA[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[9]  (
    .i(\PWMA/RemaTxNum[9]_keep ),
    .o(pnumcntA[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_dir  (
    .i(\PWMA/dir_keep ),
    .o(dir_pad[10]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[0]  (
    .i(\PWMA/pnumr[0]_keep ),
    .o(\PWMA/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[10]  (
    .i(\PWMA/pnumr[10]_keep ),
    .o(\PWMA/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[11]  (
    .i(\PWMA/pnumr[11]_keep ),
    .o(\PWMA/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[12]  (
    .i(\PWMA/pnumr[12]_keep ),
    .o(\PWMA/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[13]  (
    .i(\PWMA/pnumr[13]_keep ),
    .o(\PWMA/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[14]  (
    .i(\PWMA/pnumr[14]_keep ),
    .o(\PWMA/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[15]  (
    .i(\PWMA/pnumr[15]_keep ),
    .o(\PWMA/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[16]  (
    .i(\PWMA/pnumr[16]_keep ),
    .o(\PWMA/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[17]  (
    .i(\PWMA/pnumr[17]_keep ),
    .o(\PWMA/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[18]  (
    .i(\PWMA/pnumr[18]_keep ),
    .o(\PWMA/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[19]  (
    .i(\PWMA/pnumr[19]_keep ),
    .o(\PWMA/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[1]  (
    .i(\PWMA/pnumr[1]_keep ),
    .o(\PWMA/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[20]  (
    .i(\PWMA/pnumr[20]_keep ),
    .o(\PWMA/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[21]  (
    .i(\PWMA/pnumr[21]_keep ),
    .o(\PWMA/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[22]  (
    .i(\PWMA/pnumr[22]_keep ),
    .o(\PWMA/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[23]  (
    .i(\PWMA/pnumr[23]_keep ),
    .o(\PWMA/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[24]  (
    .i(\PWMA/pnumr[24]_keep ),
    .o(\PWMA/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[25]  (
    .i(\PWMA/pnumr[25]_keep ),
    .o(\PWMA/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[26]  (
    .i(\PWMA/pnumr[26]_keep ),
    .o(\PWMA/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[27]  (
    .i(\PWMA/pnumr[27]_keep ),
    .o(\PWMA/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[28]  (
    .i(\PWMA/pnumr[28]_keep ),
    .o(\PWMA/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[29]  (
    .i(\PWMA/pnumr[29]_keep ),
    .o(\PWMA/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[2]  (
    .i(\PWMA/pnumr[2]_keep ),
    .o(\PWMA/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[30]  (
    .i(\PWMA/pnumr[30]_keep ),
    .o(\PWMA/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[31]  (
    .i(\PWMA/pnumr[31]_keep ),
    .o(\PWMA/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[3]  (
    .i(\PWMA/pnumr[3]_keep ),
    .o(\PWMA/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[4]  (
    .i(\PWMA/pnumr[4]_keep ),
    .o(\PWMA/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[5]  (
    .i(\PWMA/pnumr[5]_keep ),
    .o(\PWMA/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[6]  (
    .i(\PWMA/pnumr[6]_keep ),
    .o(\PWMA/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[7]  (
    .i(\PWMA/pnumr[7]_keep ),
    .o(\PWMA/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[8]  (
    .i(\PWMA/pnumr[8]_keep ),
    .o(\PWMA/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[9]  (
    .i(\PWMA/pnumr[9]_keep ),
    .o(\PWMA/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pwm  (
    .i(\PWMA/pwm_keep ),
    .o(pwm_pad[10]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_stopreq  (
    .i(\PWMA/stopreq_keep ),
    .o(\PWMA/stopreq ));  // src/OnePWM.v(14)
  EF2_PHY_MSLICE #(
    //.LUT0("(D*~(C)*~((~0*~(B*A)))+D*C*~((~0*~(B*A)))+~(D)*C*(~0*~(B*A))+D*C*(~0*~(B*A)))"),
    //.LUT1("(D*~(C)*~((~1*~(B*A)))+D*C*~((~1*~(B*A)))+~(D)*C*(~1*~(B*A))+D*C*(~1*~(B*A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111100001110000),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMA/dir_reg  (
    .a({\PWMA/n24 ,\PWMA/n24 }),
    .b({\PWMA/n25_neg_lutinv ,\PWMA/n25_neg_lutinv }),
    .c({dir_pad[10],dir_pad[10]}),
    .clk(clk100m),
    .d({\PWMA/pnumr [31],\PWMA/pnumr [31]}),
    .mi({open_n16658,pwm_start_stop[26]}),
    .q({open_n16665,\PWMA/dir_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("~(~0*~(D*C*B*A))"),
    //.LUT1("~(~1*~(D*C*B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b1111111111111111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMA/pwm_reg  (
    .a({_al_u1538_o,_al_u1538_o}),
    .b({_al_u1545_o,_al_u1545_o}),
    .c({_al_u1547_o,_al_u1547_o}),
    .clk(clk100m),
    .d({_al_u1549_o,_al_u1549_o}),
    .mi({open_n16677,pwm_pad[10]}),
    .sr(\PWMA/u14_sel_is_1_o ),
    .q({open_n16683,\PWMA/pwm_keep }));  // src/OnePWM.v(45)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMA/reg0_b0|PWMA/reg0_b9  (
    .b({\PWMA/n12 [0],\PWMA/n12 [9]}),
    .c({freqA[0],freqA[9]}),
    .clk(clk100m),
    .d({\PWMA/n0_lutinv ,\PWMA/n0_lutinv }),
    .sr(\PWMA/n11 ),
    .q({\PWMA/FreCnt [0],\PWMA/FreCnt [9]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMA/reg0_b10|PWMA/reg0_b8  (
    .b({\PWMA/n12 [10],\PWMA/n12 [8]}),
    .c({freqA[10],freqA[8]}),
    .clk(clk100m),
    .d({\PWMA/n0_lutinv ,\PWMA/n0_lutinv }),
    .sr(\PWMA/n11 ),
    .q({\PWMA/FreCnt [10],\PWMA/FreCnt [8]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMA/reg0_b11|PWMA/reg0_b7  (
    .b({\PWMA/n12 [11],\PWMA/n12 [7]}),
    .c({freqA[11],freqA[7]}),
    .clk(clk100m),
    .d({\PWMA/n0_lutinv ,\PWMA/n0_lutinv }),
    .sr(\PWMA/n11 ),
    .q({\PWMA/FreCnt [11],\PWMA/FreCnt [7]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMA/reg0_b13|PWMA/reg0_b5  (
    .b({\PWMA/n12 [13],\PWMA/n12 [5]}),
    .c({freqA[13],freqA[5]}),
    .clk(clk100m),
    .d({\PWMA/n0_lutinv ,\PWMA/n0_lutinv }),
    .sr(\PWMA/n11 ),
    .q({\PWMA/FreCnt [13],\PWMA/FreCnt [5]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMA/reg0_b14|PWMA/reg0_b3  (
    .b({\PWMA/n12 [14],\PWMA/n12 [3]}),
    .c({freqA[14],freqA[3]}),
    .clk(clk100m),
    .d({\PWMA/n0_lutinv ,\PWMA/n0_lutinv }),
    .sr(\PWMA/n11 ),
    .q({\PWMA/FreCnt [14],\PWMA/FreCnt [3]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMA/reg0_b16|PWMA/reg0_b19  (
    .b({\PWMA/n12 [16],\PWMA/n12 [19]}),
    .c({freqA[16],freqA[19]}),
    .clk(clk100m),
    .d({\PWMA/n0_lutinv ,\PWMA/n0_lutinv }),
    .sr(\PWMA/n11 ),
    .q({\PWMA/FreCnt [16],\PWMA/FreCnt [19]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMA/reg0_b18|PWMA/reg0_b17  (
    .b(\PWMA/n12 [18:17]),
    .c(freqA[18:17]),
    .clk(clk100m),
    .d({\PWMA/n0_lutinv ,\PWMA/n0_lutinv }),
    .sr(\PWMA/n11 ),
    .q(\PWMA/FreCnt [18:17]));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMA/reg0_b20|PWMA/reg0_b6  (
    .b({\PWMA/n12 [20],\PWMA/n12 [6]}),
    .c({freqA[20],freqA[6]}),
    .clk(clk100m),
    .d({\PWMA/n0_lutinv ,\PWMA/n0_lutinv }),
    .sr(\PWMA/n11 ),
    .q({\PWMA/FreCnt [20],\PWMA/FreCnt [6]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMA/reg0_b21|PWMA/reg0_b4  (
    .b({\PWMA/n12 [21],\PWMA/n12 [4]}),
    .c({freqA[21],freqA[4]}),
    .clk(clk100m),
    .d({\PWMA/n0_lutinv ,\PWMA/n0_lutinv }),
    .sr(\PWMA/n11 ),
    .q({\PWMA/FreCnt [21],\PWMA/FreCnt [4]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMA/reg0_b22|PWMA/reg0_b26  (
    .b({\PWMA/n12 [22],\PWMA/n12 [26]}),
    .c({freqA[22],freqA[26]}),
    .clk(clk100m),
    .d({\PWMA/n0_lutinv ,\PWMA/n0_lutinv }),
    .sr(\PWMA/n11 ),
    .q({\PWMA/FreCnt [22],\PWMA/FreCnt [26]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMA/reg0_b24|PWMA/reg0_b25  (
    .b({\PWMA/n12 [24],\PWMA/n12 [25]}),
    .c({freqA[24],freqA[25]}),
    .clk(clk100m),
    .d({\PWMA/n0_lutinv ,\PWMA/n0_lutinv }),
    .sr(\PWMA/n11 ),
    .q({\PWMA/FreCnt [24],\PWMA/FreCnt [25]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(D*~B)*~(C*~A))"),
    //.LUT1("(~C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000110010101111),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMA/reg1_b10|PWMA/reg1_b20  (
    .a({open_n16928,\PWMA/FreCnt [17]}),
    .b({open_n16929,\PWMA/FreCnt [19]}),
    .c({\PWMA/FreCntr [10],\PWMA/FreCntr [18]}),
    .ce(\PWMA/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMA/FreCnt [9],\PWMA/FreCntr [20]}),
    .mi({freqA[10],freqA[20]}),
    .f({_al_u2558_o,_al_u2565_o}),
    .q({\PWMA/FreCntr [10],\PWMA/FreCntr [20]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(~(D*~B)*~(C*~A))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(~(D*~B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b1000110010101111),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000110010101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMA/reg1_b11|PWMA/reg1_b9  (
    .a({\PWMA/FreCnt [10],_al_u1535_o}),
    .b({\PWMA/FreCnt [5],\PWMA/FreCnt [11]}),
    .c({\PWMA/FreCntr [11],\PWMA/FreCnt [9]}),
    .ce(\PWMA/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMA/FreCntr [6],\PWMA/FreCntr [11]}),
    .e({open_n16944,\PWMA/FreCntr [9]}),
    .mi({freqA[11],freqA[9]}),
    .f({_al_u2567_o,_al_u1536_o}),
    .q({\PWMA/FreCntr [11],\PWMA/FreCntr [9]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1000010000100001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMA/reg1_b12|PWMA/reg1_b7  (
    .a({\PWMA/FreCnt [11],open_n16961}),
    .b({\PWMA/FreCnt [6],open_n16962}),
    .c({\PWMA/FreCntr [12],pwm_state_read[10]}),
    .ce(\PWMA/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMA/FreCntr [7],\PWMA/n0_lutinv }),
    .mi({freqA[12],freqA[7]}),
    .f({_al_u2571_o,\PWMA/n24 }),
    .q({\PWMA/FreCntr [12],\PWMA/FreCntr [7]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*~C)*~(D*~B))"),
    //.LUTF1("(~(D*~B)*~(~C*A))"),
    //.LUTG0("(A*~(1*~C)*~(D*~B))"),
    //.LUTG1("(~(D*~B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000100010101010),
    .INIT_LUTF1(16'b1100010011110101),
    .INIT_LUTG0(16'b1000000010100000),
    .INIT_LUTG1(16'b1100010011110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMA/reg1_b18|PWMA/reg1_b8  (
    .a({\PWMA/FreCnt [17],_al_u2573_o}),
    .b({\PWMA/FreCnt [8],\PWMA/FreCnt [13]}),
    .c({\PWMA/FreCntr [18],\PWMA/FreCnt [7]}),
    .ce(\PWMA/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMA/FreCntr [9],\PWMA/FreCntr [14]}),
    .e({open_n16977,\PWMA/FreCntr [8]}),
    .mi({freqA[18],freqA[8]}),
    .f({_al_u2573_o,_al_u2574_o}),
    .q({\PWMA/FreCntr [18],\PWMA/FreCntr [8]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(D@B)*~(C@A))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(~(D@B)*~(C@A))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000010000100001),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000010000100001),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMA/reg1_b22|PWMA/reg1_b15  (
    .a({\PWMA/FreCnt [22],\PWMA/FreCnt [14]}),
    .b({\PWMA/FreCnt [23],\PWMA/FreCnt [21]}),
    .c({\PWMA/FreCntr [22],\PWMA/FreCntr [15]}),
    .ce(\PWMA/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d(\PWMA/FreCntr [23:22]),
    .mi({freqA[22],freqA[15]}),
    .f({_al_u1533_o,_al_u2569_o}),
    .q({\PWMA/FreCntr [22],\PWMA/FreCntr [15]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(~0*C)*~(D*~B))"),
    //.LUTF1("(~(D*~B)*~(C*~A))"),
    //.LUTG0("(A*~(~1*C)*~(D*~B))"),
    //.LUTG1("(~(D*~B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000001010),
    .INIT_LUTF1(16'b1000110010101111),
    .INIT_LUTG0(16'b1000100010101010),
    .INIT_LUTG1(16'b1000110010101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMA/reg1_b24|PWMA/reg1_b13  (
    .a({\PWMA/FreCnt [23],_al_u2565_o}),
    .b({\PWMA/FreCnt [3],\PWMA/FreCnt [12]}),
    .c({\PWMA/FreCntr [24],\PWMA/FreCnt [23]}),
    .ce(\PWMA/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMA/FreCntr [4],\PWMA/FreCntr [13]}),
    .e({open_n17012,\PWMA/FreCntr [24]}),
    .mi({freqA[24],freqA[13]}),
    .f({_al_u2560_o,_al_u2566_o}),
    .q({\PWMA/FreCntr [24],\PWMA/FreCntr [13]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~C*~(0@B)*~(~D*A))"),
    //.LUTF1("(A*~(0@C)*~(D@B))"),
    //.LUTG0("(~C*~(1@B)*~(~D*A))"),
    //.LUTG1("(A*~(1@C)*~(D@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001100000001),
    .INIT_LUTF1(16'b0000100000000010),
    .INIT_LUTG0(16'b0000110000000100),
    .INIT_LUTG1(16'b1000000000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMA/reg1_b26|PWMA/reg1_b14  (
    .a({_al_u1546_o,\PWMA/FreCnt [13]}),
    .b({\PWMA/FreCnt [20],\PWMA/FreCnt [25]}),
    .c({\PWMA/FreCnt [26],\PWMA/FreCnt [26]}),
    .ce(\PWMA/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMA/FreCntr [20],\PWMA/FreCntr [14]}),
    .e({\PWMA/FreCntr [26],\PWMA/FreCntr [26]}),
    .mi({freqA[26],freqA[14]}),
    .f({_al_u1547_o,_al_u2575_o}),
    .q({\PWMA/FreCntr [26],\PWMA/FreCntr [14]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMA/reg1_b5|PWMA/reg1_b1  (
    .a({\PWMA/FreCnt [18],_al_u2563_o}),
    .b({\PWMA/FreCnt [5],\PWMA/FreCnt [0]}),
    .c({\PWMA/FreCntr [18],\PWMA/FreCnt [4]}),
    .ce(\PWMA/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMA/FreCntr [5],\PWMA/FreCntr [1]}),
    .e({open_n17045,\PWMA/FreCntr [5]}),
    .mi({freqA[5],freqA[1]}),
    .f({_al_u1537_o,_al_u2564_o}),
    .q({\PWMA/FreCntr [5],\PWMA/FreCntr [1]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~D*B)*~(C*~A))"),
    //.LUT1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111100100011),
    .INIT_LUT1(16'b1000010000100001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMA/reg1_b6|PWMA/reg1_b16  (
    .a({\PWMA/FreCnt [6],\PWMA/FreCnt [15]}),
    .b({\PWMA/FreCnt [7],\PWMA/FreCnt [5]}),
    .c({\PWMA/FreCntr [6],\PWMA/FreCntr [16]}),
    .ce(\PWMA/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d(\PWMA/FreCntr [7:6]),
    .mi({freqA[6],freqA[16]}),
    .f({_al_u1535_o,_al_u2562_o}),
    .q({\PWMA/FreCntr [6],\PWMA/FreCntr [16]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011100010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMA/reg2_b0|PWMA/reg2_b7  (
    .a({\PWMA/pnumr [0],\PWMA/pnumr [7]}),
    .b({pnumA[0],pnumA[32]}),
    .c({pnumA[32],pnumA[7]}),
    .clk(clk100m),
    .d({pwm_start_stop[26],pwm_start_stop[26]}),
    .q({\PWMA/pnumr[0]_keep ,\PWMA/pnumr[7]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMA/reg2_b10|PWMA/reg3_b10  (
    .a({\PWMA/pnumr [10],_al_u2549_o}),
    .b({pnumA[10],\PWMA/n24 }),
    .c({pnumA[32],pnumcntA[10]}),
    .clk(clk100m),
    .d({pwm_start_stop[26],\PWMA/pnumr [10]}),
    .e({open_n17096,pwm_start_stop[26]}),
    .q({\PWMA/pnumr[10]_keep ,\PWMA/RemaTxNum[10]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMA/reg2_b11|PWMA/reg3_b11  (
    .a({\PWMA/pnumr [11],_al_u2547_o}),
    .b({pnumA[11],\PWMA/n24 }),
    .c({pnumA[32],pnumcntA[11]}),
    .clk(clk100m),
    .d({pwm_start_stop[26],\PWMA/pnumr [11]}),
    .e({open_n17118,pwm_start_stop[26]}),
    .q({\PWMA/pnumr[11]_keep ,\PWMA/RemaTxNum[11]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011100010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMA/reg2_b12|PWMA/reg2_b6  (
    .a({\PWMA/pnumr [12],\PWMA/pnumr [6]}),
    .b({pnumA[12],pnumA[32]}),
    .c({pnumA[32],pnumA[6]}),
    .clk(clk100m),
    .d({pwm_start_stop[26],pwm_start_stop[26]}),
    .q({\PWMA/pnumr[12]_keep ,\PWMA/pnumr[6]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMA/reg2_b13|PWMA/reg2_b3  (
    .a({\PWMA/pnumr [13],\PWMA/pnumr [3]}),
    .b({pnumA[13],pnumA[3]}),
    .c({pnumA[32],pnumA[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[26],pwm_start_stop[26]}),
    .q({\PWMA/pnumr[13]_keep ,\PWMA/pnumr[3]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMA/reg2_b14|PWMA/reg3_b14  (
    .a({\PWMA/pnumr [14],_al_u2541_o}),
    .b({pnumA[14],\PWMA/n24 }),
    .c({pnumA[32],pnumcntA[14]}),
    .clk(clk100m),
    .d({pwm_start_stop[26],\PWMA/pnumr [14]}),
    .e({open_n17182,pwm_start_stop[26]}),
    .q({\PWMA/pnumr[14]_keep ,\PWMA/RemaTxNum[14]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMA/reg2_b15|PWMA/reg3_b15  (
    .a({\PWMA/pnumr [15],_al_u2539_o}),
    .b({pnumA[15],\PWMA/n24 }),
    .c({pnumA[32],pnumcntA[15]}),
    .clk(clk100m),
    .d({pwm_start_stop[26],\PWMA/pnumr [15]}),
    .e({open_n17204,pwm_start_stop[26]}),
    .q({\PWMA/pnumr[15]_keep ,\PWMA/RemaTxNum[15]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMA/reg2_b16|PWMA/reg2_b23  (
    .a({\PWMA/pnumr [16],\PWMA/pnumr [23]}),
    .b({pnumA[16],pnumA[23]}),
    .c({pnumA[32],pnumA[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[26],pwm_start_stop[26]}),
    .q({\PWMA/pnumr[16]_keep ,\PWMA/pnumr[23]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMA/reg2_b17|PWMA/reg2_b20  (
    .a({\PWMA/pnumr [17],\PWMA/pnumr [20]}),
    .b({pnumA[17],pnumA[20]}),
    .c({pnumA[32],pnumA[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[26],pwm_start_stop[26]}),
    .q({\PWMA/pnumr[17]_keep ,\PWMA/pnumr[20]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMA/reg2_b18|PWMA/reg3_b18  (
    .a({\PWMA/pnumr [18],_al_u2533_o}),
    .b({pnumA[18],\PWMA/n24 }),
    .c({pnumA[32],pnumcntA[18]}),
    .clk(clk100m),
    .d({pwm_start_stop[26],\PWMA/pnumr [18]}),
    .e({open_n17268,pwm_start_stop[26]}),
    .q({\PWMA/pnumr[18]_keep ,\PWMA/RemaTxNum[18]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMA/reg2_b19|PWMA/reg3_b19  (
    .a({\PWMA/pnumr [19],_al_u2531_o}),
    .b({pnumA[19],\PWMA/n24 }),
    .c({pnumA[32],pnumcntA[19]}),
    .clk(clk100m),
    .d({pwm_start_stop[26],\PWMA/pnumr [19]}),
    .e({open_n17290,pwm_start_stop[26]}),
    .q({\PWMA/pnumr[19]_keep ,\PWMA/RemaTxNum[19]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMA/reg2_b1|PWMA/reg2_b2  (
    .a({\PWMA/pnumr [1],\PWMA/pnumr [2]}),
    .b({pnumA[1],pnumA[2]}),
    .c({pnumA[32],pnumA[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[26],pwm_start_stop[26]}),
    .q({\PWMA/pnumr[1]_keep ,\PWMA/pnumr[2]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMA/reg2_b21|PWMA/reg3_b21  (
    .a({\PWMA/pnumr [21],_al_u2525_o}),
    .b({pnumA[21],\PWMA/n24 }),
    .c({pnumA[32],pnumcntA[21]}),
    .clk(clk100m),
    .d({pwm_start_stop[26],\PWMA/pnumr [21]}),
    .e({open_n17331,pwm_start_stop[26]}),
    .q({\PWMA/pnumr[21]_keep ,\PWMA/RemaTxNum[21]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMA/reg2_b22|PWMA/reg3_b22  (
    .a({\PWMA/pnumr [22],_al_u2523_o}),
    .b({pnumA[22],\PWMA/n24 }),
    .c({pnumA[32],pnumcntA[22]}),
    .clk(clk100m),
    .d({pwm_start_stop[26],\PWMA/pnumr [22]}),
    .e({open_n17353,pwm_start_stop[26]}),
    .q({\PWMA/pnumr[22]_keep ,\PWMA/RemaTxNum[22]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMA/reg2_b24|PWMA/reg2_b31  (
    .a({\PWMA/pnumr [24],\PWMA/pnumr [31]}),
    .b({pnumA[24],pnumA[31]}),
    .c({pnumA[32],pnumA[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[26],pwm_start_stop[26]}),
    .q({\PWMA/pnumr[24]_keep ,\PWMA/pnumr[31]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMA/reg2_b25|PWMA/reg2_b30  (
    .a({\PWMA/pnumr [25],\PWMA/pnumr [30]}),
    .b({pnumA[25],pnumA[30]}),
    .c({pnumA[32],pnumA[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[26],pwm_start_stop[26]}),
    .q({\PWMA/pnumr[25]_keep ,\PWMA/pnumr[30]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMA/reg2_b26|PWMA/reg2_b29  (
    .a({\PWMA/pnumr [26],\PWMA/pnumr [29]}),
    .b({pnumA[26],pnumA[29]}),
    .c({pnumA[32],pnumA[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[26],pwm_start_stop[26]}),
    .q({\PWMA/pnumr[26]_keep ,\PWMA/pnumr[29]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMA/reg2_b27|PWMA/reg2_b28  (
    .a({\PWMA/pnumr [27],\PWMA/pnumr [28]}),
    .b({pnumA[27],pnumA[28]}),
    .c({pnumA[32],pnumA[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[26],pwm_start_stop[26]}),
    .q({\PWMA/pnumr[27]_keep ,\PWMA/pnumr[28]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMA/reg2_b4|PWMA/reg3_b4  (
    .a({\PWMA/pnumr [4],_al_u2517_o}),
    .b({pnumA[32],\PWMA/n24 }),
    .c({pnumA[4],pnumcntA[4]}),
    .clk(clk100m),
    .d({pwm_start_stop[26],\PWMA/pnumr [4]}),
    .e({open_n17455,pwm_start_stop[26]}),
    .q({\PWMA/pnumr[4]_keep ,\PWMA/RemaTxNum[4]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMA/reg2_b5|PWMA/reg3_b5  (
    .a({\PWMA/pnumr [5],_al_u2515_o}),
    .b({pnumA[32],\PWMA/n24 }),
    .c({pnumA[5],pnumcntA[5]}),
    .clk(clk100m),
    .d({pwm_start_stop[26],\PWMA/pnumr [5]}),
    .e({open_n17477,pwm_start_stop[26]}),
    .q({\PWMA/pnumr[5]_keep ,\PWMA/RemaTxNum[5]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMA/reg2_b8|PWMA/reg3_b8  (
    .a({\PWMA/pnumr [8],_al_u2509_o}),
    .b({pnumA[32],\PWMA/n24 }),
    .c({pnumA[8],pnumcntA[8]}),
    .clk(clk100m),
    .d({pwm_start_stop[26],\PWMA/pnumr [8]}),
    .e({open_n17499,pwm_start_stop[26]}),
    .q({\PWMA/pnumr[8]_keep ,\PWMA/RemaTxNum[8]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMA/reg2_b9|PWMA/reg3_b9  (
    .a({\PWMA/pnumr [9],_al_u2507_o}),
    .b({pnumA[32],\PWMA/n24 }),
    .c({pnumA[9],pnumcntA[9]}),
    .clk(clk100m),
    .d({pwm_start_stop[26],\PWMA/pnumr [9]}),
    .e({open_n17521,pwm_start_stop[26]}),
    .q({\PWMA/pnumr[9]_keep ,\PWMA/RemaTxNum[9]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMA/reg3_b0  (
    .a({_al_u2553_o,_al_u2553_o}),
    .b({\PWMA/n24 ,\PWMA/n24 }),
    .c({pnumcntA[0],pnumcntA[0]}),
    .clk(clk100m),
    .d({\PWMA/pnumr [0],\PWMA/pnumr [0]}),
    .mi({open_n17553,pwm_start_stop[26]}),
    .q({open_n17560,\PWMA/RemaTxNum[0]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMA/reg3_b1  (
    .a({_al_u2551_o,_al_u2551_o}),
    .b({\PWMA/n24 ,\PWMA/n24 }),
    .c({pnumcntA[1],pnumcntA[1]}),
    .clk(clk100m),
    .d({\PWMA/pnumr [1],\PWMA/pnumr [1]}),
    .mi({open_n17572,pwm_start_stop[26]}),
    .q({open_n17579,\PWMA/RemaTxNum[1]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMA/reg3_b12  (
    .a({_al_u2545_o,_al_u2545_o}),
    .b({\PWMA/n24 ,\PWMA/n24 }),
    .c({pnumcntA[12],pnumcntA[12]}),
    .clk(clk100m),
    .d({\PWMA/pnumr [12],\PWMA/pnumr [12]}),
    .mi({open_n17591,pwm_start_stop[26]}),
    .q({open_n17598,\PWMA/RemaTxNum[12]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMA/reg3_b13  (
    .a({_al_u2543_o,_al_u2543_o}),
    .b({\PWMA/n24 ,\PWMA/n24 }),
    .c({pnumcntA[13],pnumcntA[13]}),
    .clk(clk100m),
    .d({\PWMA/pnumr [13],\PWMA/pnumr [13]}),
    .mi({open_n17610,pwm_start_stop[26]}),
    .q({open_n17617,\PWMA/RemaTxNum[13]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMA/reg3_b16  (
    .a({_al_u2537_o,_al_u2537_o}),
    .b({\PWMA/n24 ,\PWMA/n24 }),
    .c({pnumcntA[16],pnumcntA[16]}),
    .clk(clk100m),
    .d({\PWMA/pnumr [16],\PWMA/pnumr [16]}),
    .mi({open_n17629,pwm_start_stop[26]}),
    .q({open_n17636,\PWMA/RemaTxNum[16]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMA/reg3_b17  (
    .a({_al_u2535_o,_al_u2535_o}),
    .b({\PWMA/n24 ,\PWMA/n24 }),
    .c({pnumcntA[17],pnumcntA[17]}),
    .clk(clk100m),
    .d({\PWMA/pnumr [17],\PWMA/pnumr [17]}),
    .mi({open_n17648,pwm_start_stop[26]}),
    .q({open_n17655,\PWMA/RemaTxNum[17]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMA/reg3_b2  (
    .a({_al_u2529_o,_al_u2529_o}),
    .b({\PWMA/n24 ,\PWMA/n24 }),
    .c({pnumcntA[2],pnumcntA[2]}),
    .clk(clk100m),
    .d({\PWMA/pnumr [2],\PWMA/pnumr [2]}),
    .mi({open_n17667,pwm_start_stop[26]}),
    .q({open_n17674,\PWMA/RemaTxNum[2]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMA/reg3_b20  (
    .a({_al_u2527_o,_al_u2527_o}),
    .b({\PWMA/n24 ,\PWMA/n24 }),
    .c({pnumcntA[20],pnumcntA[20]}),
    .clk(clk100m),
    .d({\PWMA/pnumr [20],\PWMA/pnumr [20]}),
    .mi({open_n17686,pwm_start_stop[26]}),
    .q({open_n17693,\PWMA/RemaTxNum[20]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMA/reg3_b23  (
    .a({_al_u2521_o,_al_u2521_o}),
    .b({\PWMA/n24 ,\PWMA/n24 }),
    .c({pnumcntA[23],pnumcntA[23]}),
    .clk(clk100m),
    .d({\PWMA/pnumr [23],\PWMA/pnumr [23]}),
    .mi({open_n17705,pwm_start_stop[26]}),
    .q({open_n17712,\PWMA/RemaTxNum[23]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMA/reg3_b3  (
    .a({_al_u2519_o,_al_u2519_o}),
    .b({\PWMA/n24 ,\PWMA/n24 }),
    .c({pnumcntA[3],pnumcntA[3]}),
    .clk(clk100m),
    .d({\PWMA/pnumr [3],\PWMA/pnumr [3]}),
    .mi({open_n17724,pwm_start_stop[26]}),
    .q({open_n17731,\PWMA/RemaTxNum[3]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMA/reg3_b6  (
    .a({_al_u2513_o,_al_u2513_o}),
    .b({\PWMA/n24 ,\PWMA/n24 }),
    .c({pnumcntA[6],pnumcntA[6]}),
    .clk(clk100m),
    .d({\PWMA/pnumr [6],\PWMA/pnumr [6]}),
    .mi({open_n17743,pwm_start_stop[26]}),
    .q({open_n17750,\PWMA/RemaTxNum[6]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMA/reg3_b7  (
    .a({_al_u2511_o,_al_u2511_o}),
    .b({\PWMA/n24 ,\PWMA/n24 }),
    .c({pnumcntA[7],pnumcntA[7]}),
    .clk(clk100m),
    .d({\PWMA/pnumr [7],\PWMA/pnumr [7]}),
    .mi({open_n17762,pwm_start_stop[26]}),
    .q({open_n17769,\PWMA/RemaTxNum[7]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \PWMA/stopreq_reg  (
    .c({open_n17774,\PWMA/stopreq }),
    .clk(clk100m),
    .d({open_n17776,\PWMA/n0_lutinv }),
    .sr(pwm_start_stop[10]),
    .q({open_n17794,\PWMA/stopreq_keep }));  // src/OnePWM.v(15)
  EF2_PHY_LSLICE #(
    //.MACRO("PWMA/sub0/ucin_al_u3433"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWMA/sub0/u11_al_u3436  (
    .a({\PWMA/FreCnt [13],\PWMA/FreCnt [11]}),
    .b({\PWMA/FreCnt [14],\PWMA/FreCnt [12]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWMA/sub0/c11 ),
    .f({\PWMA/n12 [13],\PWMA/n12 [11]}),
    .fco(\PWMA/sub0/c15 ),
    .fx({\PWMA/n12 [14],\PWMA/n12 [12]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWMA/sub0/ucin_al_u3433"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWMA/sub0/u15_al_u3437  (
    .a({\PWMA/FreCnt [17],\PWMA/FreCnt [15]}),
    .b({\PWMA/FreCnt [18],\PWMA/FreCnt [16]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWMA/sub0/c15 ),
    .f({\PWMA/n12 [17],\PWMA/n12 [15]}),
    .fco(\PWMA/sub0/c19 ),
    .fx({\PWMA/n12 [18],\PWMA/n12 [16]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWMA/sub0/ucin_al_u3433"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWMA/sub0/u19_al_u3438  (
    .a({\PWMA/FreCnt [21],\PWMA/FreCnt [19]}),
    .b({\PWMA/FreCnt [22],\PWMA/FreCnt [20]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWMA/sub0/c19 ),
    .f({\PWMA/n12 [21],\PWMA/n12 [19]}),
    .fco(\PWMA/sub0/c23 ),
    .fx({\PWMA/n12 [22],\PWMA/n12 [20]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWMA/sub0/ucin_al_u3433"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWMA/sub0/u23_al_u3439  (
    .a({\PWMA/FreCnt [25],\PWMA/FreCnt [23]}),
    .b({\PWMA/FreCnt [26],\PWMA/FreCnt [24]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWMA/sub0/c23 ),
    .f({\PWMA/n12 [25],\PWMA/n12 [23]}),
    .fx({\PWMA/n12 [26],\PWMA/n12 [24]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWMA/sub0/ucin_al_u3433"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWMA/sub0/u3_al_u3434  (
    .a({\PWMA/FreCnt [5],\PWMA/FreCnt [3]}),
    .b({\PWMA/FreCnt [6],\PWMA/FreCnt [4]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWMA/sub0/c3 ),
    .f({\PWMA/n12 [5],\PWMA/n12 [3]}),
    .fco(\PWMA/sub0/c7 ),
    .fx({\PWMA/n12 [6],\PWMA/n12 [4]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWMA/sub0/ucin_al_u3433"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWMA/sub0/u7_al_u3435  (
    .a({\PWMA/FreCnt [9],\PWMA/FreCnt [7]}),
    .b({\PWMA/FreCnt [10],\PWMA/FreCnt [8]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWMA/sub0/c7 ),
    .f({\PWMA/n12 [9],\PWMA/n12 [7]}),
    .fco(\PWMA/sub0/c11 ),
    .fx({\PWMA/n12 [10],\PWMA/n12 [8]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWMA/sub0/ucin_al_u3433"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h0005),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWMA/sub0/ucin_al_u3433  (
    .a({\PWMA/FreCnt [1],1'b0}),
    .b({\PWMA/FreCnt [2],\PWMA/FreCnt [0]}),
    .c(2'b11),
    .d(2'b01),
    .e(2'b01),
    .f({\PWMA/n12 [1],open_n17921}),
    .fco(\PWMA/sub0/c3 ),
    .fx({\PWMA/n12 [2],\PWMA/n12 [0]}));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMA/sub1/u0|PWMA/sub1/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("SUB_CARRY"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000101),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMA/sub1/u0|PWMA/sub1/ucin  (
    .a({pnumcntA[0],1'b0}),
    .b({1'b1,open_n17924}),
    .clk(clk100m),
    .mi(\U_AHB/h2h_hwdata [30:29]),
    .sr(\U_AHB/n63 ),
    .f({\PWMA/n26 [0],open_n17940}),
    .fco(\PWMA/sub1/c1 ),
    .q(pnum8[30:29]));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMA/sub1/u0|PWMA/sub1/ucin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMA/sub1/u10|PWMA/sub1/u9  (
    .a(pnumcntA[10:9]),
    .b(2'b00),
    .fci(\PWMA/sub1/c9 ),
    .f(\PWMA/n26 [10:9]),
    .fco(\PWMA/sub1/c11 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMA/sub1/u0|PWMA/sub1/ucin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMA/sub1/u12|PWMA/sub1/u11  (
    .a(pnumcntA[12:11]),
    .b(2'b00),
    .fci(\PWMA/sub1/c11 ),
    .f(\PWMA/n26 [12:11]),
    .fco(\PWMA/sub1/c13 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMA/sub1/u0|PWMA/sub1/ucin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMA/sub1/u14|PWMA/sub1/u13  (
    .a(pnumcntA[14:13]),
    .b(2'b00),
    .fci(\PWMA/sub1/c13 ),
    .f(\PWMA/n26 [14:13]),
    .fco(\PWMA/sub1/c15 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMA/sub1/u0|PWMA/sub1/ucin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMA/sub1/u16|PWMA/sub1/u15  (
    .a(pnumcntA[16:15]),
    .b(2'b00),
    .fci(\PWMA/sub1/c15 ),
    .f(\PWMA/n26 [16:15]),
    .fco(\PWMA/sub1/c17 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMA/sub1/u0|PWMA/sub1/ucin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMA/sub1/u18|PWMA/sub1/u17  (
    .a(pnumcntA[18:17]),
    .b(2'b00),
    .fci(\PWMA/sub1/c17 ),
    .f(\PWMA/n26 [18:17]),
    .fco(\PWMA/sub1/c19 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMA/sub1/u0|PWMA/sub1/ucin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMA/sub1/u20|PWMA/sub1/u19  (
    .a(pnumcntA[20:19]),
    .b(2'b00),
    .fci(\PWMA/sub1/c19 ),
    .f(\PWMA/n26 [20:19]),
    .fco(\PWMA/sub1/c21 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMA/sub1/u0|PWMA/sub1/ucin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMA/sub1/u22|PWMA/sub1/u21  (
    .a(pnumcntA[22:21]),
    .b(2'b00),
    .fci(\PWMA/sub1/c21 ),
    .f(\PWMA/n26 [22:21]),
    .fco(\PWMA/sub1/c23 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMA/sub1/u0|PWMA/sub1/ucin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMA/sub1/u23_al_u3478  (
    .a({open_n18097,pnumcntA[23]}),
    .b({open_n18098,1'b0}),
    .fci(\PWMA/sub1/c23 ),
    .f({open_n18117,\PWMA/n26 [23]}));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMA/sub1/u0|PWMA/sub1/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMA/sub1/u2|PWMA/sub1/u1  (
    .a(pnumcntA[2:1]),
    .b(2'b00),
    .fci(\PWMA/sub1/c1 ),
    .f(\PWMA/n26 [2:1]),
    .fco(\PWMA/sub1/c3 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMA/sub1/u0|PWMA/sub1/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMA/sub1/u4|PWMA/sub1/u3  (
    .a(pnumcntA[4:3]),
    .b(2'b00),
    .fci(\PWMA/sub1/c3 ),
    .f(\PWMA/n26 [4:3]),
    .fco(\PWMA/sub1/c5 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMA/sub1/u0|PWMA/sub1/ucin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMA/sub1/u6|PWMA/sub1/u5  (
    .a(pnumcntA[6:5]),
    .b(2'b00),
    .fci(\PWMA/sub1/c5 ),
    .f(\PWMA/n26 [6:5]),
    .fco(\PWMA/sub1/c7 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMA/sub1/u0|PWMA/sub1/ucin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMA/sub1/u8|PWMA/sub1/u7  (
    .a(pnumcntA[8:7]),
    .b(2'b00),
    .fci(\PWMA/sub1/c7 ),
    .f(\PWMA/n26 [8:7]),
    .fco(\PWMA/sub1/c9 ));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[0]  (
    .i(\PWMB/RemaTxNum[0]_keep ),
    .o(pnumcntB[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[10]  (
    .i(\PWMB/RemaTxNum[10]_keep ),
    .o(pnumcntB[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[11]  (
    .i(\PWMB/RemaTxNum[11]_keep ),
    .o(pnumcntB[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[12]  (
    .i(\PWMB/RemaTxNum[12]_keep ),
    .o(pnumcntB[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[13]  (
    .i(\PWMB/RemaTxNum[13]_keep ),
    .o(pnumcntB[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[14]  (
    .i(\PWMB/RemaTxNum[14]_keep ),
    .o(pnumcntB[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[15]  (
    .i(\PWMB/RemaTxNum[15]_keep ),
    .o(pnumcntB[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[16]  (
    .i(\PWMB/RemaTxNum[16]_keep ),
    .o(pnumcntB[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[17]  (
    .i(\PWMB/RemaTxNum[17]_keep ),
    .o(pnumcntB[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[18]  (
    .i(\PWMB/RemaTxNum[18]_keep ),
    .o(pnumcntB[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[19]  (
    .i(\PWMB/RemaTxNum[19]_keep ),
    .o(pnumcntB[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[1]  (
    .i(\PWMB/RemaTxNum[1]_keep ),
    .o(pnumcntB[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[20]  (
    .i(\PWMB/RemaTxNum[20]_keep ),
    .o(pnumcntB[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[21]  (
    .i(\PWMB/RemaTxNum[21]_keep ),
    .o(pnumcntB[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[22]  (
    .i(\PWMB/RemaTxNum[22]_keep ),
    .o(pnumcntB[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[23]  (
    .i(\PWMB/RemaTxNum[23]_keep ),
    .o(pnumcntB[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[2]  (
    .i(\PWMB/RemaTxNum[2]_keep ),
    .o(pnumcntB[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[3]  (
    .i(\PWMB/RemaTxNum[3]_keep ),
    .o(pnumcntB[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[4]  (
    .i(\PWMB/RemaTxNum[4]_keep ),
    .o(pnumcntB[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[5]  (
    .i(\PWMB/RemaTxNum[5]_keep ),
    .o(pnumcntB[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[6]  (
    .i(\PWMB/RemaTxNum[6]_keep ),
    .o(pnumcntB[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[7]  (
    .i(\PWMB/RemaTxNum[7]_keep ),
    .o(pnumcntB[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[8]  (
    .i(\PWMB/RemaTxNum[8]_keep ),
    .o(pnumcntB[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[9]  (
    .i(\PWMB/RemaTxNum[9]_keep ),
    .o(pnumcntB[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_dir  (
    .i(\PWMB/dir_keep ),
    .o(dir_pad[11]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[0]  (
    .i(\PWMB/pnumr[0]_keep ),
    .o(\PWMB/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[10]  (
    .i(\PWMB/pnumr[10]_keep ),
    .o(\PWMB/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[11]  (
    .i(\PWMB/pnumr[11]_keep ),
    .o(\PWMB/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[12]  (
    .i(\PWMB/pnumr[12]_keep ),
    .o(\PWMB/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[13]  (
    .i(\PWMB/pnumr[13]_keep ),
    .o(\PWMB/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[14]  (
    .i(\PWMB/pnumr[14]_keep ),
    .o(\PWMB/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[15]  (
    .i(\PWMB/pnumr[15]_keep ),
    .o(\PWMB/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[16]  (
    .i(\PWMB/pnumr[16]_keep ),
    .o(\PWMB/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[17]  (
    .i(\PWMB/pnumr[17]_keep ),
    .o(\PWMB/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[18]  (
    .i(\PWMB/pnumr[18]_keep ),
    .o(\PWMB/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[19]  (
    .i(\PWMB/pnumr[19]_keep ),
    .o(\PWMB/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[1]  (
    .i(\PWMB/pnumr[1]_keep ),
    .o(\PWMB/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[20]  (
    .i(\PWMB/pnumr[20]_keep ),
    .o(\PWMB/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[21]  (
    .i(\PWMB/pnumr[21]_keep ),
    .o(\PWMB/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[22]  (
    .i(\PWMB/pnumr[22]_keep ),
    .o(\PWMB/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[23]  (
    .i(\PWMB/pnumr[23]_keep ),
    .o(\PWMB/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[24]  (
    .i(\PWMB/pnumr[24]_keep ),
    .o(\PWMB/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[25]  (
    .i(\PWMB/pnumr[25]_keep ),
    .o(\PWMB/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[26]  (
    .i(\PWMB/pnumr[26]_keep ),
    .o(\PWMB/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[27]  (
    .i(\PWMB/pnumr[27]_keep ),
    .o(\PWMB/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[28]  (
    .i(\PWMB/pnumr[28]_keep ),
    .o(\PWMB/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[29]  (
    .i(\PWMB/pnumr[29]_keep ),
    .o(\PWMB/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[2]  (
    .i(\PWMB/pnumr[2]_keep ),
    .o(\PWMB/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[30]  (
    .i(\PWMB/pnumr[30]_keep ),
    .o(\PWMB/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[31]  (
    .i(\PWMB/pnumr[31]_keep ),
    .o(\PWMB/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[3]  (
    .i(\PWMB/pnumr[3]_keep ),
    .o(\PWMB/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[4]  (
    .i(\PWMB/pnumr[4]_keep ),
    .o(\PWMB/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[5]  (
    .i(\PWMB/pnumr[5]_keep ),
    .o(\PWMB/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[6]  (
    .i(\PWMB/pnumr[6]_keep ),
    .o(\PWMB/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[7]  (
    .i(\PWMB/pnumr[7]_keep ),
    .o(\PWMB/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[8]  (
    .i(\PWMB/pnumr[8]_keep ),
    .o(\PWMB/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[9]  (
    .i(\PWMB/pnumr[9]_keep ),
    .o(\PWMB/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pwm  (
    .i(\PWMB/pwm_keep ),
    .o(pwm_pad[11]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_stopreq  (
    .i(\PWMB/stopreq_keep ),
    .o(\PWMB/stopreq ));  // src/OnePWM.v(14)
  EF2_PHY_MSLICE #(
    //.LUT0("(D*~(C)*~((~0*~(B*A)))+D*C*~((~0*~(B*A)))+~(D)*C*(~0*~(B*A))+D*C*(~0*~(B*A)))"),
    //.LUT1("(D*~(C)*~((~1*~(B*A)))+D*C*~((~1*~(B*A)))+~(D)*C*(~1*~(B*A))+D*C*(~1*~(B*A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111100001110000),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/dir_reg  (
    .a({\PWMB/n24 ,\PWMB/n24 }),
    .b({\PWMB/n25_neg_lutinv ,\PWMB/n25_neg_lutinv }),
    .c({dir_pad[11],dir_pad[11]}),
    .clk(clk100m),
    .d({\PWMB/pnumr [31],\PWMB/pnumr [31]}),
    .mi({open_n18222,pwm_start_stop[27]}),
    .q({open_n18229,\PWMB/dir_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("~(~0*~(D*C*B*A))"),
    //.LUT1("~(~1*~(D*C*B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b1111111111111111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMB/pwm_reg  (
    .a({_al_u1556_o,_al_u1556_o}),
    .b({_al_u1562_o,_al_u1562_o}),
    .c({_al_u1564_o,_al_u1564_o}),
    .clk(clk100m),
    .d({_al_u1566_o,_al_u1566_o}),
    .mi({open_n18241,pwm_pad[11]}),
    .sr(\PWMB/u14_sel_is_1_o ),
    .q({open_n18247,\PWMB/pwm_keep }));  // src/OnePWM.v(45)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMB/reg0_b0|PWMB/reg0_b15  (
    .b({\PWMB/n12 [0],\PWMB/n12 [15]}),
    .c({freqB[0],freqB[15]}),
    .clk(clk100m),
    .d({\PWMB/n0_lutinv ,\PWMB/n0_lutinv }),
    .sr(\PWMB/n11 ),
    .q({\PWMB/FreCnt [0],\PWMB/FreCnt [15]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMB/reg0_b10|PWMB/reg0_b9  (
    .b(\PWMB/n12 [10:9]),
    .c(freqB[10:9]),
    .clk(clk100m),
    .d({\PWMB/n0_lutinv ,\PWMB/n0_lutinv }),
    .sr(\PWMB/n11 ),
    .q(\PWMB/FreCnt [10:9]));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMB/reg0_b11|PWMB/reg0_b8  (
    .b({\PWMB/n12 [11],\PWMB/n12 [8]}),
    .c({freqB[11],freqB[8]}),
    .clk(clk100m),
    .d({\PWMB/n0_lutinv ,\PWMB/n0_lutinv }),
    .sr(\PWMB/n11 ),
    .q({\PWMB/FreCnt [11],\PWMB/FreCnt [8]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMB/reg0_b12|PWMB/reg0_b7  (
    .b({\PWMB/n12 [12],\PWMB/n12 [7]}),
    .c({freqB[12],freqB[7]}),
    .clk(clk100m),
    .d({\PWMB/n0_lutinv ,\PWMB/n0_lutinv }),
    .sr(\PWMB/n11 ),
    .q({\PWMB/FreCnt [12],\PWMB/FreCnt [7]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMB/reg0_b13|PWMB/reg0_b5  (
    .b({\PWMB/n12 [13],\PWMB/n12 [5]}),
    .c({freqB[13],freqB[5]}),
    .clk(clk100m),
    .d({\PWMB/n0_lutinv ,\PWMB/n0_lutinv }),
    .sr(\PWMB/n11 ),
    .q({\PWMB/FreCnt [13],\PWMB/FreCnt [5]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMB/reg0_b14|PWMB/reg0_b3  (
    .b({\PWMB/n12 [14],\PWMB/n12 [3]}),
    .c({freqB[14],freqB[3]}),
    .clk(clk100m),
    .d({\PWMB/n0_lutinv ,\PWMB/n0_lutinv }),
    .sr(\PWMB/n11 ),
    .q({\PWMB/FreCnt [14],\PWMB/FreCnt [3]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMB/reg0_b16|PWMB/reg0_b25  (
    .b({\PWMB/n12 [16],\PWMB/n12 [25]}),
    .c({freqB[16],freqB[25]}),
    .clk(clk100m),
    .d({\PWMB/n0_lutinv ,\PWMB/n0_lutinv }),
    .sr(\PWMB/n11 ),
    .q({\PWMB/FreCnt [16],\PWMB/FreCnt [25]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMB/reg0_b17|PWMB/reg0_b23  (
    .b({\PWMB/n12 [17],\PWMB/n12 [23]}),
    .c({freqB[17],freqB[23]}),
    .clk(clk100m),
    .d({\PWMB/n0_lutinv ,\PWMB/n0_lutinv }),
    .sr(\PWMB/n11 ),
    .q({\PWMB/FreCnt [17],\PWMB/FreCnt [23]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMB/reg0_b18|PWMB/reg0_b21  (
    .b({\PWMB/n12 [18],\PWMB/n12 [21]}),
    .c({freqB[18],freqB[21]}),
    .clk(clk100m),
    .d({\PWMB/n0_lutinv ,\PWMB/n0_lutinv }),
    .sr(\PWMB/n11 ),
    .q({\PWMB/FreCnt [18],\PWMB/FreCnt [21]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMB/reg0_b20|PWMB/reg0_b1  (
    .b({\PWMB/n12 [20],\PWMB/n12 [1]}),
    .c({freqB[20],freqB[1]}),
    .clk(clk100m),
    .d({\PWMB/n0_lutinv ,\PWMB/n0_lutinv }),
    .sr(\PWMB/n11 ),
    .q({\PWMB/FreCnt [20],\PWMB/FreCnt [1]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMB/reg0_b22|PWMB/reg0_b6  (
    .b({\PWMB/n12 [22],\PWMB/n12 [6]}),
    .c({freqB[22],freqB[6]}),
    .clk(clk100m),
    .d({\PWMB/n0_lutinv ,\PWMB/n0_lutinv }),
    .sr(\PWMB/n11 ),
    .q({\PWMB/FreCnt [22],\PWMB/FreCnt [6]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMB/reg0_b24|PWMB/reg0_b4  (
    .b({\PWMB/n12 [24],\PWMB/n12 [4]}),
    .c({freqB[24],freqB[4]}),
    .clk(clk100m),
    .d({\PWMB/n0_lutinv ,\PWMB/n0_lutinv }),
    .sr(\PWMB/n11 ),
    .q({\PWMB/FreCnt [24],\PWMB/FreCnt [4]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMB/reg0_b2|PWMB/reg0_b26  (
    .b({\PWMB/n12 [2],\PWMB/n12 [26]}),
    .c({freqB[2],freqB[26]}),
    .clk(clk100m),
    .d({\PWMB/n0_lutinv ,\PWMB/n0_lutinv }),
    .sr(\PWMB/n11 ),
    .q({\PWMB/FreCnt [2],\PWMB/FreCnt [26]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(~A*~(~D*C)*~(0@B))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(~A*~(~D*C)*~(1@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b0001000100000001),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b0100010000000100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg1_b10|PWMB/reg1_b17  (
    .a({_al_u2656_o,_al_u1553_o}),
    .b({\PWMB/FreCnt [16],\PWMB/FreCnt [17]}),
    .c(\PWMB/FreCnt [9:8]),
    .ce(\PWMB/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMB/FreCntr [10],\PWMB/FreCntr [17]}),
    .e({\PWMB/FreCntr [17],\PWMB/FreCntr [8]}),
    .mi({freqB[10],freqB[17]}),
    .f({_al_u2657_o,_al_u1554_o}),
    .q({\PWMB/FreCntr [10],\PWMB/FreCntr [17]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*~C)*~(D*~B))"),
    //.LUTF1("(A*~(~0*C)*~(D*~B))"),
    //.LUTG0("(A*~(1*~C)*~(D*~B))"),
    //.LUTG1("(A*~(~1*C)*~(D*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000100010101010),
    .INIT_LUTF1(16'b0000100000001010),
    .INIT_LUTG0(16'b1000000010100000),
    .INIT_LUTG1(16'b1000100010101010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg1_b11|PWMB/reg1_b4  (
    .a({_al_u2638_o,_al_u2634_o}),
    .b({\PWMB/FreCnt [10],\PWMB/FreCnt [17]}),
    .c({\PWMB/FreCnt [3],\PWMB/FreCnt [3]}),
    .ce(\PWMB/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMB/FreCntr [11],\PWMB/FreCntr [18]}),
    .e({\PWMB/FreCntr [4],\PWMB/FreCntr [4]}),
    .mi({freqB[11],freqB[4]}),
    .f({_al_u2639_o,_al_u2635_o}),
    .q({\PWMB/FreCntr [11],\PWMB/FreCntr [4]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~C*~(0@B)*~(~D*A))"),
    //.LUTF1("(~A*~(0@C)*~(D*~B))"),
    //.LUTG0("(~C*~(1@B)*~(~D*A))"),
    //.LUTG1("(~A*~(1@C)*~(D*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001100000001),
    .INIT_LUTF1(16'b0000010000000101),
    .INIT_LUTG0(16'b0000110000000100),
    .INIT_LUTG1(16'b0100000001010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg1_b12|PWMB/reg1_b3  (
    .a({_al_u2648_o,\PWMB/FreCnt [11]}),
    .b({\PWMB/FreCnt [11],\PWMB/FreCnt [2]}),
    .c({\PWMB/FreCnt [18],\PWMB/FreCnt [26]}),
    .ce(\PWMB/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMB/FreCntr [12],\PWMB/FreCntr [12]}),
    .e({\PWMB/FreCntr [19],\PWMB/FreCntr [3]}),
    .mi({freqB[12],freqB[3]}),
    .f({_al_u2649_o,_al_u2642_o}),
    .q({\PWMB/FreCntr [12],\PWMB/FreCntr [3]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(C*B*A*~(0@D))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(C*B*A*~(1@D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg1_b13|PWMB/reg1_b19  (
    .a({_al_u2637_o,_al_u1559_o}),
    .b({_al_u2639_o,\PWMB/FreCnt [13]}),
    .c({_al_u2640_o,\PWMB/FreCnt [19]}),
    .ce(\PWMB/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMB/FreCnt [12],\PWMB/FreCntr [13]}),
    .e({\PWMB/FreCntr [13],\PWMB/FreCntr [19]}),
    .mi({freqB[13],freqB[19]}),
    .f({_al_u2641_o,_al_u1560_o}),
    .q({\PWMB/FreCntr [13],\PWMB/FreCntr [19]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~A*~(~0*C)*~(D@B))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(~A*~(~1*C)*~(D@B))"),
    //.LUTG1("(C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010000000001),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0100010000010001),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg1_b16|PWMB/reg1_b14  (
    .a({open_n18596,_al_u2651_o}),
    .b({open_n18597,\PWMB/FreCnt [13]}),
    .c({\PWMB/FreCntr [16],\PWMB/FreCnt [15]}),
    .ce(\PWMB/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMB/FreCnt [15],\PWMB/FreCntr [14]}),
    .e({open_n18598,\PWMB/FreCntr [16]}),
    .mi({freqB[16],freqB[14]}),
    .f({_al_u2656_o,_al_u2652_o}),
    .q({\PWMB/FreCntr [16],\PWMB/FreCntr [14]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(D*~(C@B))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(D*~(C@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1100001100000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1100001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg1_b1|PWMB/reg1_b0  (
    .b({\PWMB/FreCnt [0],open_n18617}),
    .c({\PWMB/FreCntr [1],\PWMB/n11 }),
    .ce(\PWMB/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({_al_u2644_o,\PWMB/n0_lutinv }),
    .mi(freqB[1:0]),
    .f({_al_u2645_o,\PWMB/mux3_b0_sel_is_3_o }),
    .q(\PWMB/FreCntr [1:0]));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~D*B)*~(C*~A))"),
    //.LUT1("(~C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111100100011),
    .INIT_LUT1(16'b0000111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg1_b20|PWMB/reg1_b9  (
    .a({open_n18636,\PWMB/FreCnt [19]}),
    .b({open_n18637,\PWMB/FreCnt [8]}),
    .c({\PWMB/FreCntr [20],\PWMB/FreCntr [20]}),
    .ce(\PWMB/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMB/FreCnt [19],\PWMB/FreCntr [9]}),
    .mi({freqB[20],freqB[9]}),
    .f({_al_u2648_o,_al_u2634_o}),
    .q({\PWMB/FreCntr [20],\PWMB/FreCntr [9]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(C*~B)*~(~D*A))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(~(C*~B)*~(~D*A))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100111101000101),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1100111101000101),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg1_b21|PWMB/reg1_b24  (
    .a({\PWMB/FreCnt [20],\PWMB/FreCnt [23]}),
    .b({\PWMB/FreCnt [6],\PWMB/FreCnt [9]}),
    .c({\PWMB/FreCntr [21],\PWMB/FreCntr [10]}),
    .ce(\PWMB/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMB/FreCntr [7],\PWMB/FreCntr [24]}),
    .mi({freqB[21],freqB[24]}),
    .f({_al_u2644_o,_al_u2654_o}),
    .q({\PWMB/FreCntr [21],\PWMB/FreCntr [24]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg1_b23|PWMB/reg1_b15  (
    .a({\PWMB/FreCnt [22],_al_u2652_o}),
    .b({\PWMB/FreCnt [23],\PWMB/FreCnt [14]}),
    .c({\PWMB/FreCntr [22],\PWMB/FreCnt [22]}),
    .ce(\PWMB/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMB/FreCntr [23],\PWMB/FreCntr [15]}),
    .e({open_n18670,\PWMB/FreCntr [23]}),
    .mi({freqB[23],freqB[15]}),
    .f({_al_u1553_o,_al_u2653_o}),
    .q({\PWMB/FreCntr [23],\PWMB/FreCntr [15]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(A*~(0@C)*~(D@B))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(A*~(1@C)*~(D@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b0000100000000010),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000000000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg1_b25|PWMB/reg1_b5  (
    .a({_al_u2642_o,_al_u1551_o}),
    .b({\PWMB/FreCnt [24],\PWMB/FreCnt [18]}),
    .c({\PWMB/FreCnt [4],\PWMB/FreCnt [5]}),
    .ce(\PWMB/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMB/FreCntr [25],\PWMB/FreCntr [18]}),
    .e({\PWMB/FreCntr [5],\PWMB/FreCntr [5]}),
    .mi({freqB[25],freqB[5]}),
    .f({_al_u2643_o,_al_u1552_o}),
    .q({\PWMB/FreCntr [25],\PWMB/FreCntr [5]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(~0*C)*~(~D*B))"),
    //.LUTF1("(~(~D*B)*~(C*~A))"),
    //.LUTG0("(A*~(~1*C)*~(~D*B))"),
    //.LUTG1("(~(~D*B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101000000010),
    .INIT_LUTF1(16'b1010111100100011),
    .INIT_LUTG0(16'b1010101000100010),
    .INIT_LUTG1(16'b1010111100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg1_b26|PWMB/reg1_b18  (
    .a({\PWMB/FreCnt [25],_al_u2646_o}),
    .b({\PWMB/FreCnt [7],\PWMB/FreCnt [17]}),
    .c({\PWMB/FreCntr [26],\PWMB/FreCnt [25]}),
    .ce(\PWMB/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMB/FreCntr [8],\PWMB/FreCntr [18]}),
    .e({open_n18703,\PWMB/FreCntr [26]}),
    .mi({freqB[26],freqB[18]}),
    .f({_al_u2638_o,_al_u2647_o}),
    .q({\PWMB/FreCntr [26],\PWMB/FreCntr [18]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(~0*C)*~(D*~B))"),
    //.LUTF1("(~(D*~B)*~(~C*A))"),
    //.LUTG0("(A*~(~1*C)*~(D*~B))"),
    //.LUTG1("(~(D*~B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000001010),
    .INIT_LUTF1(16'b1100010011110101),
    .INIT_LUTG0(16'b1000100010101010),
    .INIT_LUTG1(16'b1100010011110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg1_b6|PWMB/reg1_b2  (
    .a({\PWMB/FreCnt [21],_al_u2654_o}),
    .b({\PWMB/FreCnt [5],\PWMB/FreCnt [1]}),
    .c({\PWMB/FreCntr [22],\PWMB/FreCnt [5]}),
    .ce(\PWMB/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMB/FreCntr [6],\PWMB/FreCntr [2]}),
    .e({open_n18720,\PWMB/FreCntr [6]}),
    .mi({freqB[6],freqB[2]}),
    .f({_al_u2636_o,_al_u2655_o}),
    .q({\PWMB/FreCntr [6],\PWMB/FreCntr [2]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(D*~B)*~(C*~A))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(~(D*~B)*~(C*~A))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000110010101111),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000110010101111),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg1_b7|PWMB/reg1_b8  (
    .a({\PWMB/FreCnt [7],\PWMB/FreCnt [7]}),
    .b(\PWMB/FreCnt [9:8]),
    .c({\PWMB/FreCntr [7],\PWMB/FreCntr [8]}),
    .ce(\PWMB/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMB/FreCntr [9],\PWMB/FreCntr [9]}),
    .mi({freqB[7],freqB[8]}),
    .f({_al_u1563_o,_al_u2646_o}),
    .q({\PWMB/FreCntr [7],\PWMB/FreCntr [8]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg2_b0|PWMB/reg3_b0  (
    .a({\PWMB/pnumr [0],_al_u2632_o}),
    .b({pnumB[0],\PWMB/n24 }),
    .c({pnumB[32],pnumcntB[0]}),
    .clk(clk100m),
    .d({pwm_start_stop[27],\PWMB/pnumr [0]}),
    .e({open_n18756,pwm_start_stop[27]}),
    .q({\PWMB/pnumr[0]_keep ,\PWMB/RemaTxNum[0]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011100010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011100010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg2_b10|PWMB/reg2_b8  (
    .a({\PWMB/pnumr [10],\PWMB/pnumr [8]}),
    .b({pnumB[10],pnumB[32]}),
    .c({pnumB[32],pnumB[8]}),
    .clk(clk100m),
    .d({pwm_start_stop[27],pwm_start_stop[27]}),
    .q({\PWMB/pnumr[10]_keep ,\PWMB/pnumr[8]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg2_b11|PWMB/reg3_b11  (
    .a({\PWMB/pnumr [11],_al_u2626_o}),
    .b({pnumB[11],\PWMB/n24 }),
    .c({pnumB[32],pnumcntB[11]}),
    .clk(clk100m),
    .d({pwm_start_stop[27],\PWMB/pnumr [11]}),
    .e({open_n18801,pwm_start_stop[27]}),
    .q({\PWMB/pnumr[11]_keep ,\PWMB/RemaTxNum[11]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg2_b12|PWMB/reg3_b12  (
    .a({\PWMB/pnumr [12],_al_u2624_o}),
    .b({pnumB[12],\PWMB/n24 }),
    .c({pnumB[32],pnumcntB[12]}),
    .clk(clk100m),
    .d({pwm_start_stop[27],\PWMB/pnumr [12]}),
    .e({open_n18823,pwm_start_stop[27]}),
    .q({\PWMB/pnumr[12]_keep ,\PWMB/RemaTxNum[12]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011100010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011100010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg2_b13|PWMB/reg2_b7  (
    .a({\PWMB/pnumr [13],\PWMB/pnumr [7]}),
    .b({pnumB[13],pnumB[32]}),
    .c({pnumB[32],pnumB[7]}),
    .clk(clk100m),
    .d({pwm_start_stop[27],pwm_start_stop[27]}),
    .q({\PWMB/pnumr[13]_keep ,\PWMB/pnumr[7]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011100010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg2_b14|PWMB/reg2_b4  (
    .a({\PWMB/pnumr [14],\PWMB/pnumr [4]}),
    .b({pnumB[14],pnumB[32]}),
    .c({pnumB[32],pnumB[4]}),
    .clk(clk100m),
    .d({pwm_start_stop[27],pwm_start_stop[27]}),
    .q({\PWMB/pnumr[14]_keep ,\PWMB/pnumr[4]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg2_b15|PWMB/reg3_b15  (
    .a({\PWMB/pnumr [15],_al_u2618_o}),
    .b({pnumB[15],\PWMB/n24 }),
    .c({pnumB[32],pnumcntB[15]}),
    .clk(clk100m),
    .d({pwm_start_stop[27],\PWMB/pnumr [15]}),
    .e({open_n18887,pwm_start_stop[27]}),
    .q({\PWMB/pnumr[15]_keep ,\PWMB/RemaTxNum[15]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg2_b16|PWMB/reg3_b16  (
    .a({\PWMB/pnumr [16],_al_u2616_o}),
    .b({pnumB[16],\PWMB/n24 }),
    .c({pnumB[32],pnumcntB[16]}),
    .clk(clk100m),
    .d({pwm_start_stop[27],\PWMB/pnumr [16]}),
    .e({open_n18909,pwm_start_stop[27]}),
    .q({\PWMB/pnumr[16]_keep ,\PWMB/RemaTxNum[16]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg2_b17|PWMB/reg2_b3  (
    .a({\PWMB/pnumr [17],\PWMB/pnumr [3]}),
    .b({pnumB[17],pnumB[3]}),
    .c({pnumB[32],pnumB[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[27],pwm_start_stop[27]}),
    .q({\PWMB/pnumr[17]_keep ,\PWMB/pnumr[3]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg2_b18|PWMB/reg2_b21  (
    .a({\PWMB/pnumr [18],\PWMB/pnumr [21]}),
    .b({pnumB[18],pnumB[21]}),
    .c({pnumB[32],pnumB[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[27],pwm_start_stop[27]}),
    .q({\PWMB/pnumr[18]_keep ,\PWMB/pnumr[21]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg2_b19|PWMB/reg3_b19  (
    .a({\PWMB/pnumr [19],_al_u2610_o}),
    .b({pnumB[19],\PWMB/n24 }),
    .c({pnumB[32],pnumcntB[19]}),
    .clk(clk100m),
    .d({pwm_start_stop[27],\PWMB/pnumr [19]}),
    .e({open_n18973,pwm_start_stop[27]}),
    .q({\PWMB/pnumr[19]_keep ,\PWMB/RemaTxNum[19]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg2_b1|PWMB/reg2_b20  (
    .a({\PWMB/pnumr [1],\PWMB/pnumr [20]}),
    .b({pnumB[1],pnumB[20]}),
    .c({pnumB[32],pnumB[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[27],pwm_start_stop[27]}),
    .q({\PWMB/pnumr[1]_keep ,\PWMB/pnumr[20]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg2_b22|PWMB/reg3_b22  (
    .a({\PWMB/pnumr [22],_al_u2602_o}),
    .b({pnumB[22],\PWMB/n24 }),
    .c({pnumB[32],pnumcntB[22]}),
    .clk(clk100m),
    .d({pwm_start_stop[27],\PWMB/pnumr [22]}),
    .e({open_n19018,pwm_start_stop[27]}),
    .q({\PWMB/pnumr[22]_keep ,\PWMB/RemaTxNum[22]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg2_b23|PWMB/reg3_b23  (
    .a({\PWMB/pnumr [23],_al_u2600_o}),
    .b({pnumB[23],\PWMB/n24 }),
    .c({pnumB[32],pnumcntB[23]}),
    .clk(clk100m),
    .d({pwm_start_stop[27],\PWMB/pnumr [23]}),
    .e({open_n19040,pwm_start_stop[27]}),
    .q({\PWMB/pnumr[23]_keep ,\PWMB/RemaTxNum[23]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg2_b24|PWMB/reg2_b31  (
    .a({\PWMB/pnumr [24],\PWMB/pnumr [31]}),
    .b({pnumB[24],pnumB[31]}),
    .c({pnumB[32],pnumB[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[27],pwm_start_stop[27]}),
    .q({\PWMB/pnumr[24]_keep ,\PWMB/pnumr[31]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg2_b25|PWMB/reg2_b30  (
    .a({\PWMB/pnumr [25],\PWMB/pnumr [30]}),
    .b({pnumB[25],pnumB[30]}),
    .c({pnumB[32],pnumB[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[27],pwm_start_stop[27]}),
    .q({\PWMB/pnumr[25]_keep ,\PWMB/pnumr[30]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg2_b26|PWMB/reg2_b29  (
    .a({\PWMB/pnumr [26],\PWMB/pnumr [29]}),
    .b({pnumB[26],pnumB[29]}),
    .c({pnumB[32],pnumB[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[27],pwm_start_stop[27]}),
    .q({\PWMB/pnumr[26]_keep ,\PWMB/pnumr[29]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg2_b27|PWMB/reg2_b28  (
    .a({\PWMB/pnumr [27],\PWMB/pnumr [28]}),
    .b({pnumB[27],pnumB[28]}),
    .c({pnumB[32],pnumB[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[27],pwm_start_stop[27]}),
    .q({\PWMB/pnumr[27]_keep ,\PWMB/pnumr[28]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg2_b2|PWMB/reg3_b2  (
    .a({\PWMB/pnumr [2],_al_u2608_o}),
    .b({pnumB[2],\PWMB/n24 }),
    .c({pnumB[32],pnumcntB[2]}),
    .clk(clk100m),
    .d({pwm_start_stop[27],\PWMB/pnumr [2]}),
    .e({open_n19142,pwm_start_stop[27]}),
    .q({\PWMB/pnumr[2]_keep ,\PWMB/RemaTxNum[2]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg2_b5|PWMB/reg3_b5  (
    .a({\PWMB/pnumr [5],_al_u2594_o}),
    .b({pnumB[32],\PWMB/n24 }),
    .c({pnumB[5],pnumcntB[5]}),
    .clk(clk100m),
    .d({pwm_start_stop[27],\PWMB/pnumr [5]}),
    .e({open_n19164,pwm_start_stop[27]}),
    .q({\PWMB/pnumr[5]_keep ,\PWMB/RemaTxNum[5]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg2_b6|PWMB/reg3_b6  (
    .a({\PWMB/pnumr [6],_al_u2592_o}),
    .b({pnumB[32],\PWMB/n24 }),
    .c({pnumB[6],pnumcntB[6]}),
    .clk(clk100m),
    .d({pwm_start_stop[27],\PWMB/pnumr [6]}),
    .e({open_n19186,pwm_start_stop[27]}),
    .q({\PWMB/pnumr[6]_keep ,\PWMB/RemaTxNum[6]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg2_b9|PWMB/reg3_b9  (
    .a({\PWMB/pnumr [9],_al_u2586_o}),
    .b({pnumB[32],\PWMB/n24 }),
    .c({pnumB[9],pnumcntB[9]}),
    .clk(clk100m),
    .d({pwm_start_stop[27],\PWMB/pnumr [9]}),
    .e({open_n19208,pwm_start_stop[27]}),
    .q({\PWMB/pnumr[9]_keep ,\PWMB/RemaTxNum[9]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg3_b1  (
    .a({_al_u2630_o,_al_u2630_o}),
    .b({\PWMB/n24 ,\PWMB/n24 }),
    .c({pnumcntB[1],pnumcntB[1]}),
    .clk(clk100m),
    .d({\PWMB/pnumr [1],\PWMB/pnumr [1]}),
    .mi({open_n19240,pwm_start_stop[27]}),
    .q({open_n19247,\PWMB/RemaTxNum[1]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg3_b10  (
    .a({_al_u2628_o,_al_u2628_o}),
    .b({\PWMB/n24 ,\PWMB/n24 }),
    .c({pnumcntB[10],pnumcntB[10]}),
    .clk(clk100m),
    .d({\PWMB/pnumr [10],\PWMB/pnumr [10]}),
    .mi({open_n19259,pwm_start_stop[27]}),
    .q({open_n19266,\PWMB/RemaTxNum[10]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg3_b13  (
    .a({_al_u2622_o,_al_u2622_o}),
    .b({\PWMB/n24 ,\PWMB/n24 }),
    .c({pnumcntB[13],pnumcntB[13]}),
    .clk(clk100m),
    .d({\PWMB/pnumr [13],\PWMB/pnumr [13]}),
    .mi({open_n19278,pwm_start_stop[27]}),
    .q({open_n19285,\PWMB/RemaTxNum[13]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg3_b14  (
    .a({_al_u2620_o,_al_u2620_o}),
    .b({\PWMB/n24 ,\PWMB/n24 }),
    .c({pnumcntB[14],pnumcntB[14]}),
    .clk(clk100m),
    .d({\PWMB/pnumr [14],\PWMB/pnumr [14]}),
    .mi({open_n19297,pwm_start_stop[27]}),
    .q({open_n19304,\PWMB/RemaTxNum[14]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg3_b17  (
    .a({_al_u2614_o,_al_u2614_o}),
    .b({\PWMB/n24 ,\PWMB/n24 }),
    .c({pnumcntB[17],pnumcntB[17]}),
    .clk(clk100m),
    .d({\PWMB/pnumr [17],\PWMB/pnumr [17]}),
    .mi({open_n19316,pwm_start_stop[27]}),
    .q({open_n19323,\PWMB/RemaTxNum[17]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg3_b18  (
    .a({_al_u2612_o,_al_u2612_o}),
    .b({\PWMB/n24 ,\PWMB/n24 }),
    .c({pnumcntB[18],pnumcntB[18]}),
    .clk(clk100m),
    .d({\PWMB/pnumr [18],\PWMB/pnumr [18]}),
    .mi({open_n19335,pwm_start_stop[27]}),
    .q({open_n19342,\PWMB/RemaTxNum[18]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg3_b20  (
    .a({_al_u2606_o,_al_u2606_o}),
    .b({\PWMB/n24 ,\PWMB/n24 }),
    .c({pnumcntB[20],pnumcntB[20]}),
    .clk(clk100m),
    .d({\PWMB/pnumr [20],\PWMB/pnumr [20]}),
    .mi({open_n19354,pwm_start_stop[27]}),
    .q({open_n19361,\PWMB/RemaTxNum[20]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg3_b21  (
    .a({_al_u2604_o,_al_u2604_o}),
    .b({\PWMB/n24 ,\PWMB/n24 }),
    .c({pnumcntB[21],pnumcntB[21]}),
    .clk(clk100m),
    .d({\PWMB/pnumr [21],\PWMB/pnumr [21]}),
    .mi({open_n19373,pwm_start_stop[27]}),
    .q({open_n19380,\PWMB/RemaTxNum[21]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg3_b3  (
    .a({_al_u2598_o,_al_u2598_o}),
    .b({\PWMB/n24 ,\PWMB/n24 }),
    .c({pnumcntB[3],pnumcntB[3]}),
    .clk(clk100m),
    .d({\PWMB/pnumr [3],\PWMB/pnumr [3]}),
    .mi({open_n19392,pwm_start_stop[27]}),
    .q({open_n19399,\PWMB/RemaTxNum[3]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg3_b4  (
    .a({_al_u2596_o,_al_u2596_o}),
    .b({\PWMB/n24 ,\PWMB/n24 }),
    .c({pnumcntB[4],pnumcntB[4]}),
    .clk(clk100m),
    .d({\PWMB/pnumr [4],\PWMB/pnumr [4]}),
    .mi({open_n19411,pwm_start_stop[27]}),
    .q({open_n19418,\PWMB/RemaTxNum[4]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg3_b7  (
    .a({_al_u2590_o,_al_u2590_o}),
    .b({\PWMB/n24 ,\PWMB/n24 }),
    .c({pnumcntB[7],pnumcntB[7]}),
    .clk(clk100m),
    .d({\PWMB/pnumr [7],\PWMB/pnumr [7]}),
    .mi({open_n19430,pwm_start_stop[27]}),
    .q({open_n19437,\PWMB/RemaTxNum[7]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/reg3_b8  (
    .a({_al_u2588_o,_al_u2588_o}),
    .b({\PWMB/n24 ,\PWMB/n24 }),
    .c({pnumcntB[8],pnumcntB[8]}),
    .clk(clk100m),
    .d({\PWMB/pnumr [8],\PWMB/pnumr [8]}),
    .mi({open_n19449,pwm_start_stop[27]}),
    .q({open_n19456,\PWMB/RemaTxNum[8]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_LSLICE #(
    //.MACRO("PWMB/sub0/ucin_al_u3440"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWMB/sub0/u11_al_u3443  (
    .a({\PWMB/FreCnt [13],\PWMB/FreCnt [11]}),
    .b({\PWMB/FreCnt [14],\PWMB/FreCnt [12]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWMB/sub0/c11 ),
    .f({\PWMB/n12 [13],\PWMB/n12 [11]}),
    .fco(\PWMB/sub0/c15 ),
    .fx({\PWMB/n12 [14],\PWMB/n12 [12]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWMB/sub0/ucin_al_u3440"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWMB/sub0/u15_al_u3444  (
    .a({\PWMB/FreCnt [17],\PWMB/FreCnt [15]}),
    .b({\PWMB/FreCnt [18],\PWMB/FreCnt [16]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWMB/sub0/c15 ),
    .f({\PWMB/n12 [17],\PWMB/n12 [15]}),
    .fco(\PWMB/sub0/c19 ),
    .fx({\PWMB/n12 [18],\PWMB/n12 [16]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWMB/sub0/ucin_al_u3440"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWMB/sub0/u19_al_u3445  (
    .a({\PWMB/FreCnt [21],\PWMB/FreCnt [19]}),
    .b({\PWMB/FreCnt [22],\PWMB/FreCnt [20]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWMB/sub0/c19 ),
    .f({\PWMB/n12 [21],\PWMB/n12 [19]}),
    .fco(\PWMB/sub0/c23 ),
    .fx({\PWMB/n12 [22],\PWMB/n12 [20]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWMB/sub0/ucin_al_u3440"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWMB/sub0/u23_al_u3446  (
    .a({\PWMB/FreCnt [25],\PWMB/FreCnt [23]}),
    .b({\PWMB/FreCnt [26],\PWMB/FreCnt [24]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWMB/sub0/c23 ),
    .f({\PWMB/n12 [25],\PWMB/n12 [23]}),
    .fx({\PWMB/n12 [26],\PWMB/n12 [24]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWMB/sub0/ucin_al_u3440"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWMB/sub0/u3_al_u3441  (
    .a({\PWMB/FreCnt [5],\PWMB/FreCnt [3]}),
    .b({\PWMB/FreCnt [6],\PWMB/FreCnt [4]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWMB/sub0/c3 ),
    .f({\PWMB/n12 [5],\PWMB/n12 [3]}),
    .fco(\PWMB/sub0/c7 ),
    .fx({\PWMB/n12 [6],\PWMB/n12 [4]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWMB/sub0/ucin_al_u3440"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWMB/sub0/u7_al_u3442  (
    .a({\PWMB/FreCnt [9],\PWMB/FreCnt [7]}),
    .b({\PWMB/FreCnt [10],\PWMB/FreCnt [8]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWMB/sub0/c7 ),
    .f({\PWMB/n12 [9],\PWMB/n12 [7]}),
    .fco(\PWMB/sub0/c11 ),
    .fx({\PWMB/n12 [10],\PWMB/n12 [8]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWMB/sub0/ucin_al_u3440"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h0005),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWMB/sub0/ucin_al_u3440  (
    .a({\PWMB/FreCnt [1],1'b0}),
    .b({\PWMB/FreCnt [2],\PWMB/FreCnt [0]}),
    .c(2'b11),
    .d(2'b01),
    .e(2'b01),
    .f({\PWMB/n12 [1],open_n19583}),
    .fco(\PWMB/sub0/c3 ),
    .fx({\PWMB/n12 [2],\PWMB/n12 [0]}));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMB/sub1/u0|PWMB/sub1/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("SUB_CARRY"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000101),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMB/sub1/u0|PWMB/sub1/ucin  (
    .a({pnumcntB[0],1'b0}),
    .b({1'b1,open_n19586}),
    .ce(\U_AHB/n8 ),
    .clk(clk100m),
    .mi(\U_AHB/h2h_hwdata [26:25]),
    .f({\PWMB/n26 [0],open_n19602}),
    .fco(\PWMB/sub1/c1 ),
    .q(freq2[26:25]));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMB/sub1/u0|PWMB/sub1/ucin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMB/sub1/u10|PWMB/sub1/u9  (
    .a(pnumcntB[10:9]),
    .b(2'b00),
    .fci(\PWMB/sub1/c9 ),
    .f(\PWMB/n26 [10:9]),
    .fco(\PWMB/sub1/c11 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMB/sub1/u0|PWMB/sub1/ucin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMB/sub1/u12|PWMB/sub1/u11  (
    .a(pnumcntB[12:11]),
    .b(2'b00),
    .fci(\PWMB/sub1/c11 ),
    .f(\PWMB/n26 [12:11]),
    .fco(\PWMB/sub1/c13 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMB/sub1/u0|PWMB/sub1/ucin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMB/sub1/u14|PWMB/sub1/u13  (
    .a(pnumcntB[14:13]),
    .b(2'b00),
    .fci(\PWMB/sub1/c13 ),
    .f(\PWMB/n26 [14:13]),
    .fco(\PWMB/sub1/c15 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMB/sub1/u0|PWMB/sub1/ucin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMB/sub1/u16|PWMB/sub1/u15  (
    .a(pnumcntB[16:15]),
    .b(2'b00),
    .fci(\PWMB/sub1/c15 ),
    .f(\PWMB/n26 [16:15]),
    .fco(\PWMB/sub1/c17 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMB/sub1/u0|PWMB/sub1/ucin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMB/sub1/u18|PWMB/sub1/u17  (
    .a(pnumcntB[18:17]),
    .b(2'b00),
    .fci(\PWMB/sub1/c17 ),
    .f(\PWMB/n26 [18:17]),
    .fco(\PWMB/sub1/c19 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMB/sub1/u0|PWMB/sub1/ucin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMB/sub1/u20|PWMB/sub1/u19  (
    .a(pnumcntB[20:19]),
    .b(2'b00),
    .fci(\PWMB/sub1/c19 ),
    .f(\PWMB/n26 [20:19]),
    .fco(\PWMB/sub1/c21 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMB/sub1/u0|PWMB/sub1/ucin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMB/sub1/u22|PWMB/sub1/u21  (
    .a(pnumcntB[22:21]),
    .b(2'b00),
    .fci(\PWMB/sub1/c21 ),
    .f(\PWMB/n26 [22:21]),
    .fco(\PWMB/sub1/c23 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMB/sub1/u0|PWMB/sub1/ucin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMB/sub1/u23_al_u3479  (
    .a({open_n19759,pnumcntB[23]}),
    .b({open_n19760,1'b0}),
    .fci(\PWMB/sub1/c23 ),
    .f({open_n19779,\PWMB/n26 [23]}));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMB/sub1/u0|PWMB/sub1/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMB/sub1/u2|PWMB/sub1/u1  (
    .a(pnumcntB[2:1]),
    .b(2'b00),
    .fci(\PWMB/sub1/c1 ),
    .f(\PWMB/n26 [2:1]),
    .fco(\PWMB/sub1/c3 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMB/sub1/u0|PWMB/sub1/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMB/sub1/u4|PWMB/sub1/u3  (
    .a(pnumcntB[4:3]),
    .b(2'b00),
    .fci(\PWMB/sub1/c3 ),
    .f(\PWMB/n26 [4:3]),
    .fco(\PWMB/sub1/c5 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMB/sub1/u0|PWMB/sub1/ucin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMB/sub1/u6|PWMB/sub1/u5  (
    .a(pnumcntB[6:5]),
    .b(2'b00),
    .fci(\PWMB/sub1/c5 ),
    .f(\PWMB/n26 [6:5]),
    .fco(\PWMB/sub1/c7 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMB/sub1/u0|PWMB/sub1/ucin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMB/sub1/u8|PWMB/sub1/u7  (
    .a(pnumcntB[8:7]),
    .b(2'b00),
    .fci(\PWMB/sub1/c7 ),
    .f(\PWMB/n26 [8:7]),
    .fco(\PWMB/sub1/c9 ));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[0]  (
    .i(\PWMC/RemaTxNum[0]_keep ),
    .o(pnumcntC[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[10]  (
    .i(\PWMC/RemaTxNum[10]_keep ),
    .o(pnumcntC[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[11]  (
    .i(\PWMC/RemaTxNum[11]_keep ),
    .o(pnumcntC[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[12]  (
    .i(\PWMC/RemaTxNum[12]_keep ),
    .o(pnumcntC[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[13]  (
    .i(\PWMC/RemaTxNum[13]_keep ),
    .o(pnumcntC[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[14]  (
    .i(\PWMC/RemaTxNum[14]_keep ),
    .o(pnumcntC[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[15]  (
    .i(\PWMC/RemaTxNum[15]_keep ),
    .o(pnumcntC[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[16]  (
    .i(\PWMC/RemaTxNum[16]_keep ),
    .o(pnumcntC[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[17]  (
    .i(\PWMC/RemaTxNum[17]_keep ),
    .o(pnumcntC[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[18]  (
    .i(\PWMC/RemaTxNum[18]_keep ),
    .o(pnumcntC[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[19]  (
    .i(\PWMC/RemaTxNum[19]_keep ),
    .o(pnumcntC[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[1]  (
    .i(\PWMC/RemaTxNum[1]_keep ),
    .o(pnumcntC[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[20]  (
    .i(\PWMC/RemaTxNum[20]_keep ),
    .o(pnumcntC[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[21]  (
    .i(\PWMC/RemaTxNum[21]_keep ),
    .o(pnumcntC[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[22]  (
    .i(\PWMC/RemaTxNum[22]_keep ),
    .o(pnumcntC[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[23]  (
    .i(\PWMC/RemaTxNum[23]_keep ),
    .o(pnumcntC[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[2]  (
    .i(\PWMC/RemaTxNum[2]_keep ),
    .o(pnumcntC[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[3]  (
    .i(\PWMC/RemaTxNum[3]_keep ),
    .o(pnumcntC[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[4]  (
    .i(\PWMC/RemaTxNum[4]_keep ),
    .o(pnumcntC[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[5]  (
    .i(\PWMC/RemaTxNum[5]_keep ),
    .o(pnumcntC[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[6]  (
    .i(\PWMC/RemaTxNum[6]_keep ),
    .o(pnumcntC[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[7]  (
    .i(\PWMC/RemaTxNum[7]_keep ),
    .o(pnumcntC[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[8]  (
    .i(\PWMC/RemaTxNum[8]_keep ),
    .o(pnumcntC[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[9]  (
    .i(\PWMC/RemaTxNum[9]_keep ),
    .o(pnumcntC[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_dir  (
    .i(\PWMC/dir_keep ),
    .o(dir_pad[12]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[0]  (
    .i(\PWMC/pnumr[0]_keep ),
    .o(\PWMC/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[10]  (
    .i(\PWMC/pnumr[10]_keep ),
    .o(\PWMC/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[11]  (
    .i(\PWMC/pnumr[11]_keep ),
    .o(\PWMC/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[12]  (
    .i(\PWMC/pnumr[12]_keep ),
    .o(\PWMC/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[13]  (
    .i(\PWMC/pnumr[13]_keep ),
    .o(\PWMC/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[14]  (
    .i(\PWMC/pnumr[14]_keep ),
    .o(\PWMC/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[15]  (
    .i(\PWMC/pnumr[15]_keep ),
    .o(\PWMC/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[16]  (
    .i(\PWMC/pnumr[16]_keep ),
    .o(\PWMC/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[17]  (
    .i(\PWMC/pnumr[17]_keep ),
    .o(\PWMC/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[18]  (
    .i(\PWMC/pnumr[18]_keep ),
    .o(\PWMC/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[19]  (
    .i(\PWMC/pnumr[19]_keep ),
    .o(\PWMC/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[1]  (
    .i(\PWMC/pnumr[1]_keep ),
    .o(\PWMC/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[20]  (
    .i(\PWMC/pnumr[20]_keep ),
    .o(\PWMC/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[21]  (
    .i(\PWMC/pnumr[21]_keep ),
    .o(\PWMC/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[22]  (
    .i(\PWMC/pnumr[22]_keep ),
    .o(\PWMC/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[23]  (
    .i(\PWMC/pnumr[23]_keep ),
    .o(\PWMC/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[24]  (
    .i(\PWMC/pnumr[24]_keep ),
    .o(\PWMC/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[25]  (
    .i(\PWMC/pnumr[25]_keep ),
    .o(\PWMC/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[26]  (
    .i(\PWMC/pnumr[26]_keep ),
    .o(\PWMC/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[27]  (
    .i(\PWMC/pnumr[27]_keep ),
    .o(\PWMC/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[28]  (
    .i(\PWMC/pnumr[28]_keep ),
    .o(\PWMC/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[29]  (
    .i(\PWMC/pnumr[29]_keep ),
    .o(\PWMC/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[2]  (
    .i(\PWMC/pnumr[2]_keep ),
    .o(\PWMC/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[30]  (
    .i(\PWMC/pnumr[30]_keep ),
    .o(\PWMC/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[31]  (
    .i(\PWMC/pnumr[31]_keep ),
    .o(\PWMC/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[3]  (
    .i(\PWMC/pnumr[3]_keep ),
    .o(\PWMC/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[4]  (
    .i(\PWMC/pnumr[4]_keep ),
    .o(\PWMC/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[5]  (
    .i(\PWMC/pnumr[5]_keep ),
    .o(\PWMC/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[6]  (
    .i(\PWMC/pnumr[6]_keep ),
    .o(\PWMC/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[7]  (
    .i(\PWMC/pnumr[7]_keep ),
    .o(\PWMC/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[8]  (
    .i(\PWMC/pnumr[8]_keep ),
    .o(\PWMC/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[9]  (
    .i(\PWMC/pnumr[9]_keep ),
    .o(\PWMC/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pwm  (
    .i(\PWMC/pwm_keep ),
    .o(pwm_pad[12]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_stopreq  (
    .i(\PWMC/stopreq_keep ),
    .o(\PWMC/stopreq ));  // src/OnePWM.v(14)
  EF2_PHY_MSLICE #(
    //.LUT0("(D*~(C)*~((~0*~(B*A)))+D*C*~((~0*~(B*A)))+~(D)*C*(~0*~(B*A))+D*C*(~0*~(B*A)))"),
    //.LUT1("(D*~(C)*~((~1*~(B*A)))+D*C*~((~1*~(B*A)))+~(D)*C*(~1*~(B*A))+D*C*(~1*~(B*A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111100001110000),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/dir_reg  (
    .a({\PWMC/n24 ,\PWMC/n24 }),
    .b({\PWMC/n25_neg_lutinv ,\PWMC/n25_neg_lutinv }),
    .c({dir_pad[12],dir_pad[12]}),
    .clk(clk100m),
    .d({\PWMC/pnumr [31],\PWMC/pnumr [31]}),
    .mi({open_n19884,pwm_start_stop[28]}),
    .q({open_n19891,\PWMC/dir_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("~(~0*~(D*C*B*A))"),
    //.LUT1("~(~1*~(D*C*B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b1111111111111111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMC/pwm_reg  (
    .a({_al_u1573_o,_al_u1573_o}),
    .b({_al_u1579_o,_al_u1579_o}),
    .c({_al_u1581_o,_al_u1581_o}),
    .clk(clk100m),
    .d({_al_u1583_o,_al_u1583_o}),
    .mi({open_n19903,pwm_pad[12]}),
    .sr(\PWMC/u14_sel_is_1_o ),
    .q({open_n19909,\PWMC/pwm_keep }));  // src/OnePWM.v(45)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMC/reg0_b0|PWMC/reg0_b21  (
    .b({\PWMC/n12 [0],\PWMC/n12 [21]}),
    .c({freqC[0],freqC[21]}),
    .clk(clk100m),
    .d({\PWMC/n0_lutinv ,\PWMC/n0_lutinv }),
    .sr(\PWMC/n11 ),
    .q({\PWMC/FreCnt [0],\PWMC/FreCnt [21]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMC/reg0_b10|PWMC/reg0_b15  (
    .b({\PWMC/n12 [10],\PWMC/n12 [15]}),
    .c({freqC[10],freqC[15]}),
    .clk(clk100m),
    .d({\PWMC/n0_lutinv ,\PWMC/n0_lutinv }),
    .sr(\PWMC/n11 ),
    .q({\PWMC/FreCnt [10],\PWMC/FreCnt [15]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMC/reg0_b11|PWMC/reg0_b7  (
    .b({\PWMC/n12 [11],\PWMC/n12 [7]}),
    .c({freqC[11],freqC[7]}),
    .clk(clk100m),
    .d({\PWMC/n0_lutinv ,\PWMC/n0_lutinv }),
    .sr(\PWMC/n11 ),
    .q({\PWMC/FreCnt [11],\PWMC/FreCnt [7]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMC/reg0_b12|PWMC/reg0_b5  (
    .b({\PWMC/n12 [12],\PWMC/n12 [5]}),
    .c({freqC[12],freqC[5]}),
    .clk(clk100m),
    .d({\PWMC/n0_lutinv ,\PWMC/n0_lutinv }),
    .sr(\PWMC/n11 ),
    .q({\PWMC/FreCnt [12],\PWMC/FreCnt [5]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMC/reg0_b13|PWMC/reg0_b3  (
    .b({\PWMC/n12 [13],\PWMC/n12 [3]}),
    .c({freqC[13],freqC[3]}),
    .clk(clk100m),
    .d({\PWMC/n0_lutinv ,\PWMC/n0_lutinv }),
    .sr(\PWMC/n11 ),
    .q({\PWMC/FreCnt [13],\PWMC/FreCnt [3]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMC/reg0_b14|PWMC/reg0_b25  (
    .b({\PWMC/n12 [14],\PWMC/n12 [25]}),
    .c({freqC[14],freqC[25]}),
    .clk(clk100m),
    .d({\PWMC/n0_lutinv ,\PWMC/n0_lutinv }),
    .sr(\PWMC/n11 ),
    .q({\PWMC/FreCnt [14],\PWMC/FreCnt [25]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMC/reg0_b16|PWMC/reg0_b23  (
    .b({\PWMC/n12 [16],\PWMC/n12 [23]}),
    .c({freqC[16],freqC[23]}),
    .clk(clk100m),
    .d({\PWMC/n0_lutinv ,\PWMC/n0_lutinv }),
    .sr(\PWMC/n11 ),
    .q({\PWMC/FreCnt [16],\PWMC/FreCnt [23]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMC/reg0_b17|PWMC/reg0_b19  (
    .b({\PWMC/n12 [17],\PWMC/n12 [19]}),
    .c({freqC[17],freqC[19]}),
    .clk(clk100m),
    .d({\PWMC/n0_lutinv ,\PWMC/n0_lutinv }),
    .sr(\PWMC/n11 ),
    .q({\PWMC/FreCnt [17],\PWMC/FreCnt [19]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMC/reg0_b18|PWMC/reg0_b9  (
    .b({\PWMC/n12 [18],\PWMC/n12 [9]}),
    .c({freqC[18],freqC[9]}),
    .clk(clk100m),
    .d({\PWMC/n0_lutinv ,\PWMC/n0_lutinv }),
    .sr(\PWMC/n11 ),
    .q({\PWMC/FreCnt [18],\PWMC/FreCnt [9]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMC/reg0_b1|PWMC/reg0_b8  (
    .b({\PWMC/n12 [1],\PWMC/n12 [8]}),
    .c({freqC[1],freqC[8]}),
    .clk(clk100m),
    .d({\PWMC/n0_lutinv ,\PWMC/n0_lutinv }),
    .sr(\PWMC/n11 ),
    .q({\PWMC/FreCnt [1],\PWMC/FreCnt [8]}));  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMC/reg0_b2  (
    .b({open_n20140,\PWMC/n12 [2]}),
    .c({open_n20141,freqC[2]}),
    .clk(clk100m),
    .d({open_n20143,\PWMC/n0_lutinv }),
    .sr(\PWMC/n11 ),
    .q({open_n20165,\PWMC/FreCnt [2]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMC/reg0_b20|PWMC/reg0_b6  (
    .b({\PWMC/n12 [20],\PWMC/n12 [6]}),
    .c({freqC[20],freqC[6]}),
    .clk(clk100m),
    .d({\PWMC/n0_lutinv ,\PWMC/n0_lutinv }),
    .sr(\PWMC/n11 ),
    .q({\PWMC/FreCnt [20],\PWMC/FreCnt [6]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMC/reg0_b22|PWMC/reg0_b4  (
    .b({\PWMC/n12 [22],\PWMC/n12 [4]}),
    .c({freqC[22],freqC[4]}),
    .clk(clk100m),
    .d({\PWMC/n0_lutinv ,\PWMC/n0_lutinv }),
    .sr(\PWMC/n11 ),
    .q({\PWMC/FreCnt [22],\PWMC/FreCnt [4]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMC/reg0_b24|PWMC/reg0_b26  (
    .b({\PWMC/n12 [24],\PWMC/n12 [26]}),
    .c({freqC[24],freqC[26]}),
    .clk(clk100m),
    .d({\PWMC/n0_lutinv ,\PWMC/n0_lutinv }),
    .sr(\PWMC/n11 ),
    .q({\PWMC/FreCnt [24],\PWMC/FreCnt [26]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(A*~(D@C)*~(0@B))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(A*~(D@C)*~(1@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b0010000000000010),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg1_b10|PWMC/reg1_b7  (
    .a({_al_u2734_o,_al_u1570_o}),
    .b({\PWMC/FreCnt [6],\PWMC/FreCnt [7]}),
    .c({\PWMC/FreCnt [9],\PWMC/FreCnt [9]}),
    .ce(\PWMC/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMC/FreCntr [10],\PWMC/FreCntr [7]}),
    .e({\PWMC/FreCntr [7],\PWMC/FreCntr [9]}),
    .mi({freqC[10],freqC[7]}),
    .f({_al_u2735_o,_al_u1571_o}),
    .q({\PWMC/FreCntr [10],\PWMC/FreCntr [7]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(D*~B)*~(~C*A))"),
    //.LUT1("(~(~D*B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100010011110101),
    .INIT_LUT1(16'b1010111100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg1_b11|PWMC/reg1_b18  (
    .a({\PWMC/FreCnt [10],\PWMC/FreCnt [17]}),
    .b({\PWMC/FreCnt [3],\PWMC/FreCnt [21]}),
    .c({\PWMC/FreCntr [11],\PWMC/FreCntr [18]}),
    .ce(\PWMC/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMC/FreCntr [4],\PWMC/FreCntr [22]}),
    .mi({freqC[11],freqC[18]}),
    .f({_al_u2728_o,_al_u2720_o}),
    .q({\PWMC/FreCntr [11],\PWMC/FreCntr [18]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(~0*C)*~(D*~B))"),
    //.LUTF1("(~C*~(~0*B)*~(D@A))"),
    //.LUTG0("(A*~(~1*C)*~(D*~B))"),
    //.LUTG1("(~C*~(~1*B)*~(D@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000001010),
    .INIT_LUTF1(16'b0000001000000001),
    .INIT_LUTG0(16'b1000100010101010),
    .INIT_LUTG1(16'b0000101000000101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg1_b12|PWMC/reg1_b17  (
    .a({\PWMC/FreCnt [11],_al_u2728_o}),
    .b({\PWMC/FreCnt [16],\PWMC/FreCnt [16]}),
    .c({\PWMC/FreCnt [26],\PWMC/FreCnt [7]}),
    .ce(\PWMC/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMC/FreCntr [12],\PWMC/FreCntr [17]}),
    .e({\PWMC/FreCntr [17],\PWMC/FreCntr [8]}),
    .mi({freqC[12],freqC[17]}),
    .f({_al_u2730_o,_al_u2729_o}),
    .q({\PWMC/FreCntr [12],\PWMC/FreCntr [17]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(D@B)*~(C@A))"),
    //.LUTF1("(D*~(C@B))"),
    //.LUTG0("(~(D@B)*~(C@A))"),
    //.LUTG1("(D*~(C@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000010000100001),
    .INIT_LUTF1(16'b1100001100000000),
    .INIT_LUTG0(16'b1000010000100001),
    .INIT_LUTG1(16'b1100001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg1_b14|PWMC/reg1_b4  (
    .a({open_n20276,\PWMC/FreCnt [16]}),
    .b({\PWMC/FreCnt [13],\PWMC/FreCnt [4]}),
    .c({\PWMC/FreCntr [14],\PWMC/FreCntr [16]}),
    .ce(\PWMC/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({_al_u2724_o,\PWMC/FreCntr [4]}),
    .mi({freqC[14],freqC[4]}),
    .f({_al_u2725_o,_al_u1568_o}),
    .q({\PWMC/FreCntr [14],\PWMC/FreCntr [4]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg1_b15|PWMC/reg1_b5  (
    .a({\PWMC/FreCnt [14],_al_u1568_o}),
    .b({\PWMC/FreCnt [4],\PWMC/FreCnt [18]}),
    .c({\PWMC/FreCntr [15],\PWMC/FreCnt [5]}),
    .ce(\PWMC/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMC/FreCntr [5],\PWMC/FreCntr [18]}),
    .e({open_n20295,\PWMC/FreCntr [5]}),
    .mi({freqC[15],freqC[5]}),
    .f({_al_u2724_o,_al_u1569_o}),
    .q({\PWMC/FreCntr [15],\PWMC/FreCntr [5]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*B*A*~(0@D))"),
    //.LUTF1("(~(D*~B)*~(~C*A))"),
    //.LUTG0("(C*B*A*~(1@D))"),
    //.LUTG1("(~(D*~B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b1100010011110101),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b1100010011110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg1_b16|PWMC/reg1_b25  (
    .a({\PWMC/FreCnt [15],_al_u2719_o}),
    .b({\PWMC/FreCnt [17],_al_u2721_o}),
    .c({\PWMC/FreCntr [16],_al_u2722_o}),
    .ce(\PWMC/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMC/FreCntr [18],\PWMC/FreCnt [24]}),
    .e({open_n20312,\PWMC/FreCntr [25]}),
    .mi({freqC[16],freqC[25]}),
    .f({_al_u2722_o,_al_u2723_o}),
    .q({\PWMC/FreCntr [16],\PWMC/FreCntr [25]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1000010000100001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg1_b1|PWMC/reg1_b9  (
    .a({\PWMC/FreCnt [0],open_n20329}),
    .b({\PWMC/FreCnt [8],open_n20330}),
    .c({\PWMC/FreCntr [1],pwm_state_read[12]}),
    .ce(\PWMC/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMC/FreCntr [9],\PWMC/n0_lutinv }),
    .mi({freqC[1],freqC[9]}),
    .f({_al_u2734_o,\PWMC/n24 }),
    .q({\PWMC/FreCntr [1],\PWMC/FreCntr [9]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(~(D*~B)*~(C*~A))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(~(D*~B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b1000110010101111),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000110010101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg1_b20|PWMC/reg1_b8  (
    .a({\PWMC/FreCnt [19],_al_u1580_o}),
    .b({\PWMC/FreCnt [7],\PWMC/FreCnt [24]}),
    .c({\PWMC/FreCntr [20],\PWMC/FreCnt [8]}),
    .ce(\PWMC/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMC/FreCntr [8],\PWMC/FreCntr [24]}),
    .e({open_n20345,\PWMC/FreCntr [8]}),
    .mi({freqC[20],freqC[8]}),
    .f({_al_u2732_o,_al_u1581_o}),
    .q({\PWMC/FreCntr [20],\PWMC/FreCntr [8]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg1_b22|PWMC/reg1_b21  (
    .a({\PWMC/FreCnt [22],_al_u2726_o}),
    .b({\PWMC/FreCnt [23],\PWMC/FreCnt [20]}),
    .c({\PWMC/FreCntr [22],\PWMC/FreCnt [22]}),
    .ce(\PWMC/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMC/FreCntr [23],\PWMC/FreCntr [21]}),
    .e({open_n20362,\PWMC/FreCntr [23]}),
    .mi(freqC[22:21]),
    .f({_al_u1570_o,_al_u2727_o}),
    .q(\PWMC/FreCntr [22:21]));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg1_b23|PWMC/reg1_b0  (
    .b({_al_u1182_o,open_n20381}),
    .c({_al_u1184_o,\PWMC/n11 }),
    .ce(\PWMC/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({_al_u1180_o,\PWMC/n0_lutinv }),
    .mi({freqC[23],freqC[0]}),
    .f({\PWMC/n0_lutinv ,\PWMC/mux3_b0_sel_is_3_o }),
    .q({\PWMC/FreCntr [23],\PWMC/FreCntr [0]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*B*A*~(0@D))"),
    //.LUTF1("(~(D*~B)*~(C*~A))"),
    //.LUTG0("(C*B*A*~(1@D))"),
    //.LUTG1("(~(D*~B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b1000110010101111),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b1000110010101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg1_b26|PWMC/reg1_b13  (
    .a({\PWMC/FreCnt [25],_al_u2733_o}),
    .b({\PWMC/FreCnt [3],_al_u2735_o}),
    .c({\PWMC/FreCntr [26],_al_u2736_o}),
    .ce(\PWMC/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMC/FreCntr [4],\PWMC/FreCnt [12]}),
    .e({open_n20396,\PWMC/FreCntr [13]}),
    .mi({freqC[26],freqC[13]}),
    .f({_al_u2736_o,_al_u2737_o}),
    .q({\PWMC/FreCntr [26],\PWMC/FreCntr [13]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~A*~(~0*C)*~(D@B))"),
    //.LUTF1("(A*~(0@C)*~(D@B))"),
    //.LUTG0("(~A*~(~1*C)*~(D@B))"),
    //.LUTG1("(A*~(1@C)*~(D@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010000000001),
    .INIT_LUTF1(16'b0000100000000010),
    .INIT_LUTG0(16'b0100010000010001),
    .INIT_LUTG1(16'b1000000000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg1_b3|PWMC/reg1_b2  (
    .a({_al_u1582_o,_al_u2716_o}),
    .b(\PWMC/FreCnt [2:1]),
    .c({\PWMC/FreCnt [3],\PWMC/FreCnt [21]}),
    .ce(\PWMC/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMC/FreCntr [2],\PWMC/FreCntr [2]}),
    .e({\PWMC/FreCntr [3],\PWMC/FreCntr [22]}),
    .mi(freqC[3:2]),
    .f({_al_u1583_o,_al_u2717_o}),
    .q(\PWMC/FreCntr [3:2]));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*~C)*~(~D*B))"),
    //.LUTF1("(~(~D*B)*~(~C*A))"),
    //.LUTG0("(A*~(1*~C)*~(~D*B))"),
    //.LUTG1("(~(~D*B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101000100010),
    .INIT_LUTF1(16'b1111010100110001),
    .INIT_LUTG0(16'b1010000000100000),
    .INIT_LUTG1(16'b1111010100110001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg1_b6|PWMC/reg1_b24  (
    .a({\PWMC/FreCnt [10],_al_u2732_o}),
    .b({\PWMC/FreCnt [5],\PWMC/FreCnt [23]}),
    .c({\PWMC/FreCntr [11],\PWMC/FreCnt [5]}),
    .ce(\PWMC/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMC/FreCntr [6],\PWMC/FreCntr [24]}),
    .e({open_n20429,\PWMC/FreCntr [6]}),
    .mi({freqC[6],freqC[24]}),
    .f({_al_u2718_o,_al_u2733_o}),
    .q({\PWMC/FreCntr [6],\PWMC/FreCntr [24]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg2_b0|PWMC/reg3_b0  (
    .a({\PWMC/pnumr [0],_al_u2714_o}),
    .b({pnumC[0],\PWMC/n24 }),
    .c({pnumC[32],pnumcntC[0]}),
    .clk(clk100m),
    .d({pwm_start_stop[28],\PWMC/pnumr [0]}),
    .e({open_n20447,pwm_start_stop[28]}),
    .q({\PWMC/pnumr[0]_keep ,\PWMC/RemaTxNum[0]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011100010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg2_b10|PWMC/reg2_b9  (
    .a(\PWMC/pnumr [10:9]),
    .b({pnumC[10],pnumC[32]}),
    .c({pnumC[32],pnumC[9]}),
    .clk(clk100m),
    .d({pwm_start_stop[28],pwm_start_stop[28]}),
    .q({\PWMC/pnumr[10]_keep ,\PWMC/pnumr[9]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011100010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg2_b11|PWMC/reg2_b8  (
    .a({\PWMC/pnumr [11],\PWMC/pnumr [8]}),
    .b({pnumC[11],pnumC[32]}),
    .c({pnumC[32],pnumC[8]}),
    .clk(clk100m),
    .d({pwm_start_stop[28],pwm_start_stop[28]}),
    .q({\PWMC/pnumr[11]_keep ,\PWMC/pnumr[8]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg2_b12|PWMC/reg3_b12  (
    .a({\PWMC/pnumr [12],_al_u2706_o}),
    .b({pnumC[12],\PWMC/n24 }),
    .c({pnumC[32],pnumcntC[12]}),
    .clk(clk100m),
    .d({pwm_start_stop[28],\PWMC/pnumr [12]}),
    .e({open_n20507,pwm_start_stop[28]}),
    .q({\PWMC/pnumr[12]_keep ,\PWMC/RemaTxNum[12]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg2_b13|PWMC/reg3_b13  (
    .a({\PWMC/pnumr [13],_al_u2704_o}),
    .b({pnumC[13],\PWMC/n24 }),
    .c({pnumC[32],pnumcntC[13]}),
    .clk(clk100m),
    .d({pwm_start_stop[28],\PWMC/pnumr [13]}),
    .e({open_n20529,pwm_start_stop[28]}),
    .q({\PWMC/pnumr[13]_keep ,\PWMC/RemaTxNum[13]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011100010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011100010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg2_b14|PWMC/reg2_b5  (
    .a({\PWMC/pnumr [14],\PWMC/pnumr [5]}),
    .b({pnumC[14],pnumC[32]}),
    .c({pnumC[32],pnumC[5]}),
    .clk(clk100m),
    .d({pwm_start_stop[28],pwm_start_stop[28]}),
    .q({\PWMC/pnumr[14]_keep ,\PWMC/pnumr[5]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011100010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011100010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg2_b15|PWMC/reg2_b4  (
    .a({\PWMC/pnumr [15],\PWMC/pnumr [4]}),
    .b({pnumC[15],pnumC[32]}),
    .c({pnumC[32],pnumC[4]}),
    .clk(clk100m),
    .d({pwm_start_stop[28],pwm_start_stop[28]}),
    .q({\PWMC/pnumr[15]_keep ,\PWMC/pnumr[4]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg2_b16|PWMC/reg3_b16  (
    .a({\PWMC/pnumr [16],_al_u2698_o}),
    .b({pnumC[16],\PWMC/n24 }),
    .c({pnumC[32],pnumcntC[16]}),
    .clk(clk100m),
    .d({pwm_start_stop[28],\PWMC/pnumr [16]}),
    .e({open_n20597,pwm_start_stop[28]}),
    .q({\PWMC/pnumr[16]_keep ,\PWMC/RemaTxNum[16]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg2_b17|PWMC/reg3_b17  (
    .a({\PWMC/pnumr [17],_al_u2696_o}),
    .b({pnumC[17],\PWMC/n24 }),
    .c({pnumC[32],pnumcntC[17]}),
    .clk(clk100m),
    .d({pwm_start_stop[28],\PWMC/pnumr [17]}),
    .e({open_n20619,pwm_start_stop[28]}),
    .q({\PWMC/pnumr[17]_keep ,\PWMC/RemaTxNum[17]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg2_b18|PWMC/reg2_b22  (
    .a({\PWMC/pnumr [18],\PWMC/pnumr [22]}),
    .b({pnumC[18],pnumC[22]}),
    .c({pnumC[32],pnumC[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[28],pwm_start_stop[28]}),
    .q({\PWMC/pnumr[18]_keep ,\PWMC/pnumr[22]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg2_b19|PWMC/reg2_b21  (
    .a({\PWMC/pnumr [19],\PWMC/pnumr [21]}),
    .b({pnumC[19],pnumC[21]}),
    .c({pnumC[32],pnumC[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[28],pwm_start_stop[28]}),
    .q({\PWMC/pnumr[19]_keep ,\PWMC/pnumr[21]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg2_b1|PWMC/reg3_b1  (
    .a({\PWMC/pnumr [1],_al_u2712_o}),
    .b({pnumC[1],\PWMC/n24 }),
    .c({pnumC[32],pnumcntC[1]}),
    .clk(clk100m),
    .d({pwm_start_stop[28],\PWMC/pnumr [1]}),
    .e({open_n20679,pwm_start_stop[28]}),
    .q({\PWMC/pnumr[1]_keep ,\PWMC/RemaTxNum[1]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg2_b20|PWMC/reg3_b20  (
    .a({\PWMC/pnumr [20],_al_u2688_o}),
    .b({pnumC[20],\PWMC/n24 }),
    .c({pnumC[32],pnumcntC[20]}),
    .clk(clk100m),
    .d({pwm_start_stop[28],\PWMC/pnumr [20]}),
    .e({open_n20701,pwm_start_stop[28]}),
    .q({\PWMC/pnumr[20]_keep ,\PWMC/RemaTxNum[20]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg2_b23|PWMC/reg3_b23  (
    .a({\PWMC/pnumr [23],_al_u2682_o}),
    .b({pnumC[23],\PWMC/n24 }),
    .c({pnumC[32],pnumcntC[23]}),
    .clk(clk100m),
    .d({pwm_start_stop[28],\PWMC/pnumr [23]}),
    .e({open_n20723,pwm_start_stop[28]}),
    .q({\PWMC/pnumr[23]_keep ,\PWMC/RemaTxNum[23]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg2_b24|PWMC/reg2_b31  (
    .a({\PWMC/pnumr [24],\PWMC/pnumr [31]}),
    .b({pnumC[24],pnumC[31]}),
    .c({pnumC[32],pnumC[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[28],pwm_start_stop[28]}),
    .q({\PWMC/pnumr[24]_keep ,\PWMC/pnumr[31]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg2_b25|PWMC/reg2_b30  (
    .a({\PWMC/pnumr [25],\PWMC/pnumr [30]}),
    .b({pnumC[25],pnumC[30]}),
    .c({pnumC[32],pnumC[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[28],pwm_start_stop[28]}),
    .q({\PWMC/pnumr[25]_keep ,\PWMC/pnumr[30]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg2_b26|PWMC/reg2_b29  (
    .a({\PWMC/pnumr [26],\PWMC/pnumr [29]}),
    .b({pnumC[26],pnumC[29]}),
    .c({pnumC[32],pnumC[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[28],pwm_start_stop[28]}),
    .q({\PWMC/pnumr[26]_keep ,\PWMC/pnumr[29]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg2_b27|PWMC/reg2_b28  (
    .a({\PWMC/pnumr [27],\PWMC/pnumr [28]}),
    .b({pnumC[27],pnumC[28]}),
    .c({pnumC[32],pnumC[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[28],pwm_start_stop[28]}),
    .q({\PWMC/pnumr[27]_keep ,\PWMC/pnumr[28]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg2_b2|PWMC/reg3_b2  (
    .a({\PWMC/pnumr [2],_al_u2690_o}),
    .b({pnumC[2],\PWMC/n24 }),
    .c({pnumC[32],pnumcntC[2]}),
    .clk(clk100m),
    .d({pwm_start_stop[28],\PWMC/pnumr [2]}),
    .e({open_n20833,pwm_start_stop[28]}),
    .q({\PWMC/pnumr[2]_keep ,\PWMC/RemaTxNum[2]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg2_b3|PWMC/reg3_b3  (
    .a({\PWMC/pnumr [3],_al_u2680_o}),
    .b({pnumC[3],\PWMC/n24 }),
    .c({pnumC[32],pnumcntC[3]}),
    .clk(clk100m),
    .d({pwm_start_stop[28],\PWMC/pnumr [3]}),
    .e({open_n20855,pwm_start_stop[28]}),
    .q({\PWMC/pnumr[3]_keep ,\PWMC/RemaTxNum[3]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg2_b6|PWMC/reg3_b6  (
    .a({\PWMC/pnumr [6],_al_u2674_o}),
    .b({pnumC[32],\PWMC/n24 }),
    .c({pnumC[6],pnumcntC[6]}),
    .clk(clk100m),
    .d({pwm_start_stop[28],\PWMC/pnumr [6]}),
    .e({open_n20877,pwm_start_stop[28]}),
    .q({\PWMC/pnumr[6]_keep ,\PWMC/RemaTxNum[6]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg2_b7|PWMC/reg3_b7  (
    .a({\PWMC/pnumr [7],_al_u2672_o}),
    .b({pnumC[32],\PWMC/n24 }),
    .c({pnumC[7],pnumcntC[7]}),
    .clk(clk100m),
    .d({pwm_start_stop[28],\PWMC/pnumr [7]}),
    .e({open_n20899,pwm_start_stop[28]}),
    .q({\PWMC/pnumr[7]_keep ,\PWMC/RemaTxNum[7]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg3_b10  (
    .a({_al_u2710_o,_al_u2710_o}),
    .b({\PWMC/n24 ,\PWMC/n24 }),
    .c({pnumcntC[10],pnumcntC[10]}),
    .clk(clk100m),
    .d({\PWMC/pnumr [10],\PWMC/pnumr [10]}),
    .mi({open_n20931,pwm_start_stop[28]}),
    .q({open_n20938,\PWMC/RemaTxNum[10]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg3_b11  (
    .a({_al_u2708_o,_al_u2708_o}),
    .b({\PWMC/n24 ,\PWMC/n24 }),
    .c({pnumcntC[11],pnumcntC[11]}),
    .clk(clk100m),
    .d({\PWMC/pnumr [11],\PWMC/pnumr [11]}),
    .mi({open_n20950,pwm_start_stop[28]}),
    .q({open_n20957,\PWMC/RemaTxNum[11]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg3_b14  (
    .a({_al_u2702_o,_al_u2702_o}),
    .b({\PWMC/n24 ,\PWMC/n24 }),
    .c({pnumcntC[14],pnumcntC[14]}),
    .clk(clk100m),
    .d({\PWMC/pnumr [14],\PWMC/pnumr [14]}),
    .mi({open_n20969,pwm_start_stop[28]}),
    .q({open_n20976,\PWMC/RemaTxNum[14]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg3_b15  (
    .a({_al_u2700_o,_al_u2700_o}),
    .b({\PWMC/n24 ,\PWMC/n24 }),
    .c({pnumcntC[15],pnumcntC[15]}),
    .clk(clk100m),
    .d({\PWMC/pnumr [15],\PWMC/pnumr [15]}),
    .mi({open_n20988,pwm_start_stop[28]}),
    .q({open_n20995,\PWMC/RemaTxNum[15]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg3_b18  (
    .a({_al_u2694_o,_al_u2694_o}),
    .b({\PWMC/n24 ,\PWMC/n24 }),
    .c({pnumcntC[18],pnumcntC[18]}),
    .clk(clk100m),
    .d({\PWMC/pnumr [18],\PWMC/pnumr [18]}),
    .mi({open_n21007,pwm_start_stop[28]}),
    .q({open_n21014,\PWMC/RemaTxNum[18]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg3_b19  (
    .a({_al_u2692_o,_al_u2692_o}),
    .b({\PWMC/n24 ,\PWMC/n24 }),
    .c({pnumcntC[19],pnumcntC[19]}),
    .clk(clk100m),
    .d({\PWMC/pnumr [19],\PWMC/pnumr [19]}),
    .mi({open_n21026,pwm_start_stop[28]}),
    .q({open_n21033,\PWMC/RemaTxNum[19]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg3_b21  (
    .a({_al_u2686_o,_al_u2686_o}),
    .b({\PWMC/n24 ,\PWMC/n24 }),
    .c({pnumcntC[21],pnumcntC[21]}),
    .clk(clk100m),
    .d({\PWMC/pnumr [21],\PWMC/pnumr [21]}),
    .mi({open_n21045,pwm_start_stop[28]}),
    .q({open_n21052,\PWMC/RemaTxNum[21]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg3_b22  (
    .a({_al_u2684_o,_al_u2684_o}),
    .b({\PWMC/n24 ,\PWMC/n24 }),
    .c({pnumcntC[22],pnumcntC[22]}),
    .clk(clk100m),
    .d({\PWMC/pnumr [22],\PWMC/pnumr [22]}),
    .mi({open_n21064,pwm_start_stop[28]}),
    .q({open_n21071,\PWMC/RemaTxNum[22]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg3_b4  (
    .a({_al_u2678_o,_al_u2678_o}),
    .b({\PWMC/n24 ,\PWMC/n24 }),
    .c({pnumcntC[4],pnumcntC[4]}),
    .clk(clk100m),
    .d({\PWMC/pnumr [4],\PWMC/pnumr [4]}),
    .mi({open_n21083,pwm_start_stop[28]}),
    .q({open_n21090,\PWMC/RemaTxNum[4]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg3_b5  (
    .a({_al_u2676_o,_al_u2676_o}),
    .b({\PWMC/n24 ,\PWMC/n24 }),
    .c({pnumcntC[5],pnumcntC[5]}),
    .clk(clk100m),
    .d({\PWMC/pnumr [5],\PWMC/pnumr [5]}),
    .mi({open_n21102,pwm_start_stop[28]}),
    .q({open_n21109,\PWMC/RemaTxNum[5]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg3_b8  (
    .a({_al_u2670_o,_al_u2670_o}),
    .b({\PWMC/n24 ,\PWMC/n24 }),
    .c({pnumcntC[8],pnumcntC[8]}),
    .clk(clk100m),
    .d({\PWMC/pnumr [8],\PWMC/pnumr [8]}),
    .mi({open_n21121,pwm_start_stop[28]}),
    .q({open_n21128,\PWMC/RemaTxNum[8]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/reg3_b9  (
    .a({_al_u2668_o,_al_u2668_o}),
    .b({\PWMC/n24 ,\PWMC/n24 }),
    .c({pnumcntC[9],pnumcntC[9]}),
    .clk(clk100m),
    .d({\PWMC/pnumr [9],\PWMC/pnumr [9]}),
    .mi({open_n21140,pwm_start_stop[28]}),
    .q({open_n21147,\PWMC/RemaTxNum[9]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_LSLICE #(
    //.MACRO("PWMC/sub0/ucin_al_u3447"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWMC/sub0/u11_al_u3450  (
    .a({\PWMC/FreCnt [13],\PWMC/FreCnt [11]}),
    .b({\PWMC/FreCnt [14],\PWMC/FreCnt [12]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWMC/sub0/c11 ),
    .f({\PWMC/n12 [13],\PWMC/n12 [11]}),
    .fco(\PWMC/sub0/c15 ),
    .fx({\PWMC/n12 [14],\PWMC/n12 [12]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWMC/sub0/ucin_al_u3447"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWMC/sub0/u15_al_u3451  (
    .a({\PWMC/FreCnt [17],\PWMC/FreCnt [15]}),
    .b({\PWMC/FreCnt [18],\PWMC/FreCnt [16]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWMC/sub0/c15 ),
    .f({\PWMC/n12 [17],\PWMC/n12 [15]}),
    .fco(\PWMC/sub0/c19 ),
    .fx({\PWMC/n12 [18],\PWMC/n12 [16]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWMC/sub0/ucin_al_u3447"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWMC/sub0/u19_al_u3452  (
    .a({\PWMC/FreCnt [21],\PWMC/FreCnt [19]}),
    .b({\PWMC/FreCnt [22],\PWMC/FreCnt [20]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWMC/sub0/c19 ),
    .f({\PWMC/n12 [21],\PWMC/n12 [19]}),
    .fco(\PWMC/sub0/c23 ),
    .fx({\PWMC/n12 [22],\PWMC/n12 [20]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWMC/sub0/ucin_al_u3447"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWMC/sub0/u23_al_u3453  (
    .a({\PWMC/FreCnt [25],\PWMC/FreCnt [23]}),
    .b({\PWMC/FreCnt [26],\PWMC/FreCnt [24]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWMC/sub0/c23 ),
    .f({\PWMC/n12 [25],\PWMC/n12 [23]}),
    .fx({\PWMC/n12 [26],\PWMC/n12 [24]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWMC/sub0/ucin_al_u3447"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWMC/sub0/u3_al_u3448  (
    .a({\PWMC/FreCnt [5],\PWMC/FreCnt [3]}),
    .b({\PWMC/FreCnt [6],\PWMC/FreCnt [4]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWMC/sub0/c3 ),
    .f({\PWMC/n12 [5],\PWMC/n12 [3]}),
    .fco(\PWMC/sub0/c7 ),
    .fx({\PWMC/n12 [6],\PWMC/n12 [4]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWMC/sub0/ucin_al_u3447"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWMC/sub0/u7_al_u3449  (
    .a({\PWMC/FreCnt [9],\PWMC/FreCnt [7]}),
    .b({\PWMC/FreCnt [10],\PWMC/FreCnt [8]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWMC/sub0/c7 ),
    .f({\PWMC/n12 [9],\PWMC/n12 [7]}),
    .fco(\PWMC/sub0/c11 ),
    .fx({\PWMC/n12 [10],\PWMC/n12 [8]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWMC/sub0/ucin_al_u3447"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'h0005),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/sub0/ucin_al_u3447  (
    .a({\PWMC/FreCnt [1],1'b0}),
    .b({\PWMC/FreCnt [2],\PWMC/FreCnt [0]}),
    .c(2'b11),
    .ce(\U_AHB/n28 ),
    .clk(clk100m),
    .d(2'b01),
    .e(2'b01),
    .mi({open_n21258,\U_AHB/h2h_hwdata [2]}),
    .f({\PWMC/n12 [1],open_n21271}),
    .fco(\PWMC/sub0/c3 ),
    .fx({\PWMC/n12 [2],\PWMC/n12 [0]}),
    .q({open_n21272,freqC[2]}));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMC/sub1/u0|PWMC/sub1/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("SUB_CARRY"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000101),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMC/sub1/u0|PWMC/sub1/ucin  (
    .a({pnumcntC[0],1'b0}),
    .b({1'b1,open_n21273}),
    .ce(\U_AHB/n8 ),
    .clk(clk100m),
    .mi({\U_AHB/h2h_hwdata [8],\U_AHB/h2h_hwdata [6]}),
    .f({\PWMC/n26 [0],open_n21289}),
    .fco(\PWMC/sub1/c1 ),
    .q({freq2[8],freq2[6]}));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMC/sub1/u0|PWMC/sub1/ucin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMC/sub1/u10|PWMC/sub1/u9  (
    .a(pnumcntC[10:9]),
    .b(2'b00),
    .fci(\PWMC/sub1/c9 ),
    .f(\PWMC/n26 [10:9]),
    .fco(\PWMC/sub1/c11 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMC/sub1/u0|PWMC/sub1/ucin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMC/sub1/u12|PWMC/sub1/u11  (
    .a(pnumcntC[12:11]),
    .b(2'b00),
    .fci(\PWMC/sub1/c11 ),
    .f(\PWMC/n26 [12:11]),
    .fco(\PWMC/sub1/c13 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMC/sub1/u0|PWMC/sub1/ucin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMC/sub1/u14|PWMC/sub1/u13  (
    .a(pnumcntC[14:13]),
    .b(2'b00),
    .fci(\PWMC/sub1/c13 ),
    .f(\PWMC/n26 [14:13]),
    .fco(\PWMC/sub1/c15 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMC/sub1/u0|PWMC/sub1/ucin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMC/sub1/u16|PWMC/sub1/u15  (
    .a(pnumcntC[16:15]),
    .b(2'b00),
    .fci(\PWMC/sub1/c15 ),
    .f(\PWMC/n26 [16:15]),
    .fco(\PWMC/sub1/c17 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMC/sub1/u0|PWMC/sub1/ucin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMC/sub1/u18|PWMC/sub1/u17  (
    .a(pnumcntC[18:17]),
    .b(2'b00),
    .fci(\PWMC/sub1/c17 ),
    .f(\PWMC/n26 [18:17]),
    .fco(\PWMC/sub1/c19 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMC/sub1/u0|PWMC/sub1/ucin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMC/sub1/u20|PWMC/sub1/u19  (
    .a(pnumcntC[20:19]),
    .b(2'b00),
    .fci(\PWMC/sub1/c19 ),
    .f(\PWMC/n26 [20:19]),
    .fco(\PWMC/sub1/c21 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMC/sub1/u0|PWMC/sub1/ucin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMC/sub1/u22|PWMC/sub1/u21  (
    .a(pnumcntC[22:21]),
    .b(2'b00),
    .fci(\PWMC/sub1/c21 ),
    .f(\PWMC/n26 [22:21]),
    .fco(\PWMC/sub1/c23 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMC/sub1/u0|PWMC/sub1/ucin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMC/sub1/u23_al_u3480  (
    .a({open_n21446,pnumcntC[23]}),
    .b({open_n21447,1'b0}),
    .fci(\PWMC/sub1/c23 ),
    .f({open_n21466,\PWMC/n26 [23]}));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMC/sub1/u0|PWMC/sub1/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMC/sub1/u2|PWMC/sub1/u1  (
    .a(pnumcntC[2:1]),
    .b(2'b00),
    .fci(\PWMC/sub1/c1 ),
    .f(\PWMC/n26 [2:1]),
    .fco(\PWMC/sub1/c3 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMC/sub1/u0|PWMC/sub1/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMC/sub1/u4|PWMC/sub1/u3  (
    .a(pnumcntC[4:3]),
    .b(2'b00),
    .fci(\PWMC/sub1/c3 ),
    .f(\PWMC/n26 [4:3]),
    .fco(\PWMC/sub1/c5 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMC/sub1/u0|PWMC/sub1/ucin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMC/sub1/u6|PWMC/sub1/u5  (
    .a(pnumcntC[6:5]),
    .b(2'b00),
    .fci(\PWMC/sub1/c5 ),
    .f(\PWMC/n26 [6:5]),
    .fco(\PWMC/sub1/c7 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMC/sub1/u0|PWMC/sub1/ucin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMC/sub1/u8|PWMC/sub1/u7  (
    .a(pnumcntC[8:7]),
    .b(2'b00),
    .fci(\PWMC/sub1/c7 ),
    .f(\PWMC/n26 [8:7]),
    .fco(\PWMC/sub1/c9 ));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[0]  (
    .i(\PWMD/RemaTxNum[0]_keep ),
    .o(pnumcntD[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[10]  (
    .i(\PWMD/RemaTxNum[10]_keep ),
    .o(pnumcntD[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[11]  (
    .i(\PWMD/RemaTxNum[11]_keep ),
    .o(pnumcntD[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[12]  (
    .i(\PWMD/RemaTxNum[12]_keep ),
    .o(pnumcntD[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[13]  (
    .i(\PWMD/RemaTxNum[13]_keep ),
    .o(pnumcntD[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[14]  (
    .i(\PWMD/RemaTxNum[14]_keep ),
    .o(pnumcntD[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[15]  (
    .i(\PWMD/RemaTxNum[15]_keep ),
    .o(pnumcntD[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[16]  (
    .i(\PWMD/RemaTxNum[16]_keep ),
    .o(pnumcntD[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[17]  (
    .i(\PWMD/RemaTxNum[17]_keep ),
    .o(pnumcntD[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[18]  (
    .i(\PWMD/RemaTxNum[18]_keep ),
    .o(pnumcntD[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[19]  (
    .i(\PWMD/RemaTxNum[19]_keep ),
    .o(pnumcntD[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[1]  (
    .i(\PWMD/RemaTxNum[1]_keep ),
    .o(pnumcntD[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[20]  (
    .i(\PWMD/RemaTxNum[20]_keep ),
    .o(pnumcntD[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[21]  (
    .i(\PWMD/RemaTxNum[21]_keep ),
    .o(pnumcntD[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[22]  (
    .i(\PWMD/RemaTxNum[22]_keep ),
    .o(pnumcntD[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[23]  (
    .i(\PWMD/RemaTxNum[23]_keep ),
    .o(pnumcntD[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[2]  (
    .i(\PWMD/RemaTxNum[2]_keep ),
    .o(pnumcntD[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[3]  (
    .i(\PWMD/RemaTxNum[3]_keep ),
    .o(pnumcntD[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[4]  (
    .i(\PWMD/RemaTxNum[4]_keep ),
    .o(pnumcntD[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[5]  (
    .i(\PWMD/RemaTxNum[5]_keep ),
    .o(pnumcntD[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[6]  (
    .i(\PWMD/RemaTxNum[6]_keep ),
    .o(pnumcntD[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[7]  (
    .i(\PWMD/RemaTxNum[7]_keep ),
    .o(pnumcntD[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[8]  (
    .i(\PWMD/RemaTxNum[8]_keep ),
    .o(pnumcntD[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[9]  (
    .i(\PWMD/RemaTxNum[9]_keep ),
    .o(pnumcntD[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_dir  (
    .i(\PWMD/dir_keep ),
    .o(dir_pad[13]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[0]  (
    .i(\PWMD/pnumr[0]_keep ),
    .o(\PWMD/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[10]  (
    .i(\PWMD/pnumr[10]_keep ),
    .o(\PWMD/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[11]  (
    .i(\PWMD/pnumr[11]_keep ),
    .o(\PWMD/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[12]  (
    .i(\PWMD/pnumr[12]_keep ),
    .o(\PWMD/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[13]  (
    .i(\PWMD/pnumr[13]_keep ),
    .o(\PWMD/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[14]  (
    .i(\PWMD/pnumr[14]_keep ),
    .o(\PWMD/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[15]  (
    .i(\PWMD/pnumr[15]_keep ),
    .o(\PWMD/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[16]  (
    .i(\PWMD/pnumr[16]_keep ),
    .o(\PWMD/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[17]  (
    .i(\PWMD/pnumr[17]_keep ),
    .o(\PWMD/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[18]  (
    .i(\PWMD/pnumr[18]_keep ),
    .o(\PWMD/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[19]  (
    .i(\PWMD/pnumr[19]_keep ),
    .o(\PWMD/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[1]  (
    .i(\PWMD/pnumr[1]_keep ),
    .o(\PWMD/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[20]  (
    .i(\PWMD/pnumr[20]_keep ),
    .o(\PWMD/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[21]  (
    .i(\PWMD/pnumr[21]_keep ),
    .o(\PWMD/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[22]  (
    .i(\PWMD/pnumr[22]_keep ),
    .o(\PWMD/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[23]  (
    .i(\PWMD/pnumr[23]_keep ),
    .o(\PWMD/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[24]  (
    .i(\PWMD/pnumr[24]_keep ),
    .o(\PWMD/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[25]  (
    .i(\PWMD/pnumr[25]_keep ),
    .o(\PWMD/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[26]  (
    .i(\PWMD/pnumr[26]_keep ),
    .o(\PWMD/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[27]  (
    .i(\PWMD/pnumr[27]_keep ),
    .o(\PWMD/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[28]  (
    .i(\PWMD/pnumr[28]_keep ),
    .o(\PWMD/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[29]  (
    .i(\PWMD/pnumr[29]_keep ),
    .o(\PWMD/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[2]  (
    .i(\PWMD/pnumr[2]_keep ),
    .o(\PWMD/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[30]  (
    .i(\PWMD/pnumr[30]_keep ),
    .o(\PWMD/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[31]  (
    .i(\PWMD/pnumr[31]_keep ),
    .o(\PWMD/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[3]  (
    .i(\PWMD/pnumr[3]_keep ),
    .o(\PWMD/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[4]  (
    .i(\PWMD/pnumr[4]_keep ),
    .o(\PWMD/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[5]  (
    .i(\PWMD/pnumr[5]_keep ),
    .o(\PWMD/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[6]  (
    .i(\PWMD/pnumr[6]_keep ),
    .o(\PWMD/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[7]  (
    .i(\PWMD/pnumr[7]_keep ),
    .o(\PWMD/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[8]  (
    .i(\PWMD/pnumr[8]_keep ),
    .o(\PWMD/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[9]  (
    .i(\PWMD/pnumr[9]_keep ),
    .o(\PWMD/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pwm  (
    .i(\PWMD/pwm_keep ),
    .o(pwm_pad[13]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_stopreq  (
    .i(\PWMD/stopreq_keep ),
    .o(\PWMD/stopreq ));  // src/OnePWM.v(14)
  EF2_PHY_MSLICE #(
    //.LUT0("(D*~(C)*~((~0*~(B*A)))+D*C*~((~0*~(B*A)))+~(D)*C*(~0*~(B*A))+D*C*(~0*~(B*A)))"),
    //.LUT1("(D*~(C)*~((~1*~(B*A)))+D*C*~((~1*~(B*A)))+~(D)*C*(~1*~(B*A))+D*C*(~1*~(B*A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111100001110000),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/dir_reg  (
    .a({\PWMD/n24 ,\PWMD/n24 }),
    .b({\PWMD/n25_neg_lutinv ,\PWMD/n25_neg_lutinv }),
    .c({dir_pad[13],dir_pad[13]}),
    .clk(clk100m),
    .d({\PWMD/pnumr [31],\PWMD/pnumr [31]}),
    .mi({open_n21571,pwm_start_stop[29]}),
    .q({open_n21578,\PWMD/dir_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("~(~0*~(D*C*B*A))"),
    //.LUT1("~(~1*~(D*C*B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b1111111111111111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMD/pwm_reg  (
    .a({_al_u1590_o,_al_u1590_o}),
    .b({_al_u1596_o,_al_u1596_o}),
    .c({_al_u1598_o,_al_u1598_o}),
    .clk(clk100m),
    .d({_al_u1600_o,_al_u1600_o}),
    .mi({open_n21590,pwm_pad[13]}),
    .sr(\PWMD/u14_sel_is_1_o ),
    .q({open_n21596,\PWMD/pwm_keep }));  // src/OnePWM.v(45)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMD/reg0_b0|PWMD/reg0_b8  (
    .b({\PWMD/n12 [0],\PWMD/n12 [8]}),
    .c({freqD[0],freqD[8]}),
    .clk(clk100m),
    .d({\PWMD/n0_lutinv ,\PWMD/n0_lutinv }),
    .sr(\PWMD/n11 ),
    .q({\PWMD/FreCnt [0],\PWMD/FreCnt [8]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMD/reg0_b10|PWMD/reg0_b7  (
    .b({\PWMD/n12 [10],\PWMD/n12 [7]}),
    .c({freqD[10],freqD[7]}),
    .clk(clk100m),
    .d({\PWMD/n0_lutinv ,\PWMD/n0_lutinv }),
    .sr(\PWMD/n11 ),
    .q({\PWMD/FreCnt [10],\PWMD/FreCnt [7]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMD/reg0_b11|PWMD/reg0_b17  (
    .b({\PWMD/n12 [11],\PWMD/n12 [17]}),
    .c({freqD[11],freqD[17]}),
    .clk(clk100m),
    .d({\PWMD/n0_lutinv ,\PWMD/n0_lutinv }),
    .sr(\PWMD/n11 ),
    .q({\PWMD/FreCnt [11],\PWMD/FreCnt [17]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMD/reg0_b14|PWMD/reg0_b13  (
    .b(\PWMD/n12 [14:13]),
    .c(freqD[14:13]),
    .clk(clk100m),
    .d({\PWMD/n0_lutinv ,\PWMD/n0_lutinv }),
    .sr(\PWMD/n11 ),
    .q(\PWMD/FreCnt [14:13]));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMD/reg0_b16|PWMD/reg0_b9  (
    .b({\PWMD/n12 [16],\PWMD/n12 [9]}),
    .c({freqD[16],freqD[9]}),
    .clk(clk100m),
    .d({\PWMD/n0_lutinv ,\PWMD/n0_lutinv }),
    .sr(\PWMD/n11 ),
    .q({\PWMD/FreCnt [16],\PWMD/FreCnt [9]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMD/reg0_b18|PWMD/reg0_b5  (
    .b({\PWMD/n12 [18],\PWMD/n12 [5]}),
    .c({freqD[18],freqD[5]}),
    .clk(clk100m),
    .d({\PWMD/n0_lutinv ,\PWMD/n0_lutinv }),
    .sr(\PWMD/n11 ),
    .q({\PWMD/FreCnt [18],\PWMD/FreCnt [5]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMD/reg0_b20|PWMD/reg0_b4  (
    .b({\PWMD/n12 [20],\PWMD/n12 [4]}),
    .c({freqD[20],freqD[4]}),
    .clk(clk100m),
    .d({\PWMD/n0_lutinv ,\PWMD/n0_lutinv }),
    .sr(\PWMD/n11 ),
    .q({\PWMD/FreCnt [20],\PWMD/FreCnt [4]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMD/reg0_b21|PWMD/reg0_b3  (
    .b({\PWMD/n12 [21],\PWMD/n12 [3]}),
    .c({freqD[21],freqD[3]}),
    .clk(clk100m),
    .d({\PWMD/n0_lutinv ,\PWMD/n0_lutinv }),
    .sr(\PWMD/n11 ),
    .q({\PWMD/FreCnt [21],\PWMD/FreCnt [3]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMD/reg0_b22|PWMD/reg0_b25  (
    .b({\PWMD/n12 [22],\PWMD/n12 [25]}),
    .c({freqD[22],freqD[25]}),
    .clk(clk100m),
    .d({\PWMD/n0_lutinv ,\PWMD/n0_lutinv }),
    .sr(\PWMD/n11 ),
    .q({\PWMD/FreCnt [22],\PWMD/FreCnt [25]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMD/reg0_b2|PWMD/reg0_b24  (
    .b({\PWMD/n12 [2],\PWMD/n12 [24]}),
    .c({freqD[2],freqD[24]}),
    .clk(clk100m),
    .d({\PWMD/n0_lutinv ,\PWMD/n0_lutinv }),
    .sr(\PWMD/n11 ),
    .q({\PWMD/FreCnt [2],\PWMD/FreCnt [24]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*B*A*~(0@D))"),
    //.LUTF1("(~(C@B)*~(D@A))"),
    //.LUTG0("(C*B*A*~(1@D))"),
    //.LUTG1("(~(C@B)*~(D@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b1000001001000001),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b1000001001000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg1_b10|PWMD/reg1_b12  (
    .a({\PWMD/FreCnt [22],_al_u2797_o}),
    .b({\PWMD/FreCnt [9],_al_u2798_o}),
    .c({\PWMD/FreCntr [10],_al_u2799_o}),
    .ce(\PWMD/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMD/FreCntr [23],\PWMD/FreCnt [11]}),
    .e({open_n21805,\PWMD/FreCntr [12]}),
    .mi({freqD[10],freqD[12]}),
    .f({_al_u2798_o,_al_u2800_o}),
    .q({\PWMD/FreCntr [10],\PWMD/FreCntr [12]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~A*~(~0*C)*~(D@B))"),
    //.LUTF1("(~(~D*B)*~(C*~A))"),
    //.LUTG0("(~A*~(~1*C)*~(D@B))"),
    //.LUTG1("(~(~D*B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010000000001),
    .INIT_LUTF1(16'b1010111100100011),
    .INIT_LUTG0(16'b0100010000010001),
    .INIT_LUTG1(16'b1010111100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg1_b13|PWMD/reg1_b11  (
    .a({\PWMD/FreCnt [12],_al_u2809_o}),
    .b({\PWMD/FreCnt [8],\PWMD/FreCnt [10]}),
    .c({\PWMD/FreCntr [13],\PWMD/FreCnt [12]}),
    .ce(\PWMD/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMD/FreCntr [9],\PWMD/FreCntr [11]}),
    .e({open_n21822,\PWMD/FreCntr [13]}),
    .mi({freqD[13],freqD[11]}),
    .f({_al_u2795_o,_al_u2810_o}),
    .q({\PWMD/FreCntr [13],\PWMD/FreCntr [11]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(D*~B)*~(~C*A))"),
    //.LUTF1("(~(~D*B)*~(C*~A))"),
    //.LUTG0("(~(D*~B)*~(~C*A))"),
    //.LUTG1("(~(~D*B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100010011110101),
    .INIT_LUTF1(16'b1010111100100011),
    .INIT_LUTG0(16'b1100010011110101),
    .INIT_LUTG1(16'b1010111100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg1_b16|PWMD/reg1_b20  (
    .a({\PWMD/FreCnt [15],\PWMD/FreCnt [15]}),
    .b({\PWMD/FreCnt [19],\PWMD/FreCnt [19]}),
    .c({\PWMD/FreCntr [16],\PWMD/FreCntr [16]}),
    .ce(\PWMD/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMD/FreCntr [20],\PWMD/FreCntr [20]}),
    .mi({freqD[16],freqD[20]}),
    .f({_al_u2811_o,_al_u2799_o}),
    .q({\PWMD/FreCntr [16],\PWMD/FreCntr [20]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(D@B)*~(C@A))"),
    //.LUT1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000010000100001),
    .INIT_LUT1(16'b1000010000100001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg1_b17|PWMD/reg1_b4  (
    .a({\PWMD/FreCnt [16],\PWMD/FreCnt [16]}),
    .b({\PWMD/FreCnt [2],\PWMD/FreCnt [4]}),
    .c(\PWMD/FreCntr [17:16]),
    .ce(\PWMD/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMD/FreCntr [3],\PWMD/FreCntr [4]}),
    .mi({freqD[17],freqD[4]}),
    .f({_al_u2803_o,_al_u1585_o}),
    .q({\PWMD/FreCntr [17],\PWMD/FreCntr [4]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(~C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg1_b18|PWMD/reg1_b9  (
    .c({\PWMD/FreCntr [18],\PWMD/FreCntr [9]}),
    .ce(\PWMD/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMD/FreCnt [17],\PWMD/FreCnt [8]}),
    .mi({freqD[18],freqD[9]}),
    .f({_al_u2809_o,_al_u2813_o}),
    .q({\PWMD/FreCntr [18],\PWMD/FreCntr [9]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*~C)*~(D*~B))"),
    //.LUTF1("(A*~(~0*C)*~(D@B))"),
    //.LUTG0("(A*~(1*~C)*~(D*~B))"),
    //.LUTG1("(A*~(~1*C)*~(D@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000100010101010),
    .INIT_LUTF1(16'b0000100000000010),
    .INIT_LUTG0(16'b1000000010100000),
    .INIT_LUTG1(16'b1000100000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg1_b19|PWMD/reg1_b8  (
    .a({_al_u2796_o,_al_u2795_o}),
    .b({\PWMD/FreCnt [18],\PWMD/FreCnt [1]}),
    .c({\PWMD/FreCnt [7],\PWMD/FreCnt [7]}),
    .ce(\PWMD/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMD/FreCntr [19],\PWMD/FreCntr [2]}),
    .e({\PWMD/FreCntr [8],\PWMD/FreCntr [8]}),
    .mi({freqD[19],freqD[8]}),
    .f({_al_u2797_o,_al_u2796_o}),
    .q({\PWMD/FreCntr [19],\PWMD/FreCntr [8]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~A*~(0@C)*~(D*~B))"),
    //.LUTF1("(~C*D)"),
    //.LUTG0("(~A*~(1@C)*~(D*~B))"),
    //.LUTG1("(~C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010000000101),
    .INIT_LUTF1(16'b0000111100000000),
    .INIT_LUTG0(16'b0100000001010000),
    .INIT_LUTG1(16'b0000111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg1_b1|PWMD/reg1_b22  (
    .a({open_n21909,_al_u2813_o}),
    .b({open_n21910,\PWMD/FreCnt [0]}),
    .c({\PWMD/FreCntr [1],\PWMD/FreCnt [21]}),
    .ce(\PWMD/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMD/FreCnt [0],\PWMD/FreCntr [1]}),
    .e({open_n21911,\PWMD/FreCntr [22]}),
    .mi({freqD[1],freqD[22]}),
    .f({_al_u2815_o,_al_u2814_o}),
    .q({\PWMD/FreCntr [1],\PWMD/FreCntr [22]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~A*~(~0*C)*~(D@B))"),
    //.LUTF1("(~(D*~B)*~(C*~A))"),
    //.LUTG0("(~A*~(~1*C)*~(D@B))"),
    //.LUTG1("(~(D*~B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010000000001),
    .INIT_LUTF1(16'b1000110010101111),
    .INIT_LUTG0(16'b0100010000010001),
    .INIT_LUTG1(16'b1000110010101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg1_b24|PWMD/reg1_b15  (
    .a({\PWMD/FreCnt [17],_al_u2815_o}),
    .b({\PWMD/FreCnt [23],\PWMD/FreCnt [14]}),
    .c({\PWMD/FreCntr [18],\PWMD/FreCnt [23]}),
    .ce(\PWMD/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMD/FreCntr [24],\PWMD/FreCntr [15]}),
    .e({open_n21928,\PWMD/FreCntr [24]}),
    .mi({freqD[24],freqD[15]}),
    .f({_al_u2805_o,_al_u2816_o}),
    .q({\PWMD/FreCntr [24],\PWMD/FreCntr [15]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~B*~(0@C)*~(D*~A))"),
    //.LUTF1("(A*~(~D*C)*~(~0*B))"),
    //.LUTG0("(~B*~(1@C)*~(D*~A))"),
    //.LUTG1("(A*~(~D*C)*~(~1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001000000011),
    .INIT_LUTF1(16'b0010001000000010),
    .INIT_LUTG0(16'b0010000000110000),
    .INIT_LUTG1(16'b1010101000001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg1_b2|PWMD/reg1_b14  (
    .a({_al_u2805_o,\PWMD/FreCnt [13]}),
    .b({\PWMD/FreCnt [1],\PWMD/FreCnt [26]}),
    .c({\PWMD/FreCnt [13],\PWMD/FreCnt [3]}),
    .ce(\PWMD/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMD/FreCntr [14],\PWMD/FreCntr [14]}),
    .e({\PWMD/FreCntr [2],\PWMD/FreCntr [4]}),
    .mi({freqD[2],freqD[14]}),
    .f({_al_u2806_o,_al_u2807_o}),
    .q({\PWMD/FreCntr [2],\PWMD/FreCntr [14]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(D@B)*~(C@A))"),
    //.LUT1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000010000100001),
    .INIT_LUT1(16'b1000010000100001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg1_b5|PWMD/reg1_b7  (
    .a({\PWMD/FreCnt [4],\PWMD/FreCnt [7]}),
    .b({\PWMD/FreCnt [6],\PWMD/FreCnt [9]}),
    .c({\PWMD/FreCntr [5],\PWMD/FreCntr [7]}),
    .ce(\PWMD/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMD/FreCntr [7],\PWMD/FreCntr [9]}),
    .mi({freqD[5],freqD[7]}),
    .f({_al_u2801_o,_al_u1597_o}),
    .q({\PWMD/FreCntr [5],\PWMD/FreCntr [7]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(D*~(C@B))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(D*~(C@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b1100001100000000),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1100001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg1_b6|PWMD/reg1_b26  (
    .a({open_n21975,_al_u2803_o}),
    .b({\PWMD/FreCnt [6],\PWMD/FreCnt [25]}),
    .c({\PWMD/FreCntr [6],\PWMD/FreCnt [5]}),
    .ce(\PWMD/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({_al_u1591_o,\PWMD/FreCntr [26]}),
    .e({open_n21976,\PWMD/FreCntr [6]}),
    .mi({freqD[6],freqD[26]}),
    .f({_al_u1592_o,_al_u2804_o}),
    .q({\PWMD/FreCntr [6],\PWMD/FreCntr [26]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011100010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011100010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg2_b0|PWMD/reg2_b9  (
    .a({\PWMD/pnumr [0],\PWMD/pnumr [9]}),
    .b({pnumD[0],pnumD[32]}),
    .c({pnumD[32],pnumD[9]}),
    .clk(clk100m),
    .d({pwm_start_stop[29],pwm_start_stop[29]}),
    .q({\PWMD/pnumr[0]_keep ,\PWMD/pnumr[9]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg2_b10|PWMD/reg3_b10  (
    .a({\PWMD/pnumr [10],_al_u2789_o}),
    .b({pnumD[10],\PWMD/n24 }),
    .c({pnumD[32],pnumcntD[10]}),
    .clk(clk100m),
    .d({pwm_start_stop[29],\PWMD/pnumr [10]}),
    .e({open_n22017,pwm_start_stop[29]}),
    .q({\PWMD/pnumr[10]_keep ,\PWMD/RemaTxNum[10]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011100010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011100010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg2_b11|PWMD/reg2_b6  (
    .a({\PWMD/pnumr [11],\PWMD/pnumr [6]}),
    .b({pnumD[11],pnumD[32]}),
    .c({pnumD[32],pnumD[6]}),
    .clk(clk100m),
    .d({pwm_start_stop[29],pwm_start_stop[29]}),
    .q({\PWMD/pnumr[11]_keep ,\PWMD/pnumr[6]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011100010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg2_b12|PWMD/reg2_b5  (
    .a({\PWMD/pnumr [12],\PWMD/pnumr [5]}),
    .b({pnumD[12],pnumD[32]}),
    .c({pnumD[32],pnumD[5]}),
    .clk(clk100m),
    .d({pwm_start_stop[29],pwm_start_stop[29]}),
    .q({\PWMD/pnumr[12]_keep ,\PWMD/pnumr[5]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg2_b13|PWMD/reg3_b13  (
    .a({\PWMD/pnumr [13],_al_u2783_o}),
    .b({pnumD[13],\PWMD/n24 }),
    .c({pnumD[32],pnumcntD[13]}),
    .clk(clk100m),
    .d({pwm_start_stop[29],\PWMD/pnumr [13]}),
    .e({open_n22081,pwm_start_stop[29]}),
    .q({\PWMD/pnumr[13]_keep ,\PWMD/RemaTxNum[13]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg2_b14|PWMD/reg3_b14  (
    .a({\PWMD/pnumr [14],_al_u2781_o}),
    .b({pnumD[14],\PWMD/n24 }),
    .c({pnumD[32],pnumcntD[14]}),
    .clk(clk100m),
    .d({pwm_start_stop[29],\PWMD/pnumr [14]}),
    .e({open_n22103,pwm_start_stop[29]}),
    .q({\PWMD/pnumr[14]_keep ,\PWMD/RemaTxNum[14]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg2_b15|PWMD/reg2_b23  (
    .a({\PWMD/pnumr [15],\PWMD/pnumr [23]}),
    .b({pnumD[15],pnumD[23]}),
    .c({pnumD[32],pnumD[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[29],pwm_start_stop[29]}),
    .q({\PWMD/pnumr[15]_keep ,\PWMD/pnumr[23]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg2_b16|PWMD/reg2_b22  (
    .a({\PWMD/pnumr [16],\PWMD/pnumr [22]}),
    .b({pnumD[16],pnumD[22]}),
    .c({pnumD[32],pnumD[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[29],pwm_start_stop[29]}),
    .q({\PWMD/pnumr[16]_keep ,\PWMD/pnumr[22]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg2_b17|PWMD/reg3_b17  (
    .a({\PWMD/pnumr [17],_al_u2775_o}),
    .b({pnumD[17],\PWMD/n24 }),
    .c({pnumD[32],pnumcntD[17]}),
    .clk(clk100m),
    .d({pwm_start_stop[29],\PWMD/pnumr [17]}),
    .e({open_n22167,pwm_start_stop[29]}),
    .q({\PWMD/pnumr[17]_keep ,\PWMD/RemaTxNum[17]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg2_b18|PWMD/reg3_b18  (
    .a({\PWMD/pnumr [18],_al_u2773_o}),
    .b({pnumD[18],\PWMD/n24 }),
    .c({pnumD[32],pnumcntD[18]}),
    .clk(clk100m),
    .d({pwm_start_stop[29],\PWMD/pnumr [18]}),
    .e({open_n22189,pwm_start_stop[29]}),
    .q({\PWMD/pnumr[18]_keep ,\PWMD/RemaTxNum[18]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg2_b19|PWMD/reg2_b2  (
    .a({\PWMD/pnumr [19],\PWMD/pnumr [2]}),
    .b({pnumD[19],pnumD[2]}),
    .c({pnumD[32],pnumD[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[29],pwm_start_stop[29]}),
    .q({\PWMD/pnumr[19]_keep ,\PWMD/pnumr[2]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg2_b1|PWMD/reg3_b1  (
    .a({\PWMD/pnumr [1],_al_u2791_o}),
    .b({pnumD[1],\PWMD/n24 }),
    .c({pnumD[32],pnumcntD[1]}),
    .clk(clk100m),
    .d({pwm_start_stop[29],\PWMD/pnumr [1]}),
    .e({open_n22234,pwm_start_stop[29]}),
    .q({\PWMD/pnumr[1]_keep ,\PWMD/RemaTxNum[1]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg2_b20|PWMD/reg3_b20  (
    .a({\PWMD/pnumr [20],_al_u2767_o}),
    .b({pnumD[20],\PWMD/n24 }),
    .c({pnumD[32],pnumcntD[20]}),
    .clk(clk100m),
    .d({pwm_start_stop[29],\PWMD/pnumr [20]}),
    .e({open_n22256,pwm_start_stop[29]}),
    .q({\PWMD/pnumr[20]_keep ,\PWMD/RemaTxNum[20]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg2_b21|PWMD/reg3_b21  (
    .a({\PWMD/pnumr [21],_al_u2765_o}),
    .b({pnumD[21],\PWMD/n24 }),
    .c({pnumD[32],pnumcntD[21]}),
    .clk(clk100m),
    .d({pwm_start_stop[29],\PWMD/pnumr [21]}),
    .e({open_n22278,pwm_start_stop[29]}),
    .q({\PWMD/pnumr[21]_keep ,\PWMD/RemaTxNum[21]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg2_b24|PWMD/reg2_b31  (
    .a({\PWMD/pnumr [24],\PWMD/pnumr [31]}),
    .b({pnumD[24],pnumD[31]}),
    .c({pnumD[32],pnumD[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[29],pwm_start_stop[29]}),
    .q({\PWMD/pnumr[24]_keep ,\PWMD/pnumr[31]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg2_b25|PWMD/reg2_b30  (
    .a({\PWMD/pnumr [25],\PWMD/pnumr [30]}),
    .b({pnumD[25],pnumD[30]}),
    .c({pnumD[32],pnumD[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[29],pwm_start_stop[29]}),
    .q({\PWMD/pnumr[25]_keep ,\PWMD/pnumr[30]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg2_b26|PWMD/reg2_b29  (
    .a({\PWMD/pnumr [26],\PWMD/pnumr [29]}),
    .b({pnumD[26],pnumD[29]}),
    .c({pnumD[32],pnumD[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[29],pwm_start_stop[29]}),
    .q({\PWMD/pnumr[26]_keep ,\PWMD/pnumr[29]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg2_b27|PWMD/reg2_b28  (
    .a({\PWMD/pnumr [27],\PWMD/pnumr [28]}),
    .b({pnumD[27],pnumD[28]}),
    .c({pnumD[32],pnumD[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[29],pwm_start_stop[29]}),
    .q({\PWMD/pnumr[27]_keep ,\PWMD/pnumr[28]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg2_b3|PWMD/reg3_b3  (
    .a({\PWMD/pnumr [3],_al_u2759_o}),
    .b({pnumD[3],\PWMD/n24 }),
    .c({pnumD[32],pnumcntD[3]}),
    .clk(clk100m),
    .d({pwm_start_stop[29],\PWMD/pnumr [3]}),
    .e({open_n22388,pwm_start_stop[29]}),
    .q({\PWMD/pnumr[3]_keep ,\PWMD/RemaTxNum[3]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg2_b4|PWMD/reg3_b4  (
    .a({\PWMD/pnumr [4],_al_u2757_o}),
    .b({pnumD[32],\PWMD/n24 }),
    .c({pnumD[4],pnumcntD[4]}),
    .clk(clk100m),
    .d({pwm_start_stop[29],\PWMD/pnumr [4]}),
    .e({open_n22410,pwm_start_stop[29]}),
    .q({\PWMD/pnumr[4]_keep ,\PWMD/RemaTxNum[4]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg2_b7|PWMD/reg3_b7  (
    .a({\PWMD/pnumr [7],_al_u2751_o}),
    .b({pnumD[32],\PWMD/n24 }),
    .c({pnumD[7],pnumcntD[7]}),
    .clk(clk100m),
    .d({pwm_start_stop[29],\PWMD/pnumr [7]}),
    .e({open_n22432,pwm_start_stop[29]}),
    .q({\PWMD/pnumr[7]_keep ,\PWMD/RemaTxNum[7]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg2_b8|PWMD/reg3_b8  (
    .a({\PWMD/pnumr [8],_al_u2749_o}),
    .b({pnumD[32],\PWMD/n24 }),
    .c({pnumD[8],pnumcntD[8]}),
    .clk(clk100m),
    .d({pwm_start_stop[29],\PWMD/pnumr [8]}),
    .e({open_n22454,pwm_start_stop[29]}),
    .q({\PWMD/pnumr[8]_keep ,\PWMD/RemaTxNum[8]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg3_b0  (
    .a({_al_u2793_o,_al_u2793_o}),
    .b({\PWMD/n24 ,\PWMD/n24 }),
    .c({pnumcntD[0],pnumcntD[0]}),
    .clk(clk100m),
    .d({\PWMD/pnumr [0],\PWMD/pnumr [0]}),
    .mi({open_n22486,pwm_start_stop[29]}),
    .q({open_n22493,\PWMD/RemaTxNum[0]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg3_b11  (
    .a({_al_u2787_o,_al_u2787_o}),
    .b({\PWMD/n24 ,\PWMD/n24 }),
    .c({pnumcntD[11],pnumcntD[11]}),
    .clk(clk100m),
    .d({\PWMD/pnumr [11],\PWMD/pnumr [11]}),
    .mi({open_n22505,pwm_start_stop[29]}),
    .q({open_n22512,\PWMD/RemaTxNum[11]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg3_b12  (
    .a({_al_u2785_o,_al_u2785_o}),
    .b({\PWMD/n24 ,\PWMD/n24 }),
    .c({pnumcntD[12],pnumcntD[12]}),
    .clk(clk100m),
    .d({\PWMD/pnumr [12],\PWMD/pnumr [12]}),
    .mi({open_n22524,pwm_start_stop[29]}),
    .q({open_n22531,\PWMD/RemaTxNum[12]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg3_b15  (
    .a({_al_u2779_o,_al_u2779_o}),
    .b({\PWMD/n24 ,\PWMD/n24 }),
    .c({pnumcntD[15],pnumcntD[15]}),
    .clk(clk100m),
    .d({\PWMD/pnumr [15],\PWMD/pnumr [15]}),
    .mi({open_n22543,pwm_start_stop[29]}),
    .q({open_n22550,\PWMD/RemaTxNum[15]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg3_b16  (
    .a({_al_u2777_o,_al_u2777_o}),
    .b({\PWMD/n24 ,\PWMD/n24 }),
    .c({pnumcntD[16],pnumcntD[16]}),
    .clk(clk100m),
    .d({\PWMD/pnumr [16],\PWMD/pnumr [16]}),
    .mi({open_n22562,pwm_start_stop[29]}),
    .q({open_n22569,\PWMD/RemaTxNum[16]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg3_b19  (
    .a({_al_u2771_o,_al_u2771_o}),
    .b({\PWMD/n24 ,\PWMD/n24 }),
    .c({pnumcntD[19],pnumcntD[19]}),
    .clk(clk100m),
    .d({\PWMD/pnumr [19],\PWMD/pnumr [19]}),
    .mi({open_n22581,pwm_start_stop[29]}),
    .q({open_n22588,\PWMD/RemaTxNum[19]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg3_b2  (
    .a({_al_u2769_o,_al_u2769_o}),
    .b({\PWMD/n24 ,\PWMD/n24 }),
    .c({pnumcntD[2],pnumcntD[2]}),
    .clk(clk100m),
    .d({\PWMD/pnumr [2],\PWMD/pnumr [2]}),
    .mi({open_n22600,pwm_start_stop[29]}),
    .q({open_n22607,\PWMD/RemaTxNum[2]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg3_b22  (
    .a({_al_u2763_o,_al_u2763_o}),
    .b({\PWMD/n24 ,\PWMD/n24 }),
    .c({pnumcntD[22],pnumcntD[22]}),
    .clk(clk100m),
    .d({\PWMD/pnumr [22],\PWMD/pnumr [22]}),
    .mi({open_n22619,pwm_start_stop[29]}),
    .q({open_n22626,\PWMD/RemaTxNum[22]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg3_b23  (
    .a({_al_u2761_o,_al_u2761_o}),
    .b({\PWMD/n24 ,\PWMD/n24 }),
    .c({pnumcntD[23],pnumcntD[23]}),
    .clk(clk100m),
    .d({\PWMD/pnumr [23],\PWMD/pnumr [23]}),
    .mi({open_n22638,pwm_start_stop[29]}),
    .q({open_n22645,\PWMD/RemaTxNum[23]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg3_b5  (
    .a({_al_u2755_o,_al_u2755_o}),
    .b({\PWMD/n24 ,\PWMD/n24 }),
    .c({pnumcntD[5],pnumcntD[5]}),
    .clk(clk100m),
    .d({\PWMD/pnumr [5],\PWMD/pnumr [5]}),
    .mi({open_n22657,pwm_start_stop[29]}),
    .q({open_n22664,\PWMD/RemaTxNum[5]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg3_b6  (
    .a({_al_u2753_o,_al_u2753_o}),
    .b({\PWMD/n24 ,\PWMD/n24 }),
    .c({pnumcntD[6],pnumcntD[6]}),
    .clk(clk100m),
    .d({\PWMD/pnumr [6],\PWMD/pnumr [6]}),
    .mi({open_n22676,pwm_start_stop[29]}),
    .q({open_n22683,\PWMD/RemaTxNum[6]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMD/reg3_b9  (
    .a({_al_u2747_o,_al_u2747_o}),
    .b({\PWMD/n24 ,\PWMD/n24 }),
    .c({pnumcntD[9],pnumcntD[9]}),
    .clk(clk100m),
    .d({\PWMD/pnumr [9],\PWMD/pnumr [9]}),
    .mi({open_n22695,pwm_start_stop[29]}),
    .q({open_n22702,\PWMD/RemaTxNum[9]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_LSLICE #(
    //.MACRO("PWMD/sub0/ucin_al_u3454"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWMD/sub0/u11_al_u3457  (
    .a({\PWMD/FreCnt [13],\PWMD/FreCnt [11]}),
    .b({\PWMD/FreCnt [14],\PWMD/FreCnt [12]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWMD/sub0/c11 ),
    .f({\PWMD/n12 [13],\PWMD/n12 [11]}),
    .fco(\PWMD/sub0/c15 ),
    .fx({\PWMD/n12 [14],\PWMD/n12 [12]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWMD/sub0/ucin_al_u3454"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWMD/sub0/u15_al_u3458  (
    .a({\PWMD/FreCnt [17],\PWMD/FreCnt [15]}),
    .b({\PWMD/FreCnt [18],\PWMD/FreCnt [16]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWMD/sub0/c15 ),
    .f({\PWMD/n12 [17],\PWMD/n12 [15]}),
    .fco(\PWMD/sub0/c19 ),
    .fx({\PWMD/n12 [18],\PWMD/n12 [16]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWMD/sub0/ucin_al_u3454"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWMD/sub0/u19_al_u3459  (
    .a({\PWMD/FreCnt [21],\PWMD/FreCnt [19]}),
    .b({\PWMD/FreCnt [22],\PWMD/FreCnt [20]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWMD/sub0/c19 ),
    .f({\PWMD/n12 [21],\PWMD/n12 [19]}),
    .fco(\PWMD/sub0/c23 ),
    .fx({\PWMD/n12 [22],\PWMD/n12 [20]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWMD/sub0/ucin_al_u3454"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWMD/sub0/u23_al_u3460  (
    .a({\PWMD/FreCnt [25],\PWMD/FreCnt [23]}),
    .b({\PWMD/FreCnt [26],\PWMD/FreCnt [24]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWMD/sub0/c23 ),
    .f({\PWMD/n12 [25],\PWMD/n12 [23]}),
    .fx({\PWMD/n12 [26],\PWMD/n12 [24]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWMD/sub0/ucin_al_u3454"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWMD/sub0/u3_al_u3455  (
    .a({\PWMD/FreCnt [5],\PWMD/FreCnt [3]}),
    .b({\PWMD/FreCnt [6],\PWMD/FreCnt [4]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWMD/sub0/c3 ),
    .f({\PWMD/n12 [5],\PWMD/n12 [3]}),
    .fco(\PWMD/sub0/c7 ),
    .fx({\PWMD/n12 [6],\PWMD/n12 [4]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWMD/sub0/ucin_al_u3454"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWMD/sub0/u7_al_u3456  (
    .a({\PWMD/FreCnt [9],\PWMD/FreCnt [7]}),
    .b({\PWMD/FreCnt [10],\PWMD/FreCnt [8]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWMD/sub0/c7 ),
    .f({\PWMD/n12 [9],\PWMD/n12 [7]}),
    .fco(\PWMD/sub0/c11 ),
    .fx({\PWMD/n12 [10],\PWMD/n12 [8]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWMD/sub0/ucin_al_u3454"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h0005),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWMD/sub0/ucin_al_u3454  (
    .a({\PWMD/FreCnt [1],1'b0}),
    .b({\PWMD/FreCnt [2],\PWMD/FreCnt [0]}),
    .c(2'b11),
    .d(2'b01),
    .e(2'b01),
    .f({\PWMD/n12 [1],open_n22829}),
    .fco(\PWMD/sub0/c3 ),
    .fx({\PWMD/n12 [2],\PWMD/n12 [0]}));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMD/sub1/u0|PWMD/sub1/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("SUB_CARRY"),
    .INIT_LUT0(16'b0000000000000101),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMD/sub1/u0|PWMD/sub1/ucin  (
    .a({pnumcntD[0],1'b0}),
    .b({1'b1,open_n22832}),
    .f({\PWMD/n26 [0],open_n22852}),
    .fco(\PWMD/sub1/c1 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMD/sub1/u0|PWMD/sub1/ucin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMD/sub1/u10|PWMD/sub1/u9  (
    .a(pnumcntD[10:9]),
    .b(2'b00),
    .fci(\PWMD/sub1/c9 ),
    .f(\PWMD/n26 [10:9]),
    .fco(\PWMD/sub1/c11 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMD/sub1/u0|PWMD/sub1/ucin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMD/sub1/u12|PWMD/sub1/u11  (
    .a(pnumcntD[12:11]),
    .b(2'b00),
    .fci(\PWMD/sub1/c11 ),
    .f(\PWMD/n26 [12:11]),
    .fco(\PWMD/sub1/c13 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMD/sub1/u0|PWMD/sub1/ucin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMD/sub1/u14|PWMD/sub1/u13  (
    .a(pnumcntD[14:13]),
    .b(2'b00),
    .fci(\PWMD/sub1/c13 ),
    .f(\PWMD/n26 [14:13]),
    .fco(\PWMD/sub1/c15 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMD/sub1/u0|PWMD/sub1/ucin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMD/sub1/u16|PWMD/sub1/u15  (
    .a(pnumcntD[16:15]),
    .b(2'b00),
    .fci(\PWMD/sub1/c15 ),
    .f(\PWMD/n26 [16:15]),
    .fco(\PWMD/sub1/c17 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMD/sub1/u0|PWMD/sub1/ucin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMD/sub1/u18|PWMD/sub1/u17  (
    .a(pnumcntD[18:17]),
    .b(2'b00),
    .fci(\PWMD/sub1/c17 ),
    .f(\PWMD/n26 [18:17]),
    .fco(\PWMD/sub1/c19 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMD/sub1/u0|PWMD/sub1/ucin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMD/sub1/u20|PWMD/sub1/u19  (
    .a(pnumcntD[20:19]),
    .b(2'b00),
    .fci(\PWMD/sub1/c19 ),
    .f(\PWMD/n26 [20:19]),
    .fco(\PWMD/sub1/c21 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMD/sub1/u0|PWMD/sub1/ucin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMD/sub1/u22|PWMD/sub1/u21  (
    .a(pnumcntD[22:21]),
    .b(2'b00),
    .fci(\PWMD/sub1/c21 ),
    .f(\PWMD/n26 [22:21]),
    .fco(\PWMD/sub1/c23 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMD/sub1/u0|PWMD/sub1/ucin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMD/sub1/u23_al_u3481  (
    .a({open_n23011,pnumcntD[23]}),
    .b({open_n23012,1'b0}),
    .fci(\PWMD/sub1/c23 ),
    .f({open_n23031,\PWMD/n26 [23]}));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMD/sub1/u0|PWMD/sub1/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMD/sub1/u2|PWMD/sub1/u1  (
    .a(pnumcntD[2:1]),
    .b(2'b00),
    .fci(\PWMD/sub1/c1 ),
    .f(\PWMD/n26 [2:1]),
    .fco(\PWMD/sub1/c3 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMD/sub1/u0|PWMD/sub1/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMD/sub1/u4|PWMD/sub1/u3  (
    .a(pnumcntD[4:3]),
    .b(2'b00),
    .fci(\PWMD/sub1/c3 ),
    .f(\PWMD/n26 [4:3]),
    .fco(\PWMD/sub1/c5 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMD/sub1/u0|PWMD/sub1/ucin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMD/sub1/u6|PWMD/sub1/u5  (
    .a(pnumcntD[6:5]),
    .b(2'b00),
    .fci(\PWMD/sub1/c5 ),
    .f(\PWMD/n26 [6:5]),
    .fco(\PWMD/sub1/c7 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMD/sub1/u0|PWMD/sub1/ucin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMD/sub1/u8|PWMD/sub1/u7  (
    .a(pnumcntD[8:7]),
    .b(2'b00),
    .fci(\PWMD/sub1/c7 ),
    .f(\PWMD/n26 [8:7]),
    .fco(\PWMD/sub1/c9 ));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[0]  (
    .i(\PWME/RemaTxNum[0]_keep ),
    .o(pnumcntE[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[10]  (
    .i(\PWME/RemaTxNum[10]_keep ),
    .o(pnumcntE[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[11]  (
    .i(\PWME/RemaTxNum[11]_keep ),
    .o(pnumcntE[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[12]  (
    .i(\PWME/RemaTxNum[12]_keep ),
    .o(pnumcntE[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[13]  (
    .i(\PWME/RemaTxNum[13]_keep ),
    .o(pnumcntE[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[14]  (
    .i(\PWME/RemaTxNum[14]_keep ),
    .o(pnumcntE[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[15]  (
    .i(\PWME/RemaTxNum[15]_keep ),
    .o(pnumcntE[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[16]  (
    .i(\PWME/RemaTxNum[16]_keep ),
    .o(pnumcntE[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[17]  (
    .i(\PWME/RemaTxNum[17]_keep ),
    .o(pnumcntE[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[18]  (
    .i(\PWME/RemaTxNum[18]_keep ),
    .o(pnumcntE[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[19]  (
    .i(\PWME/RemaTxNum[19]_keep ),
    .o(pnumcntE[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[1]  (
    .i(\PWME/RemaTxNum[1]_keep ),
    .o(pnumcntE[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[20]  (
    .i(\PWME/RemaTxNum[20]_keep ),
    .o(pnumcntE[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[21]  (
    .i(\PWME/RemaTxNum[21]_keep ),
    .o(pnumcntE[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[22]  (
    .i(\PWME/RemaTxNum[22]_keep ),
    .o(pnumcntE[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[23]  (
    .i(\PWME/RemaTxNum[23]_keep ),
    .o(pnumcntE[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[2]  (
    .i(\PWME/RemaTxNum[2]_keep ),
    .o(pnumcntE[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[3]  (
    .i(\PWME/RemaTxNum[3]_keep ),
    .o(pnumcntE[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[4]  (
    .i(\PWME/RemaTxNum[4]_keep ),
    .o(pnumcntE[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[5]  (
    .i(\PWME/RemaTxNum[5]_keep ),
    .o(pnumcntE[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[6]  (
    .i(\PWME/RemaTxNum[6]_keep ),
    .o(pnumcntE[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[7]  (
    .i(\PWME/RemaTxNum[7]_keep ),
    .o(pnumcntE[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[8]  (
    .i(\PWME/RemaTxNum[8]_keep ),
    .o(pnumcntE[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[9]  (
    .i(\PWME/RemaTxNum[9]_keep ),
    .o(pnumcntE[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_dir  (
    .i(\PWME/dir_keep ),
    .o(dir_pad[14]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[0]  (
    .i(\PWME/pnumr[0]_keep ),
    .o(\PWME/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[10]  (
    .i(\PWME/pnumr[10]_keep ),
    .o(\PWME/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[11]  (
    .i(\PWME/pnumr[11]_keep ),
    .o(\PWME/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[12]  (
    .i(\PWME/pnumr[12]_keep ),
    .o(\PWME/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[13]  (
    .i(\PWME/pnumr[13]_keep ),
    .o(\PWME/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[14]  (
    .i(\PWME/pnumr[14]_keep ),
    .o(\PWME/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[15]  (
    .i(\PWME/pnumr[15]_keep ),
    .o(\PWME/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[16]  (
    .i(\PWME/pnumr[16]_keep ),
    .o(\PWME/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[17]  (
    .i(\PWME/pnumr[17]_keep ),
    .o(\PWME/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[18]  (
    .i(\PWME/pnumr[18]_keep ),
    .o(\PWME/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[19]  (
    .i(\PWME/pnumr[19]_keep ),
    .o(\PWME/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[1]  (
    .i(\PWME/pnumr[1]_keep ),
    .o(\PWME/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[20]  (
    .i(\PWME/pnumr[20]_keep ),
    .o(\PWME/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[21]  (
    .i(\PWME/pnumr[21]_keep ),
    .o(\PWME/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[22]  (
    .i(\PWME/pnumr[22]_keep ),
    .o(\PWME/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[23]  (
    .i(\PWME/pnumr[23]_keep ),
    .o(\PWME/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[24]  (
    .i(\PWME/pnumr[24]_keep ),
    .o(\PWME/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[25]  (
    .i(\PWME/pnumr[25]_keep ),
    .o(\PWME/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[26]  (
    .i(\PWME/pnumr[26]_keep ),
    .o(\PWME/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[27]  (
    .i(\PWME/pnumr[27]_keep ),
    .o(\PWME/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[28]  (
    .i(\PWME/pnumr[28]_keep ),
    .o(\PWME/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[29]  (
    .i(\PWME/pnumr[29]_keep ),
    .o(\PWME/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[2]  (
    .i(\PWME/pnumr[2]_keep ),
    .o(\PWME/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[30]  (
    .i(\PWME/pnumr[30]_keep ),
    .o(\PWME/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[31]  (
    .i(\PWME/pnumr[31]_keep ),
    .o(\PWME/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[3]  (
    .i(\PWME/pnumr[3]_keep ),
    .o(\PWME/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[4]  (
    .i(\PWME/pnumr[4]_keep ),
    .o(\PWME/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[5]  (
    .i(\PWME/pnumr[5]_keep ),
    .o(\PWME/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[6]  (
    .i(\PWME/pnumr[6]_keep ),
    .o(\PWME/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[7]  (
    .i(\PWME/pnumr[7]_keep ),
    .o(\PWME/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[8]  (
    .i(\PWME/pnumr[8]_keep ),
    .o(\PWME/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[9]  (
    .i(\PWME/pnumr[9]_keep ),
    .o(\PWME/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pwm  (
    .i(\PWME/pwm_keep ),
    .o(pwm_pad[14]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_stopreq  (
    .i(\PWME/stopreq_keep ),
    .o(\PWME/stopreq ));  // src/OnePWM.v(14)
  EF2_PHY_MSLICE #(
    //.LUT0("(D*~(C)*~((~0*~(B*A)))+D*C*~((~0*~(B*A)))+~(D)*C*(~0*~(B*A))+D*C*(~0*~(B*A)))"),
    //.LUT1("(D*~(C)*~((~1*~(B*A)))+D*C*~((~1*~(B*A)))+~(D)*C*(~1*~(B*A))+D*C*(~1*~(B*A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111100001110000),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/dir_reg  (
    .a({\PWME/n24 ,\PWME/n24 }),
    .b({\PWME/n25_neg_lutinv ,\PWME/n25_neg_lutinv }),
    .c({dir_pad[14],dir_pad[14]}),
    .clk(clk100m),
    .d({\PWME/pnumr [31],\PWME/pnumr [31]}),
    .mi({open_n23136,pwm_start_stop[30]}),
    .q({open_n23143,\PWME/dir_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("~(~0*~(D*C*B*A))"),
    //.LUT1("~(~1*~(D*C*B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b1111111111111111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWME/pwm_reg  (
    .a({_al_u1607_o,_al_u1607_o}),
    .b({_al_u1614_o,_al_u1614_o}),
    .c({_al_u1616_o,_al_u1616_o}),
    .clk(clk100m),
    .d({_al_u1618_o,_al_u1618_o}),
    .mi({open_n23155,pwm_pad[14]}),
    .sr(\PWME/u14_sel_is_1_o ),
    .q({open_n23161,\PWME/pwm_keep }));  // src/OnePWM.v(45)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWME/reg0_b0|PWME/reg0_b5  (
    .b({\PWME/n12 [0],\PWME/n12 [5]}),
    .c({freqE[0],freqE[5]}),
    .clk(clk100m),
    .d({\PWME/n0_lutinv ,\PWME/n0_lutinv }),
    .sr(\PWME/n11 ),
    .q({\PWME/FreCnt [0],\PWME/FreCnt [5]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWME/reg0_b10|PWME/reg0_b3  (
    .b({\PWME/n12 [10],\PWME/n12 [3]}),
    .c({freqE[10],freqE[3]}),
    .clk(clk100m),
    .d({\PWME/n0_lutinv ,\PWME/n0_lutinv }),
    .sr(\PWME/n11 ),
    .q({\PWME/FreCnt [10],\PWME/FreCnt [3]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWME/reg0_b11|PWME/reg0_b23  (
    .b({\PWME/n12 [11],\PWME/n12 [23]}),
    .c({freqE[11],freqE[23]}),
    .clk(clk100m),
    .d({\PWME/n0_lutinv ,\PWME/n0_lutinv }),
    .sr(\PWME/n11 ),
    .q({\PWME/FreCnt [11],\PWME/FreCnt [23]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWME/reg0_b14|PWME/reg0_b12  (
    .b({\PWME/n12 [14],\PWME/n12 [12]}),
    .c({freqE[14],freqE[12]}),
    .clk(clk100m),
    .d({\PWME/n0_lutinv ,\PWME/n0_lutinv }),
    .sr(\PWME/n11 ),
    .q({\PWME/FreCnt [14],\PWME/FreCnt [12]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWME/reg0_b16|PWME/reg0_b9  (
    .b({\PWME/n12 [16],\PWME/n12 [9]}),
    .c({freqE[16],freqE[9]}),
    .clk(clk100m),
    .d({\PWME/n0_lutinv ,\PWME/n0_lutinv }),
    .sr(\PWME/n11 ),
    .q({\PWME/FreCnt [16],\PWME/FreCnt [9]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWME/reg0_b18|PWME/reg0_b8  (
    .b({\PWME/n12 [18],\PWME/n12 [8]}),
    .c({freqE[18],freqE[8]}),
    .clk(clk100m),
    .d({\PWME/n0_lutinv ,\PWME/n0_lutinv }),
    .sr(\PWME/n11 ),
    .q({\PWME/FreCnt [18],\PWME/FreCnt [8]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWME/reg0_b20|PWME/reg0_b7  (
    .b({\PWME/n12 [20],\PWME/n12 [7]}),
    .c({freqE[20],freqE[7]}),
    .clk(clk100m),
    .d({\PWME/n0_lutinv ,\PWME/n0_lutinv }),
    .sr(\PWME/n11 ),
    .q({\PWME/FreCnt [20],\PWME/FreCnt [7]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWME/reg0_b22|PWME/reg0_b6  (
    .b({\PWME/n12 [22],\PWME/n12 [6]}),
    .c({freqE[22],freqE[6]}),
    .clk(clk100m),
    .d({\PWME/n0_lutinv ,\PWME/n0_lutinv }),
    .sr(\PWME/n11 ),
    .q({\PWME/FreCnt [22],\PWME/FreCnt [6]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWME/reg0_b24|PWME/reg0_b4  (
    .b({\PWME/n12 [24],\PWME/n12 [4]}),
    .c({freqE[24],freqE[4]}),
    .clk(clk100m),
    .d({\PWME/n0_lutinv ,\PWME/n0_lutinv }),
    .sr(\PWME/n11 ),
    .q({\PWME/FreCnt [24],\PWME/FreCnt [4]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWME/reg0_b25|PWME/reg0_b26  (
    .b({\PWME/n12 [25],\PWME/n12 [26]}),
    .c({freqE[25],freqE[26]}),
    .clk(clk100m),
    .d({\PWME/n0_lutinv ,\PWME/n0_lutinv }),
    .sr(\PWME/n11 ),
    .q({\PWME/FreCnt [25],\PWME/FreCnt [26]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~A*~(0@C)*~(~D*B))"),
    //.LUTF1("(~A*~(~0*C)*~(D@B))"),
    //.LUTG0("(~A*~(1@C)*~(~D*B))"),
    //.LUTG1("(~A*~(~1*C)*~(D@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010100000001),
    .INIT_LUTF1(16'b0000010000000001),
    .INIT_LUTG0(16'b0101000000010000),
    .INIT_LUTG1(16'b0100010000010001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/reg1_b13|PWME/reg1_b24  (
    .a({_al_u2875_o,_al_u1611_o}),
    .b({\PWME/FreCnt [12],\PWME/FreCnt [12]}),
    .c({\PWME/FreCnt [23],\PWME/FreCnt [24]}),
    .ce(\PWME/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d(\PWME/FreCntr [13:12]),
    .e({\PWME/FreCntr [24],\PWME/FreCntr [24]}),
    .mi({freqE[13],freqE[24]}),
    .f({_al_u2876_o,_al_u1612_o}),
    .q({\PWME/FreCntr [13],\PWME/FreCntr [24]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(~(~D*B)*~(~C*A))"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(~(~D*B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b1111010100110001),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b1111010100110001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/reg1_b15|PWME/reg1_b26  (
    .a({\PWME/FreCnt [1],open_n23398}),
    .b({\PWME/FreCnt [15],_al_u1256_o}),
    .c({\PWME/FreCntr [1],_al_u1258_o}),
    .ce(\PWME/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWME/FreCntr [15],_al_u1254_o}),
    .mi({freqE[15],freqE[26]}),
    .f({_al_u1613_o,\PWME/n0_lutinv }),
    .q({\PWME/FreCntr [15],\PWME/FreCntr [26]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*~C)*~(~D*B))"),
    //.LUTF1("(~(C*~B)*~(D*~A))"),
    //.LUTG0("(A*~(1*~C)*~(~D*B))"),
    //.LUTG1("(~(C*~B)*~(D*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101000100010),
    .INIT_LUTF1(16'b1000101011001111),
    .INIT_LUTG0(16'b1010000000100000),
    .INIT_LUTG1(16'b1000101011001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/reg1_b16|PWME/reg1_b2  (
    .a({\PWME/FreCnt [1],_al_u2893_o}),
    .b({\PWME/FreCnt [15],\PWME/FreCnt [1]}),
    .c({\PWME/FreCntr [16],\PWME/FreCnt [19]}),
    .ce(\PWME/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWME/FreCntr [2],\PWME/FreCntr [2]}),
    .e({open_n23417,\PWME/FreCntr [20]}),
    .mi({freqE[16],freqE[2]}),
    .f({_al_u2885_o,_al_u2894_o}),
    .q({\PWME/FreCntr [16],\PWME/FreCntr [2]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~A*~(0@C)*~(D*~B))"),
    //.LUTF1("(B*A*~(D@C))"),
    //.LUTG0("(~A*~(1@C)*~(D*~B))"),
    //.LUTG1("(B*A*~(D@C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010000000101),
    .INIT_LUTF1(16'b1000000000001000),
    .INIT_LUTG0(16'b0100000001010000),
    .INIT_LUTG1(16'b1000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/reg1_b17|PWME/reg1_b9  (
    .a({_al_u2882_o,_al_u2881_o}),
    .b({_al_u2883_o,\PWME/FreCnt [21]}),
    .c({\PWME/FreCnt [16],\PWME/FreCnt [8]}),
    .ce(\PWME/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWME/FreCntr [17],\PWME/FreCntr [22]}),
    .e({open_n23434,\PWME/FreCntr [9]}),
    .mi({freqE[17],freqE[9]}),
    .f({_al_u2884_o,_al_u2882_o}),
    .q({\PWME/FreCntr [17],\PWME/FreCntr [9]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~B*~(0@C)*~(~D*A))"),
    //.LUTF1("(~(~D*B)*~(C*~A))"),
    //.LUTG0("(~B*~(1@C)*~(~D*A))"),
    //.LUTG1("(~(~D*B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000001100000001),
    .INIT_LUTF1(16'b1010111100100011),
    .INIT_LUTG0(16'b0011000000010000),
    .INIT_LUTG1(16'b1010111100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/reg1_b22|PWME/reg1_b14  (
    .a({\PWME/FreCnt [13],\PWME/FreCnt [13]}),
    .b({\PWME/FreCnt [21],\PWME/FreCnt [26]}),
    .c({\PWME/FreCntr [14],\PWME/FreCnt [7]}),
    .ce(\PWME/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWME/FreCntr [22],\PWME/FreCntr [14]}),
    .e({open_n23451,\PWME/FreCntr [8]}),
    .mi({freqE[22],freqE[14]}),
    .f({_al_u2887_o,_al_u2895_o}),
    .q({\PWME/FreCntr [22],\PWME/FreCntr [14]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(~0*C)*~(D*~B))"),
    //.LUTF1("(A*~(0@C)*~(~D*B))"),
    //.LUTG0("(A*~(~1*C)*~(D*~B))"),
    //.LUTG1("(A*~(1@C)*~(~D*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000001010),
    .INIT_LUTF1(16'b0000101000000010),
    .INIT_LUTG0(16'b1000100010101010),
    .INIT_LUTG1(16'b1010000000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/reg1_b25|PWME/reg1_b11  (
    .a({_al_u2876_o,_al_u2885_o}),
    .b({\PWME/FreCnt [10],\PWME/FreCnt [10]}),
    .c({\PWME/FreCnt [24],\PWME/FreCnt [19]}),
    .ce(\PWME/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWME/FreCntr [11],\PWME/FreCntr [11]}),
    .e({\PWME/FreCntr [25],\PWME/FreCntr [20]}),
    .mi({freqE[25],freqE[11]}),
    .f({_al_u2877_o,_al_u2886_o}),
    .q({\PWME/FreCntr [25],\PWME/FreCntr [11]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*B*A*~(0@D))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(C*B*A*~(1@D))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/reg1_b3|PWME/reg1_b10  (
    .a({\PWME/FreCnt [10],_al_u2877_o}),
    .b({\PWME/FreCnt [3],_al_u2878_o}),
    .c({\PWME/FreCntr [10],_al_u2879_o}),
    .ce(\PWME/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWME/FreCntr [3],\PWME/FreCnt [9]}),
    .e({open_n23484,\PWME/FreCntr [10]}),
    .mi({freqE[3],freqE[10]}),
    .f({_al_u1609_o,_al_u2880_o}),
    .q({\PWME/FreCntr [3],\PWME/FreCntr [10]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(D*~B)*~(~C*A))"),
    //.LUT1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100010011110101),
    .INIT_LUT1(16'b1000010000100001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/reg1_b5|PWME/reg1_b18  (
    .a(\PWME/FreCnt [18:17]),
    .b({\PWME/FreCnt [5],\PWME/FreCnt [23]}),
    .c({\PWME/FreCntr [18],\PWME/FreCntr [18]}),
    .ce(\PWME/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWME/FreCntr [5],\PWME/FreCntr [24]}),
    .mi({freqE[5],freqE[18]}),
    .f({_al_u1606_o,_al_u2893_o}),
    .q({\PWME/FreCntr [5],\PWME/FreCntr [18]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~D*B)*~(~C*A))"),
    //.LUTF1("(~(~D*B)*~(C*~A))"),
    //.LUTG0("(~(~D*B)*~(~C*A))"),
    //.LUTG1("(~(~D*B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111010100110001),
    .INIT_LUTF1(16'b1010111100100011),
    .INIT_LUTG0(16'b1111010100110001),
    .INIT_LUTG1(16'b1010111100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/reg1_b6|PWME/reg1_b4  (
    .a({\PWME/FreCnt [3],\PWME/FreCnt [15]}),
    .b({\PWME/FreCnt [5],\PWME/FreCnt [3]}),
    .c({\PWME/FreCntr [4],\PWME/FreCntr [16]}),
    .ce(\PWME/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWME/FreCntr [6],\PWME/FreCntr [4]}),
    .mi({freqE[6],freqE[4]}),
    .f({_al_u2878_o,_al_u2883_o}),
    .q({\PWME/FreCntr [6],\PWME/FreCntr [4]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(D@B)*~(C@A))"),
    //.LUTF1("(D*~(C@B))"),
    //.LUTG0("(~(D@B)*~(C@A))"),
    //.LUTG1("(D*~(C@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000010000100001),
    .INIT_LUTF1(16'b1100001100000000),
    .INIT_LUTG0(16'b1000010000100001),
    .INIT_LUTG1(16'b1100001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/reg1_b7|PWME/reg1_b23  (
    .a({open_n23533,\PWME/FreCnt [22]}),
    .b({\PWME/FreCnt [6],\PWME/FreCnt [4]}),
    .c({\PWME/FreCntr [7],\PWME/FreCntr [23]}),
    .ce(\PWME/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({_al_u2889_o,\PWME/FreCntr [5]}),
    .mi({freqE[7],freqE[23]}),
    .f({_al_u2890_o,_al_u2889_o}),
    .q({\PWME/FreCntr [7],\PWME/FreCntr [23]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011100010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/reg2_b0|PWME/reg2_b7  (
    .a({\PWME/pnumr [0],\PWME/pnumr [7]}),
    .b({pnumE[0],pnumE[32]}),
    .c({pnumE[32],pnumE[7]}),
    .clk(clk100m),
    .d({pwm_start_stop[30],pwm_start_stop[30]}),
    .q({\PWME/pnumr[0]_keep ,\PWME/pnumr[7]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/reg2_b10|PWME/reg3_b10  (
    .a({\PWME/pnumr [10],_al_u2869_o}),
    .b({pnumE[10],\PWME/n24 }),
    .c({pnumE[32],pnumcntE[10]}),
    .clk(clk100m),
    .d({pwm_start_stop[30],\PWME/pnumr [10]}),
    .e({open_n23572,pwm_start_stop[30]}),
    .q({\PWME/pnumr[10]_keep ,\PWME/RemaTxNum[10]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/reg2_b11|PWME/reg3_b11  (
    .a({\PWME/pnumr [11],_al_u2867_o}),
    .b({pnumE[11],\PWME/n24 }),
    .c({pnumE[32],pnumcntE[11]}),
    .clk(clk100m),
    .d({pwm_start_stop[30],\PWME/pnumr [11]}),
    .e({open_n23594,pwm_start_stop[30]}),
    .q({\PWME/pnumr[11]_keep ,\PWME/RemaTxNum[11]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011100010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/reg2_b12|PWME/reg2_b6  (
    .a({\PWME/pnumr [12],\PWME/pnumr [6]}),
    .b({pnumE[12],pnumE[32]}),
    .c({pnumE[32],pnumE[6]}),
    .clk(clk100m),
    .d({pwm_start_stop[30],pwm_start_stop[30]}),
    .q({\PWME/pnumr[12]_keep ,\PWME/pnumr[6]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/reg2_b13|PWME/reg2_b3  (
    .a({\PWME/pnumr [13],\PWME/pnumr [3]}),
    .b({pnumE[13],pnumE[3]}),
    .c({pnumE[32],pnumE[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[30],pwm_start_stop[30]}),
    .q({\PWME/pnumr[13]_keep ,\PWME/pnumr[3]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/reg2_b14|PWME/reg3_b14  (
    .a({\PWME/pnumr [14],_al_u2861_o}),
    .b({pnumE[14],\PWME/n24 }),
    .c({pnumE[32],pnumcntE[14]}),
    .clk(clk100m),
    .d({pwm_start_stop[30],\PWME/pnumr [14]}),
    .e({open_n23658,pwm_start_stop[30]}),
    .q({\PWME/pnumr[14]_keep ,\PWME/RemaTxNum[14]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/reg2_b15|PWME/reg3_b15  (
    .a({\PWME/pnumr [15],_al_u2859_o}),
    .b({pnumE[15],\PWME/n24 }),
    .c({pnumE[32],pnumcntE[15]}),
    .clk(clk100m),
    .d({pwm_start_stop[30],\PWME/pnumr [15]}),
    .e({open_n23680,pwm_start_stop[30]}),
    .q({\PWME/pnumr[15]_keep ,\PWME/RemaTxNum[15]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/reg2_b16|PWME/reg2_b23  (
    .a({\PWME/pnumr [16],\PWME/pnumr [23]}),
    .b({pnumE[16],pnumE[23]}),
    .c({pnumE[32],pnumE[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[30],pwm_start_stop[30]}),
    .q({\PWME/pnumr[16]_keep ,\PWME/pnumr[23]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/reg2_b17|PWME/reg2_b20  (
    .a({\PWME/pnumr [17],\PWME/pnumr [20]}),
    .b({pnumE[17],pnumE[20]}),
    .c({pnumE[32],pnumE[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[30],pwm_start_stop[30]}),
    .q({\PWME/pnumr[17]_keep ,\PWME/pnumr[20]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/reg2_b18|PWME/reg3_b18  (
    .a({\PWME/pnumr [18],_al_u2853_o}),
    .b({pnumE[18],\PWME/n24 }),
    .c({pnumE[32],pnumcntE[18]}),
    .clk(clk100m),
    .d({pwm_start_stop[30],\PWME/pnumr [18]}),
    .e({open_n23744,pwm_start_stop[30]}),
    .q({\PWME/pnumr[18]_keep ,\PWME/RemaTxNum[18]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/reg2_b19|PWME/reg3_b19  (
    .a({\PWME/pnumr [19],_al_u2851_o}),
    .b({pnumE[19],\PWME/n24 }),
    .c({pnumE[32],pnumcntE[19]}),
    .clk(clk100m),
    .d({pwm_start_stop[30],\PWME/pnumr [19]}),
    .e({open_n23766,pwm_start_stop[30]}),
    .q({\PWME/pnumr[19]_keep ,\PWME/RemaTxNum[19]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/reg2_b1|PWME/reg2_b2  (
    .a({\PWME/pnumr [1],\PWME/pnumr [2]}),
    .b({pnumE[1],pnumE[2]}),
    .c({pnumE[32],pnumE[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[30],pwm_start_stop[30]}),
    .q({\PWME/pnumr[1]_keep ,\PWME/pnumr[2]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/reg2_b21|PWME/reg3_b21  (
    .a({\PWME/pnumr [21],_al_u2845_o}),
    .b({pnumE[21],\PWME/n24 }),
    .c({pnumE[32],pnumcntE[21]}),
    .clk(clk100m),
    .d({pwm_start_stop[30],\PWME/pnumr [21]}),
    .e({open_n23807,pwm_start_stop[30]}),
    .q({\PWME/pnumr[21]_keep ,\PWME/RemaTxNum[21]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/reg2_b22|PWME/reg3_b22  (
    .a({\PWME/pnumr [22],_al_u2843_o}),
    .b({pnumE[22],\PWME/n24 }),
    .c({pnumE[32],pnumcntE[22]}),
    .clk(clk100m),
    .d({pwm_start_stop[30],\PWME/pnumr [22]}),
    .e({open_n23829,pwm_start_stop[30]}),
    .q({\PWME/pnumr[22]_keep ,\PWME/RemaTxNum[22]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/reg2_b24|PWME/reg2_b31  (
    .a({\PWME/pnumr [24],\PWME/pnumr [31]}),
    .b({pnumE[24],pnumE[31]}),
    .c({pnumE[32],pnumE[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[30],pwm_start_stop[30]}),
    .q({\PWME/pnumr[24]_keep ,\PWME/pnumr[31]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/reg2_b25|PWME/reg2_b30  (
    .a({\PWME/pnumr [25],\PWME/pnumr [30]}),
    .b({pnumE[25],pnumE[30]}),
    .c({pnumE[32],pnumE[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[30],pwm_start_stop[30]}),
    .q({\PWME/pnumr[25]_keep ,\PWME/pnumr[30]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/reg2_b26|PWME/reg2_b29  (
    .a({\PWME/pnumr [26],\PWME/pnumr [29]}),
    .b({pnumE[26],pnumE[29]}),
    .c({pnumE[32],pnumE[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[30],pwm_start_stop[30]}),
    .q({\PWME/pnumr[26]_keep ,\PWME/pnumr[29]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/reg2_b27|PWME/reg2_b28  (
    .a({\PWME/pnumr [27],\PWME/pnumr [28]}),
    .b({pnumE[27],pnumE[28]}),
    .c({pnumE[32],pnumE[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[30],pwm_start_stop[30]}),
    .q({\PWME/pnumr[27]_keep ,\PWME/pnumr[28]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/reg2_b4|PWME/reg3_b4  (
    .a({\PWME/pnumr [4],_al_u2837_o}),
    .b({pnumE[32],\PWME/n24 }),
    .c({pnumE[4],pnumcntE[4]}),
    .clk(clk100m),
    .d({pwm_start_stop[30],\PWME/pnumr [4]}),
    .e({open_n23931,pwm_start_stop[30]}),
    .q({\PWME/pnumr[4]_keep ,\PWME/RemaTxNum[4]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/reg2_b5|PWME/reg3_b5  (
    .a({\PWME/pnumr [5],_al_u2835_o}),
    .b({pnumE[32],\PWME/n24 }),
    .c({pnumE[5],pnumcntE[5]}),
    .clk(clk100m),
    .d({pwm_start_stop[30],\PWME/pnumr [5]}),
    .e({open_n23953,pwm_start_stop[30]}),
    .q({\PWME/pnumr[5]_keep ,\PWME/RemaTxNum[5]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/reg2_b8|PWME/reg3_b8  (
    .a({\PWME/pnumr [8],_al_u2829_o}),
    .b({pnumE[32],\PWME/n24 }),
    .c({pnumE[8],pnumcntE[8]}),
    .clk(clk100m),
    .d({pwm_start_stop[30],\PWME/pnumr [8]}),
    .e({open_n23975,pwm_start_stop[30]}),
    .q({\PWME/pnumr[8]_keep ,\PWME/RemaTxNum[8]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/reg2_b9|PWME/reg3_b9  (
    .a({\PWME/pnumr [9],_al_u2827_o}),
    .b({pnumE[32],\PWME/n24 }),
    .c({pnumE[9],pnumcntE[9]}),
    .clk(clk100m),
    .d({pwm_start_stop[30],\PWME/pnumr [9]}),
    .e({open_n23997,pwm_start_stop[30]}),
    .q({\PWME/pnumr[9]_keep ,\PWME/RemaTxNum[9]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/reg3_b0  (
    .a({_al_u2873_o,_al_u2873_o}),
    .b({\PWME/n24 ,\PWME/n24 }),
    .c({pnumcntE[0],pnumcntE[0]}),
    .clk(clk100m),
    .d({\PWME/pnumr [0],\PWME/pnumr [0]}),
    .mi({open_n24029,pwm_start_stop[30]}),
    .q({open_n24036,\PWME/RemaTxNum[0]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/reg3_b1  (
    .a({_al_u2871_o,_al_u2871_o}),
    .b({\PWME/n24 ,\PWME/n24 }),
    .c({pnumcntE[1],pnumcntE[1]}),
    .clk(clk100m),
    .d({\PWME/pnumr [1],\PWME/pnumr [1]}),
    .mi({open_n24048,pwm_start_stop[30]}),
    .q({open_n24055,\PWME/RemaTxNum[1]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/reg3_b12  (
    .a({_al_u2865_o,_al_u2865_o}),
    .b({\PWME/n24 ,\PWME/n24 }),
    .c({pnumcntE[12],pnumcntE[12]}),
    .clk(clk100m),
    .d({\PWME/pnumr [12],\PWME/pnumr [12]}),
    .mi({open_n24067,pwm_start_stop[30]}),
    .q({open_n24074,\PWME/RemaTxNum[12]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/reg3_b13  (
    .a({_al_u2863_o,_al_u2863_o}),
    .b({\PWME/n24 ,\PWME/n24 }),
    .c({pnumcntE[13],pnumcntE[13]}),
    .clk(clk100m),
    .d({\PWME/pnumr [13],\PWME/pnumr [13]}),
    .mi({open_n24086,pwm_start_stop[30]}),
    .q({open_n24093,\PWME/RemaTxNum[13]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/reg3_b16  (
    .a({_al_u2857_o,_al_u2857_o}),
    .b({\PWME/n24 ,\PWME/n24 }),
    .c({pnumcntE[16],pnumcntE[16]}),
    .clk(clk100m),
    .d({\PWME/pnumr [16],\PWME/pnumr [16]}),
    .mi({open_n24105,pwm_start_stop[30]}),
    .q({open_n24112,\PWME/RemaTxNum[16]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/reg3_b17  (
    .a({_al_u2855_o,_al_u2855_o}),
    .b({\PWME/n24 ,\PWME/n24 }),
    .c({pnumcntE[17],pnumcntE[17]}),
    .clk(clk100m),
    .d({\PWME/pnumr [17],\PWME/pnumr [17]}),
    .mi({open_n24124,pwm_start_stop[30]}),
    .q({open_n24131,\PWME/RemaTxNum[17]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/reg3_b2  (
    .a({_al_u2849_o,_al_u2849_o}),
    .b({\PWME/n24 ,\PWME/n24 }),
    .c({pnumcntE[2],pnumcntE[2]}),
    .clk(clk100m),
    .d({\PWME/pnumr [2],\PWME/pnumr [2]}),
    .mi({open_n24143,pwm_start_stop[30]}),
    .q({open_n24150,\PWME/RemaTxNum[2]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/reg3_b20  (
    .a({_al_u2847_o,_al_u2847_o}),
    .b({\PWME/n24 ,\PWME/n24 }),
    .c({pnumcntE[20],pnumcntE[20]}),
    .clk(clk100m),
    .d({\PWME/pnumr [20],\PWME/pnumr [20]}),
    .mi({open_n24162,pwm_start_stop[30]}),
    .q({open_n24169,\PWME/RemaTxNum[20]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/reg3_b23  (
    .a({_al_u2841_o,_al_u2841_o}),
    .b({\PWME/n24 ,\PWME/n24 }),
    .c({pnumcntE[23],pnumcntE[23]}),
    .clk(clk100m),
    .d({\PWME/pnumr [23],\PWME/pnumr [23]}),
    .mi({open_n24181,pwm_start_stop[30]}),
    .q({open_n24188,\PWME/RemaTxNum[23]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/reg3_b3  (
    .a({_al_u2839_o,_al_u2839_o}),
    .b({\PWME/n24 ,\PWME/n24 }),
    .c({pnumcntE[3],pnumcntE[3]}),
    .clk(clk100m),
    .d({\PWME/pnumr [3],\PWME/pnumr [3]}),
    .mi({open_n24200,pwm_start_stop[30]}),
    .q({open_n24207,\PWME/RemaTxNum[3]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/reg3_b6  (
    .a({_al_u2833_o,_al_u2833_o}),
    .b({\PWME/n24 ,\PWME/n24 }),
    .c({pnumcntE[6],pnumcntE[6]}),
    .clk(clk100m),
    .d({\PWME/pnumr [6],\PWME/pnumr [6]}),
    .mi({open_n24219,pwm_start_stop[30]}),
    .q({open_n24226,\PWME/RemaTxNum[6]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWME/reg3_b7  (
    .a({_al_u2831_o,_al_u2831_o}),
    .b({\PWME/n24 ,\PWME/n24 }),
    .c({pnumcntE[7],pnumcntE[7]}),
    .clk(clk100m),
    .d({\PWME/pnumr [7],\PWME/pnumr [7]}),
    .mi({open_n24238,pwm_start_stop[30]}),
    .q({open_n24245,\PWME/RemaTxNum[7]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_LSLICE #(
    //.MACRO("PWME/sub0/ucin_al_u3461"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWME/sub0/u11_al_u3464  (
    .a({\PWME/FreCnt [13],\PWME/FreCnt [11]}),
    .b({\PWME/FreCnt [14],\PWME/FreCnt [12]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWME/sub0/c11 ),
    .f({\PWME/n12 [13],\PWME/n12 [11]}),
    .fco(\PWME/sub0/c15 ),
    .fx({\PWME/n12 [14],\PWME/n12 [12]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWME/sub0/ucin_al_u3461"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWME/sub0/u15_al_u3465  (
    .a({\PWME/FreCnt [17],\PWME/FreCnt [15]}),
    .b({\PWME/FreCnt [18],\PWME/FreCnt [16]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWME/sub0/c15 ),
    .f({\PWME/n12 [17],\PWME/n12 [15]}),
    .fco(\PWME/sub0/c19 ),
    .fx({\PWME/n12 [18],\PWME/n12 [16]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWME/sub0/ucin_al_u3461"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWME/sub0/u19_al_u3466  (
    .a({\PWME/FreCnt [21],\PWME/FreCnt [19]}),
    .b({\PWME/FreCnt [22],\PWME/FreCnt [20]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWME/sub0/c19 ),
    .f({\PWME/n12 [21],\PWME/n12 [19]}),
    .fco(\PWME/sub0/c23 ),
    .fx({\PWME/n12 [22],\PWME/n12 [20]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWME/sub0/ucin_al_u3461"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWME/sub0/u23_al_u3467  (
    .a({\PWME/FreCnt [25],\PWME/FreCnt [23]}),
    .b({\PWME/FreCnt [26],\PWME/FreCnt [24]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWME/sub0/c23 ),
    .f({\PWME/n12 [25],\PWME/n12 [23]}),
    .fx({\PWME/n12 [26],\PWME/n12 [24]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWME/sub0/ucin_al_u3461"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWME/sub0/u3_al_u3462  (
    .a({\PWME/FreCnt [5],\PWME/FreCnt [3]}),
    .b({\PWME/FreCnt [6],\PWME/FreCnt [4]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWME/sub0/c3 ),
    .f({\PWME/n12 [5],\PWME/n12 [3]}),
    .fco(\PWME/sub0/c7 ),
    .fx({\PWME/n12 [6],\PWME/n12 [4]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWME/sub0/ucin_al_u3461"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWME/sub0/u7_al_u3463  (
    .a({\PWME/FreCnt [9],\PWME/FreCnt [7]}),
    .b({\PWME/FreCnt [10],\PWME/FreCnt [8]}),
    .c(2'b11),
    .d(2'b00),
    .e(2'b00),
    .fci(\PWME/sub0/c7 ),
    .f({\PWME/n12 [9],\PWME/n12 [7]}),
    .fco(\PWME/sub0/c11 ),
    .fx({\PWME/n12 [10],\PWME/n12 [8]}));
  EF2_PHY_LSLICE #(
    //.MACRO("PWME/sub0/ucin_al_u3461"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h0005),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \PWME/sub0/ucin_al_u3461  (
    .a({\PWME/FreCnt [1],1'b0}),
    .b({\PWME/FreCnt [2],\PWME/FreCnt [0]}),
    .c(2'b11),
    .d(2'b01),
    .e(2'b01),
    .f({\PWME/n12 [1],open_n24372}),
    .fco(\PWME/sub0/c3 ),
    .fx({\PWME/n12 [2],\PWME/n12 [0]}));
  EF2_PHY_MSLICE #(
    //.MACRO("PWME/sub1/u0|PWME/sub1/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("SUB_CARRY"),
    .INIT_LUT0(16'b0000000000000101),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWME/sub1/u0|PWME/sub1/ucin  (
    .a({pnumcntE[0],1'b0}),
    .b({1'b1,open_n24375}),
    .f({\PWME/n26 [0],open_n24395}),
    .fco(\PWME/sub1/c1 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWME/sub1/u0|PWME/sub1/ucin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWME/sub1/u10|PWME/sub1/u9  (
    .a(pnumcntE[10:9]),
    .b(2'b00),
    .fci(\PWME/sub1/c9 ),
    .f(\PWME/n26 [10:9]),
    .fco(\PWME/sub1/c11 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWME/sub1/u0|PWME/sub1/ucin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWME/sub1/u12|PWME/sub1/u11  (
    .a(pnumcntE[12:11]),
    .b(2'b00),
    .fci(\PWME/sub1/c11 ),
    .f(\PWME/n26 [12:11]),
    .fco(\PWME/sub1/c13 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWME/sub1/u0|PWME/sub1/ucin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWME/sub1/u14|PWME/sub1/u13  (
    .a(pnumcntE[14:13]),
    .b(2'b00),
    .fci(\PWME/sub1/c13 ),
    .f(\PWME/n26 [14:13]),
    .fco(\PWME/sub1/c15 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWME/sub1/u0|PWME/sub1/ucin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWME/sub1/u16|PWME/sub1/u15  (
    .a(pnumcntE[16:15]),
    .b(2'b00),
    .fci(\PWME/sub1/c15 ),
    .f(\PWME/n26 [16:15]),
    .fco(\PWME/sub1/c17 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWME/sub1/u0|PWME/sub1/ucin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWME/sub1/u18|PWME/sub1/u17  (
    .a(pnumcntE[18:17]),
    .b(2'b00),
    .fci(\PWME/sub1/c17 ),
    .f(\PWME/n26 [18:17]),
    .fco(\PWME/sub1/c19 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWME/sub1/u0|PWME/sub1/ucin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWME/sub1/u20|PWME/sub1/u19  (
    .a(pnumcntE[20:19]),
    .b(2'b00),
    .fci(\PWME/sub1/c19 ),
    .f(\PWME/n26 [20:19]),
    .fco(\PWME/sub1/c21 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWME/sub1/u0|PWME/sub1/ucin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWME/sub1/u22|PWME/sub1/u21  (
    .a(pnumcntE[22:21]),
    .b(2'b00),
    .fci(\PWME/sub1/c21 ),
    .f(\PWME/n26 [22:21]),
    .fco(\PWME/sub1/c23 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWME/sub1/u0|PWME/sub1/ucin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWME/sub1/u23_al_u3482  (
    .a({open_n24554,pnumcntE[23]}),
    .b({open_n24555,1'b0}),
    .fci(\PWME/sub1/c23 ),
    .f({open_n24574,\PWME/n26 [23]}));
  EF2_PHY_MSLICE #(
    //.MACRO("PWME/sub1/u0|PWME/sub1/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWME/sub1/u2|PWME/sub1/u1  (
    .a(pnumcntE[2:1]),
    .b(2'b00),
    .fci(\PWME/sub1/c1 ),
    .f(\PWME/n26 [2:1]),
    .fco(\PWME/sub1/c3 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWME/sub1/u0|PWME/sub1/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWME/sub1/u4|PWME/sub1/u3  (
    .a(pnumcntE[4:3]),
    .b(2'b00),
    .fci(\PWME/sub1/c3 ),
    .f(\PWME/n26 [4:3]),
    .fco(\PWME/sub1/c5 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWME/sub1/u0|PWME/sub1/ucin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWME/sub1/u6|PWME/sub1/u5  (
    .a(pnumcntE[6:5]),
    .b(2'b00),
    .fci(\PWME/sub1/c5 ),
    .f(\PWME/n26 [6:5]),
    .fco(\PWME/sub1/c7 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWME/sub1/u0|PWME/sub1/ucin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWME/sub1/u8|PWME/sub1/u7  (
    .a(pnumcntE[8:7]),
    .b(2'b00),
    .fci(\PWME/sub1/c7 ),
    .f(\PWME/n26 [8:7]),
    .fco(\PWME/sub1/c9 ));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[0]  (
    .i(\PWMF/RemaTxNum[0]_keep ),
    .o(pnumcntF[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[10]  (
    .i(\PWMF/RemaTxNum[10]_keep ),
    .o(pnumcntF[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[11]  (
    .i(\PWMF/RemaTxNum[11]_keep ),
    .o(pnumcntF[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[12]  (
    .i(\PWMF/RemaTxNum[12]_keep ),
    .o(pnumcntF[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[13]  (
    .i(\PWMF/RemaTxNum[13]_keep ),
    .o(pnumcntF[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[14]  (
    .i(\PWMF/RemaTxNum[14]_keep ),
    .o(pnumcntF[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[15]  (
    .i(\PWMF/RemaTxNum[15]_keep ),
    .o(pnumcntF[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[16]  (
    .i(\PWMF/RemaTxNum[16]_keep ),
    .o(pnumcntF[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[17]  (
    .i(\PWMF/RemaTxNum[17]_keep ),
    .o(pnumcntF[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[18]  (
    .i(\PWMF/RemaTxNum[18]_keep ),
    .o(pnumcntF[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[19]  (
    .i(\PWMF/RemaTxNum[19]_keep ),
    .o(pnumcntF[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[1]  (
    .i(\PWMF/RemaTxNum[1]_keep ),
    .o(pnumcntF[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[20]  (
    .i(\PWMF/RemaTxNum[20]_keep ),
    .o(pnumcntF[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[21]  (
    .i(\PWMF/RemaTxNum[21]_keep ),
    .o(pnumcntF[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[22]  (
    .i(\PWMF/RemaTxNum[22]_keep ),
    .o(pnumcntF[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[23]  (
    .i(\PWMF/RemaTxNum[23]_keep ),
    .o(pnumcntF[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[2]  (
    .i(\PWMF/RemaTxNum[2]_keep ),
    .o(pnumcntF[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[3]  (
    .i(\PWMF/RemaTxNum[3]_keep ),
    .o(pnumcntF[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[4]  (
    .i(\PWMF/RemaTxNum[4]_keep ),
    .o(pnumcntF[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[5]  (
    .i(\PWMF/RemaTxNum[5]_keep ),
    .o(pnumcntF[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[6]  (
    .i(\PWMF/RemaTxNum[6]_keep ),
    .o(pnumcntF[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[7]  (
    .i(\PWMF/RemaTxNum[7]_keep ),
    .o(pnumcntF[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[8]  (
    .i(\PWMF/RemaTxNum[8]_keep ),
    .o(pnumcntF[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[9]  (
    .i(\PWMF/RemaTxNum[9]_keep ),
    .o(pnumcntF[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_dir  (
    .i(\PWMF/dir_keep ),
    .o(dir_pad[15]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[0]  (
    .i(\PWMF/pnumr[0]_keep ),
    .o(\PWMF/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[10]  (
    .i(\PWMF/pnumr[10]_keep ),
    .o(\PWMF/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[11]  (
    .i(\PWMF/pnumr[11]_keep ),
    .o(\PWMF/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[12]  (
    .i(\PWMF/pnumr[12]_keep ),
    .o(\PWMF/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[13]  (
    .i(\PWMF/pnumr[13]_keep ),
    .o(\PWMF/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[14]  (
    .i(\PWMF/pnumr[14]_keep ),
    .o(\PWMF/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[15]  (
    .i(\PWMF/pnumr[15]_keep ),
    .o(\PWMF/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[16]  (
    .i(\PWMF/pnumr[16]_keep ),
    .o(\PWMF/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[17]  (
    .i(\PWMF/pnumr[17]_keep ),
    .o(\PWMF/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[18]  (
    .i(\PWMF/pnumr[18]_keep ),
    .o(\PWMF/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[19]  (
    .i(\PWMF/pnumr[19]_keep ),
    .o(\PWMF/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[1]  (
    .i(\PWMF/pnumr[1]_keep ),
    .o(\PWMF/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[20]  (
    .i(\PWMF/pnumr[20]_keep ),
    .o(\PWMF/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[21]  (
    .i(\PWMF/pnumr[21]_keep ),
    .o(\PWMF/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[22]  (
    .i(\PWMF/pnumr[22]_keep ),
    .o(\PWMF/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[23]  (
    .i(\PWMF/pnumr[23]_keep ),
    .o(\PWMF/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[24]  (
    .i(\PWMF/pnumr[24]_keep ),
    .o(\PWMF/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[25]  (
    .i(\PWMF/pnumr[25]_keep ),
    .o(\PWMF/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[26]  (
    .i(\PWMF/pnumr[26]_keep ),
    .o(\PWMF/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[27]  (
    .i(\PWMF/pnumr[27]_keep ),
    .o(\PWMF/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[28]  (
    .i(\PWMF/pnumr[28]_keep ),
    .o(\PWMF/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[29]  (
    .i(\PWMF/pnumr[29]_keep ),
    .o(\PWMF/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[2]  (
    .i(\PWMF/pnumr[2]_keep ),
    .o(\PWMF/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[30]  (
    .i(\PWMF/pnumr[30]_keep ),
    .o(\PWMF/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[31]  (
    .i(\PWMF/pnumr[31]_keep ),
    .o(\PWMF/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[3]  (
    .i(\PWMF/pnumr[3]_keep ),
    .o(\PWMF/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[4]  (
    .i(\PWMF/pnumr[4]_keep ),
    .o(\PWMF/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[5]  (
    .i(\PWMF/pnumr[5]_keep ),
    .o(\PWMF/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[6]  (
    .i(\PWMF/pnumr[6]_keep ),
    .o(\PWMF/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[7]  (
    .i(\PWMF/pnumr[7]_keep ),
    .o(\PWMF/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[8]  (
    .i(\PWMF/pnumr[8]_keep ),
    .o(\PWMF/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[9]  (
    .i(\PWMF/pnumr[9]_keep ),
    .o(\PWMF/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pwm  (
    .i(\PWMF/pwm_keep ),
    .o(pwm_pad[15]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_stopreq  (
    .i(\PWMF/stopreq_keep ),
    .o(\PWMF/stopreq ));  // src/OnePWM.v(14)
  EF2_PHY_MSLICE #(
    //.LUT0("(D*~(C)*~((~0*~(B*A)))+D*C*~((~0*~(B*A)))+~(D)*C*(~0*~(B*A))+D*C*(~0*~(B*A)))"),
    //.LUT1("(D*~(C)*~((~1*~(B*A)))+D*C*~((~1*~(B*A)))+~(D)*C*(~1*~(B*A))+D*C*(~1*~(B*A)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111100001110000),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/dir_reg  (
    .a({\PWMF/n24 ,\PWMF/n24 }),
    .b({\PWMF/n25_neg_lutinv ,\PWMF/n25_neg_lutinv }),
    .c({dir_pad[15],dir_pad[15]}),
    .clk(clk100m),
    .d({\PWMF/pnumr [31],\PWMF/pnumr [31]}),
    .mi({open_n24679,pwm_start_stop[31]}),
    .q({open_n24686,\PWMF/dir_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("~(~0*~(D*C*B*A))"),
    //.LUT1("~(~1*~(D*C*B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b1111111111111111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMF/pwm_reg  (
    .a({_al_u1625_o,_al_u1625_o}),
    .b({_al_u1632_o,_al_u1632_o}),
    .c({_al_u1634_o,_al_u1634_o}),
    .clk(clk100m),
    .d({_al_u1636_o,_al_u1636_o}),
    .mi({open_n24698,pwm_pad[15]}),
    .sr(\PWMF/u14_sel_is_1_o ),
    .q({open_n24704,\PWMF/pwm_keep }));  // src/OnePWM.v(45)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMF/reg0_b0|PWMF/reg0_b15  (
    .b({\PWMF/n12 [0],\PWMF/n12 [15]}),
    .c({freqF[0],freqF[15]}),
    .clk(clk100m),
    .d({\PWMF/n0_lutinv ,\PWMF/n0_lutinv }),
    .sr(\PWMF/n11 ),
    .q({\PWMF/FreCnt [0],\PWMF/FreCnt [15]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMF/reg0_b10|PWMF/reg0_b1  (
    .b({\PWMF/n12 [10],\PWMF/n12 [1]}),
    .c({freqF[10],freqF[1]}),
    .clk(clk100m),
    .d({\PWMF/n0_lutinv ,\PWMF/n0_lutinv }),
    .sr(\PWMF/n11 ),
    .q({\PWMF/FreCnt [10],\PWMF/FreCnt [1]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMF/reg0_b11|PWMF/reg0_b9  (
    .b({\PWMF/n12 [11],\PWMF/n12 [9]}),
    .c({freqF[11],freqF[9]}),
    .clk(clk100m),
    .d({\PWMF/n0_lutinv ,\PWMF/n0_lutinv }),
    .sr(\PWMF/n11 ),
    .q({\PWMF/FreCnt [11],\PWMF/FreCnt [9]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMF/reg0_b12|PWMF/reg0_b8  (
    .b({\PWMF/n12 [12],\PWMF/n12 [8]}),
    .c({freqF[12],freqF[8]}),
    .clk(clk100m),
    .d({\PWMF/n0_lutinv ,\PWMF/n0_lutinv }),
    .sr(\PWMF/n11 ),
    .q({\PWMF/FreCnt [12],\PWMF/FreCnt [8]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMF/reg0_b13|PWMF/reg0_b7  (
    .b({\PWMF/n12 [13],\PWMF/n12 [7]}),
    .c({freqF[13],freqF[7]}),
    .clk(clk100m),
    .d({\PWMF/n0_lutinv ,\PWMF/n0_lutinv }),
    .sr(\PWMF/n11 ),
    .q({\PWMF/FreCnt [13],\PWMF/FreCnt [7]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMF/reg0_b14|PWMF/reg0_b5  (
    .b({\PWMF/n12 [14],\PWMF/n12 [5]}),
    .c({freqF[14],freqF[5]}),
    .clk(clk100m),
    .d({\PWMF/n0_lutinv ,\PWMF/n0_lutinv }),
    .sr(\PWMF/n11 ),
    .q({\PWMF/FreCnt [14],\PWMF/FreCnt [5]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMF/reg0_b16|PWMF/reg0_b3  (
    .b({\PWMF/n12 [16],\PWMF/n12 [3]}),
    .c({freqF[16],freqF[3]}),
    .clk(clk100m),
    .d({\PWMF/n0_lutinv ,\PWMF/n0_lutinv }),
    .sr(\PWMF/n11 ),
    .q({\PWMF/FreCnt [16],\PWMF/FreCnt [3]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMF/reg0_b17|PWMF/reg0_b25  (
    .b({\PWMF/n12 [17],\PWMF/n12 [25]}),
    .c({freqF[17],freqF[25]}),
    .clk(clk100m),
    .d({\PWMF/n0_lutinv ,\PWMF/n0_lutinv }),
    .sr(\PWMF/n11 ),
    .q({\PWMF/FreCnt [17],\PWMF/FreCnt [25]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMF/reg0_b18|PWMF/reg0_b23  (
    .b({\PWMF/n12 [18],\PWMF/n12 [23]}),
    .c({freqF[18],freqF[23]}),
    .clk(clk100m),
    .d({\PWMF/n0_lutinv ,\PWMF/n0_lutinv }),
    .sr(\PWMF/n11 ),
    .q({\PWMF/FreCnt [18],\PWMF/FreCnt [23]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMF/reg0_b19|PWMF/reg0_b21  (
    .b({\PWMF/n12 [19],\PWMF/n12 [21]}),
    .c({freqF[19],freqF[21]}),
    .clk(clk100m),
    .d({\PWMF/n0_lutinv ,\PWMF/n0_lutinv }),
    .sr(\PWMF/n11 ),
    .q({\PWMF/FreCnt [19],\PWMF/FreCnt [21]}));  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMF/reg0_b2  (
    .b({open_n24923,\PWMF/n12 [2]}),
    .c({open_n24924,freqF[2]}),
    .clk(clk100m),
    .d({open_n24926,\PWMF/n0_lutinv }),
    .sr(\PWMF/n11 ),
    .q({open_n24944,\PWMF/FreCnt [2]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMF/reg0_b20|PWMF/reg0_b6  (
    .b({\PWMF/n12 [20],\PWMF/n12 [6]}),
    .c({freqF[20],freqF[6]}),
    .clk(clk100m),
    .d({\PWMF/n0_lutinv ,\PWMF/n0_lutinv }),
    .sr(\PWMF/n11 ),
    .q({\PWMF/FreCnt [20],\PWMF/FreCnt [6]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1111000011001100),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1111000011001100),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMF/reg0_b22|PWMF/reg0_b4  (
    .b({\PWMF/n12 [22],\PWMF/n12 [4]}),
    .c({freqF[22],freqF[4]}),
    .clk(clk100m),
    .d({\PWMF/n0_lutinv ,\PWMF/n0_lutinv }),
    .sr(\PWMF/n11 ),
    .q({\PWMF/FreCnt [22],\PWMF/FreCnt [4]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111000011001100),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \PWMF/reg0_b24|PWMF/reg0_b26  (
    .b({\PWMF/n12 [24],\PWMF/n12 [26]}),
    .c({freqF[24],freqF[26]}),
    .clk(clk100m),
    .d({\PWMF/n0_lutinv ,\PWMF/n0_lutinv }),
    .sr(\PWMF/n11 ),
    .q({\PWMF/FreCnt [24],\PWMF/FreCnt [26]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*~C)*~(~0*B))"),
    //.LUTF1("(~(~C*B)*~(D*~A))"),
    //.LUTG0("(A*~(D*~C)*~(~1*B))"),
    //.LUTG1("(~(~C*B)*~(D*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010000000100010),
    .INIT_LUTF1(16'b1010001011110011),
    .INIT_LUTG0(16'b1010000010101010),
    .INIT_LUTG1(16'b1010001011110011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg1_b10|PWMF/reg1_b26  (
    .a({\PWMF/FreCnt [8],_al_u2971_o}),
    .b({\PWMF/FreCnt [9],\PWMF/FreCnt [25]}),
    .c({\PWMF/FreCntr [10],\PWMF/FreCnt [9]}),
    .ce(\PWMF/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMF/FreCntr [9],\PWMF/FreCntr [10]}),
    .e({open_n25013,\PWMF/FreCntr [26]}),
    .mi({freqF[10],freqF[26]}),
    .f({_al_u2974_o,_al_u2972_o}),
    .q({\PWMF/FreCntr [10],\PWMF/FreCntr [26]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*~C)*~(~D*B))"),
    //.LUTF1("(A*~(0*~C)*~(D*~B))"),
    //.LUTG0("(A*~(1*~C)*~(~D*B))"),
    //.LUTG1("(A*~(1*~C)*~(D*~B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101000100010),
    .INIT_LUTF1(16'b1000100010101010),
    .INIT_LUTG0(16'b1010000000100000),
    .INIT_LUTG1(16'b1000000010100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg1_b14|PWMF/reg1_b18  (
    .a({_al_u2974_o,_al_u2976_o}),
    .b({\PWMF/FreCnt [13],\PWMF/FreCnt [17]}),
    .c({\PWMF/FreCnt [17],\PWMF/FreCnt [19]}),
    .ce(\PWMF/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMF/FreCntr [14],\PWMF/FreCntr [18]}),
    .e({\PWMF/FreCntr [18],\PWMF/FreCntr [20]}),
    .mi({freqF[14],freqF[18]}),
    .f({_al_u2975_o,_al_u2977_o}),
    .q({\PWMF/FreCntr [14],\PWMF/FreCntr [18]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*B*A*~(0@D))"),
    //.LUTF1("(~(D*~B)*~(~C*A))"),
    //.LUTG0("(C*B*A*~(1@D))"),
    //.LUTG1("(~(D*~B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b1100010011110101),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b1100010011110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg1_b16|PWMF/reg1_b13  (
    .a({\PWMF/FreCnt [15],_al_u2966_o}),
    .b({\PWMF/FreCnt [25],_al_u2968_o}),
    .c({\PWMF/FreCntr [16],_al_u2969_o}),
    .ce(\PWMF/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMF/FreCntr [26],\PWMF/FreCnt [12]}),
    .e({open_n25046,\PWMF/FreCntr [13]}),
    .mi({freqF[16],freqF[13]}),
    .f({_al_u2969_o,_al_u2970_o}),
    .q({\PWMF/FreCntr [16],\PWMF/FreCntr [13]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(D*~B)*~(C*~A))"),
    //.LUTF1("(B*A*~(D@C))"),
    //.LUTG0("(~(D*~B)*~(C*~A))"),
    //.LUTG1("(B*A*~(D@C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000110010101111),
    .INIT_LUTF1(16'b1000000000001000),
    .INIT_LUTG0(16'b1000110010101111),
    .INIT_LUTG1(16'b1000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg1_b17|PWMF/reg1_b11  (
    .a({_al_u2964_o,\PWMF/FreCnt [10]}),
    .b({_al_u2965_o,\PWMF/FreCnt [21]}),
    .c({\PWMF/FreCnt [16],\PWMF/FreCntr [11]}),
    .ce(\PWMF/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMF/FreCntr [17],\PWMF/FreCntr [22]}),
    .mi({freqF[17],freqF[11]}),
    .f({_al_u2966_o,_al_u2965_o}),
    .q({\PWMF/FreCntr [17],\PWMF/FreCntr [11]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(D@B)*~(C@A))"),
    //.LUTF1("(B*A*~(D@C))"),
    //.LUTG0("(~(D@B)*~(C@A))"),
    //.LUTG1("(B*A*~(D@C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000010000100001),
    .INIT_LUTF1(16'b1000000000001000),
    .INIT_LUTG0(16'b1000010000100001),
    .INIT_LUTG1(16'b1000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg1_b21|PWMF/reg1_b19  (
    .a({_al_u1626_o,\PWMF/FreCnt [18]}),
    .b({_al_u1627_o,\PWMF/FreCnt [20]}),
    .c({\PWMF/FreCnt [21],\PWMF/FreCntr [19]}),
    .ce(\PWMF/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMF/FreCntr [21],\PWMF/FreCntr [21]}),
    .mi({freqF[21],freqF[19]}),
    .f({_al_u1628_o,_al_u2964_o}),
    .q({\PWMF/FreCntr [21],\PWMF/FreCntr [19]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~A*~(0@C)*~(~D*B))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(~A*~(1@C)*~(~D*B))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010100000001),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b0101000000010000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg1_b22|PWMF/reg1_b20  (
    .a({\PWMF/FreCnt [22],_al_u2961_o}),
    .b({\PWMF/FreCnt [23],\PWMF/FreCnt [19]}),
    .c({\PWMF/FreCntr [22],\PWMF/FreCnt [22]}),
    .ce(\PWMF/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMF/FreCntr [23],\PWMF/FreCntr [20]}),
    .e({open_n25099,\PWMF/FreCntr [23]}),
    .mi({freqF[22],freqF[20]}),
    .f({_al_u1620_o,_al_u2962_o}),
    .q({\PWMF/FreCntr [22],\PWMF/FreCntr [20]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg1_b23|PWMF/reg1_b0  (
    .b({_al_u1293_o,open_n25118}),
    .c({_al_u1295_o,\PWMF/n11 }),
    .ce(\PWMF/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({_al_u1291_o,\PWMF/n0_lutinv }),
    .mi({freqF[23],freqF[0]}),
    .f({\PWMF/n0_lutinv ,\PWMF/mux3_b0_sel_is_3_o }),
    .q({\PWMF/FreCntr [23],\PWMF/FreCntr [0]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*~C)*~(~D*B))"),
    //.LUTF1("(~(D*~B)*~(C*~A))"),
    //.LUTG0("(A*~(1*~C)*~(~D*B))"),
    //.LUTG1("(~(D*~B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101000100010),
    .INIT_LUTF1(16'b1000110010101111),
    .INIT_LUTG0(16'b1010000000100000),
    .INIT_LUTG1(16'b1000110010101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg1_b24|PWMF/reg1_b4  (
    .a({\PWMF/FreCnt [23],_al_u2967_o}),
    .b({\PWMF/FreCnt [3],\PWMF/FreCnt [3]}),
    .c({\PWMF/FreCntr [24],\PWMF/FreCnt [7]}),
    .ce(\PWMF/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMF/FreCntr [4],\PWMF/FreCntr [4]}),
    .e({open_n25137,\PWMF/FreCntr [8]}),
    .mi({freqF[24],freqF[4]}),
    .f({_al_u2971_o,_al_u2968_o}),
    .q({\PWMF/FreCntr [24],\PWMF/FreCntr [4]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*B*A*~(0@D))"),
    //.LUTF1("(~(C@B)*~(D@A))"),
    //.LUTG0("(C*B*A*~(1@D))"),
    //.LUTG1("(~(C@B)*~(D@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b1000001001000001),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b1000001001000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg1_b25|PWMF/reg1_b3  (
    .a({\PWMF/FreCnt [2],_al_u1621_o}),
    .b({\PWMF/FreCnt [24],_al_u1623_o}),
    .c({\PWMF/FreCntr [25],_al_u1624_o}),
    .ce(\PWMF/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMF/FreCntr [3],\PWMF/FreCnt [3]}),
    .e({open_n25154,\PWMF/FreCntr [3]}),
    .mi({freqF[25],freqF[3]}),
    .f({_al_u2955_o,_al_u1625_o}),
    .q({\PWMF/FreCntr [25],\PWMF/FreCntr [3]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*~C)*~(~0*B))"),
    //.LUTF1("(~(~D*B)*~(C*~A))"),
    //.LUTG0("(A*~(D*~C)*~(~1*B))"),
    //.LUTG1("(~(~D*B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010000000100010),
    .INIT_LUTF1(16'b1010111100100011),
    .INIT_LUTG0(16'b1010000010101010),
    .INIT_LUTG1(16'b1010111100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg1_b2|PWMF/reg1_b15  (
    .a({\PWMF/FreCnt [1],_al_u2959_o}),
    .b({\PWMF/FreCnt [21],\PWMF/FreCnt [1]}),
    .c({\PWMF/FreCntr [2],\PWMF/FreCnt [14]}),
    .ce(\PWMF/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMF/FreCntr [22],\PWMF/FreCntr [15]}),
    .e({open_n25171,\PWMF/FreCntr [2]}),
    .mi({freqF[2],freqF[15]}),
    .f({_al_u2976_o,_al_u2960_o}),
    .q({\PWMF/FreCntr [2],\PWMF/FreCntr [15]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(D@B)*~(C@A))"),
    //.LUT1("(D*~(C@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000010000100001),
    .INIT_LUT1(16'b1100001100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg1_b5|PWMF/reg1_b12  (
    .a({open_n25188,\PWMF/FreCnt [11]}),
    .b({\PWMF/FreCnt [4],\PWMF/FreCnt [6]}),
    .c({\PWMF/FreCntr [5],\PWMF/FreCntr [12]}),
    .ce(\PWMF/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({_al_u2957_o,\PWMF/FreCntr [7]}),
    .mi({freqF[5],freqF[12]}),
    .f({_al_u2958_o,_al_u2957_o}),
    .q({\PWMF/FreCntr [5],\PWMF/FreCntr [12]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(~0*C)*~(D@B))"),
    //.LUTF1("(~(D*~B)*~(~C*A))"),
    //.LUTG0("(A*~(~1*C)*~(D@B))"),
    //.LUTG1("(~(D*~B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b1100010011110101),
    .INIT_LUTG0(16'b1000100000100010),
    .INIT_LUTG1(16'b1100010011110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg1_b6|PWMF/reg1_b1  (
    .a({\PWMF/FreCnt [14],_al_u2972_o}),
    .b({\PWMF/FreCnt [5],\PWMF/FreCnt [0]}),
    .c({\PWMF/FreCntr [15],\PWMF/FreCnt [5]}),
    .ce(\PWMF/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMF/FreCntr [6],\PWMF/FreCntr [1]}),
    .e({open_n25203,\PWMF/FreCntr [6]}),
    .mi({freqF[6],freqF[1]}),
    .f({_al_u2954_o,_al_u2973_o}),
    .q({\PWMF/FreCntr [6],\PWMF/FreCntr [1]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~D*B)*~(C*~A))"),
    //.LUT1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010111100100011),
    .INIT_LUT1(16'b1000010000100001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg1_b7|PWMF/reg1_b8  (
    .a({\PWMF/FreCnt [6],\PWMF/FreCnt [15]}),
    .b({\PWMF/FreCnt [7],\PWMF/FreCnt [7]}),
    .c({\PWMF/FreCntr [6],\PWMF/FreCntr [16]}),
    .ce(\PWMF/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMF/FreCntr [7],\PWMF/FreCntr [8]}),
    .mi({freqF[7],freqF[8]}),
    .f({_al_u1622_o,_al_u2959_o}),
    .q({\PWMF/FreCntr [7],\PWMF/FreCntr [8]}));  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg1_b9  (
    .c({open_n25238,\PWMF/FreCntr [9]}),
    .ce(\PWMF/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({open_n25239,\PWMF/FreCnt [8]}),
    .mi({open_n25250,freqF[9]}),
    .f({open_n25252,_al_u2961_o}),
    .q({open_n25256,\PWMF/FreCntr [9]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg2_b0|PWMF/reg3_b0  (
    .a({\PWMF/pnumr [0],_al_u2952_o}),
    .b({pnumF[0],\PWMF/n24 }),
    .c({pnumF[32],pnumcntF[0]}),
    .clk(clk100m),
    .d({pwm_start_stop[31],\PWMF/pnumr [0]}),
    .e({open_n25258,pwm_start_stop[31]}),
    .q({\PWMF/pnumr[0]_keep ,\PWMF/RemaTxNum[0]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011100010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011100010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg2_b10|PWMF/reg2_b8  (
    .a({\PWMF/pnumr [10],\PWMF/pnumr [8]}),
    .b({pnumF[10],pnumF[32]}),
    .c({pnumF[32],pnumF[8]}),
    .clk(clk100m),
    .d({pwm_start_stop[31],pwm_start_stop[31]}),
    .q({\PWMF/pnumr[10]_keep ,\PWMF/pnumr[8]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg2_b11|PWMF/reg3_b11  (
    .a({\PWMF/pnumr [11],_al_u2946_o}),
    .b({pnumF[11],\PWMF/n24 }),
    .c({pnumF[32],pnumcntF[11]}),
    .clk(clk100m),
    .d({pwm_start_stop[31],\PWMF/pnumr [11]}),
    .e({open_n25303,pwm_start_stop[31]}),
    .q({\PWMF/pnumr[11]_keep ,\PWMF/RemaTxNum[11]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg2_b12|PWMF/reg3_b12  (
    .a({\PWMF/pnumr [12],_al_u2944_o}),
    .b({pnumF[12],\PWMF/n24 }),
    .c({pnumF[32],pnumcntF[12]}),
    .clk(clk100m),
    .d({pwm_start_stop[31],\PWMF/pnumr [12]}),
    .e({open_n25325,pwm_start_stop[31]}),
    .q({\PWMF/pnumr[12]_keep ,\PWMF/RemaTxNum[12]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011100010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011100010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg2_b13|PWMF/reg2_b7  (
    .a({\PWMF/pnumr [13],\PWMF/pnumr [7]}),
    .b({pnumF[13],pnumF[32]}),
    .c({pnumF[32],pnumF[7]}),
    .clk(clk100m),
    .d({pwm_start_stop[31],pwm_start_stop[31]}),
    .q({\PWMF/pnumr[13]_keep ,\PWMF/pnumr[7]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011100010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg2_b14|PWMF/reg2_b4  (
    .a({\PWMF/pnumr [14],\PWMF/pnumr [4]}),
    .b({pnumF[14],pnumF[32]}),
    .c({pnumF[32],pnumF[4]}),
    .clk(clk100m),
    .d({pwm_start_stop[31],pwm_start_stop[31]}),
    .q({\PWMF/pnumr[14]_keep ,\PWMF/pnumr[4]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg2_b15|PWMF/reg3_b15  (
    .a({\PWMF/pnumr [15],_al_u2938_o}),
    .b({pnumF[15],\PWMF/n24 }),
    .c({pnumF[32],pnumcntF[15]}),
    .clk(clk100m),
    .d({pwm_start_stop[31],\PWMF/pnumr [15]}),
    .e({open_n25389,pwm_start_stop[31]}),
    .q({\PWMF/pnumr[15]_keep ,\PWMF/RemaTxNum[15]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg2_b16|PWMF/reg3_b16  (
    .a({\PWMF/pnumr [16],_al_u2936_o}),
    .b({pnumF[16],\PWMF/n24 }),
    .c({pnumF[32],pnumcntF[16]}),
    .clk(clk100m),
    .d({pwm_start_stop[31],\PWMF/pnumr [16]}),
    .e({open_n25411,pwm_start_stop[31]}),
    .q({\PWMF/pnumr[16]_keep ,\PWMF/RemaTxNum[16]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg2_b17|PWMF/reg2_b3  (
    .a({\PWMF/pnumr [17],\PWMF/pnumr [3]}),
    .b({pnumF[17],pnumF[3]}),
    .c({pnumF[32],pnumF[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[31],pwm_start_stop[31]}),
    .q({\PWMF/pnumr[17]_keep ,\PWMF/pnumr[3]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg2_b18|PWMF/reg2_b21  (
    .a({\PWMF/pnumr [18],\PWMF/pnumr [21]}),
    .b({pnumF[18],pnumF[21]}),
    .c({pnumF[32],pnumF[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[31],pwm_start_stop[31]}),
    .q({\PWMF/pnumr[18]_keep ,\PWMF/pnumr[21]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg2_b19|PWMF/reg3_b19  (
    .a({\PWMF/pnumr [19],_al_u2930_o}),
    .b({pnumF[19],\PWMF/n24 }),
    .c({pnumF[32],pnumcntF[19]}),
    .clk(clk100m),
    .d({pwm_start_stop[31],\PWMF/pnumr [19]}),
    .e({open_n25475,pwm_start_stop[31]}),
    .q({\PWMF/pnumr[19]_keep ,\PWMF/RemaTxNum[19]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg2_b1|PWMF/reg2_b20  (
    .a({\PWMF/pnumr [1],\PWMF/pnumr [20]}),
    .b({pnumF[1],pnumF[20]}),
    .c({pnumF[32],pnumF[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[31],pwm_start_stop[31]}),
    .q({\PWMF/pnumr[1]_keep ,\PWMF/pnumr[20]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg2_b22|PWMF/reg3_b22  (
    .a({\PWMF/pnumr [22],_al_u2922_o}),
    .b({pnumF[22],\PWMF/n24 }),
    .c({pnumF[32],pnumcntF[22]}),
    .clk(clk100m),
    .d({pwm_start_stop[31],\PWMF/pnumr [22]}),
    .e({open_n25520,pwm_start_stop[31]}),
    .q({\PWMF/pnumr[22]_keep ,\PWMF/RemaTxNum[22]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg2_b23|PWMF/reg3_b23  (
    .a({\PWMF/pnumr [23],_al_u2920_o}),
    .b({pnumF[23],\PWMF/n24 }),
    .c({pnumF[32],pnumcntF[23]}),
    .clk(clk100m),
    .d({pwm_start_stop[31],\PWMF/pnumr [23]}),
    .e({open_n25542,pwm_start_stop[31]}),
    .q({\PWMF/pnumr[23]_keep ,\PWMF/RemaTxNum[23]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg2_b24|PWMF/reg2_b31  (
    .a({\PWMF/pnumr [24],\PWMF/pnumr [31]}),
    .b({pnumF[24],pnumF[31]}),
    .c({pnumF[32],pnumF[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[31],pwm_start_stop[31]}),
    .q({\PWMF/pnumr[24]_keep ,\PWMF/pnumr[31]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg2_b25|PWMF/reg2_b30  (
    .a({\PWMF/pnumr [25],\PWMF/pnumr [30]}),
    .b({pnumF[25],pnumF[30]}),
    .c({pnumF[32],pnumF[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[31],pwm_start_stop[31]}),
    .q({\PWMF/pnumr[25]_keep ,\PWMF/pnumr[30]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1100000011001010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg2_b26|PWMF/reg2_b29  (
    .a({\PWMF/pnumr [26],\PWMF/pnumr [29]}),
    .b({pnumF[26],pnumF[29]}),
    .c({pnumF[32],pnumF[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[31],pwm_start_stop[31]}),
    .q({\PWMF/pnumr[26]_keep ,\PWMF/pnumr[29]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg2_b27|PWMF/reg2_b28  (
    .a({\PWMF/pnumr [27],\PWMF/pnumr [28]}),
    .b({pnumF[27],pnumF[28]}),
    .c({pnumF[32],pnumF[32]}),
    .clk(clk100m),
    .d({pwm_start_stop[31],pwm_start_stop[31]}),
    .q({\PWMF/pnumr[27]_keep ,\PWMF/pnumr[28]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011001010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011001010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg2_b2|PWMF/reg3_b2  (
    .a({\PWMF/pnumr [2],_al_u2928_o}),
    .b({pnumF[2],\PWMF/n24 }),
    .c({pnumF[32],pnumcntF[2]}),
    .clk(clk100m),
    .d({pwm_start_stop[31],\PWMF/pnumr [2]}),
    .e({open_n25644,pwm_start_stop[31]}),
    .q({\PWMF/pnumr[2]_keep ,\PWMF/RemaTxNum[2]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg2_b5|PWMF/reg3_b5  (
    .a({\PWMF/pnumr [5],_al_u2914_o}),
    .b({pnumF[32],\PWMF/n24 }),
    .c({pnumF[5],pnumcntF[5]}),
    .clk(clk100m),
    .d({pwm_start_stop[31],\PWMF/pnumr [5]}),
    .e({open_n25666,pwm_start_stop[31]}),
    .q({\PWMF/pnumr[5]_keep ,\PWMF/RemaTxNum[5]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg2_b6|PWMF/reg3_b6  (
    .a({\PWMF/pnumr [6],_al_u2912_o}),
    .b({pnumF[32],\PWMF/n24 }),
    .c({pnumF[6],pnumcntF[6]}),
    .clk(clk100m),
    .d({pwm_start_stop[31],\PWMF/pnumr [6]}),
    .e({open_n25688,pwm_start_stop[31]}),
    .q({\PWMF/pnumr[6]_keep ,\PWMF/RemaTxNum[6]_keep }));  // src/OnePWM.v(58)
  // src/OnePWM.v(58)
  // src/OnePWM.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1100000011100010),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1100000011100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg2_b9|PWMF/reg3_b9  (
    .a({\PWMF/pnumr [9],_al_u2906_o}),
    .b({pnumF[32],\PWMF/n24 }),
    .c({pnumF[9],pnumcntF[9]}),
    .clk(clk100m),
    .d({pwm_start_stop[31],\PWMF/pnumr [9]}),
    .e({open_n25710,pwm_start_stop[31]}),
    .q({\PWMF/pnumr[9]_keep ,\PWMF/RemaTxNum[9]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg3_b1  (
    .a({_al_u2950_o,_al_u2950_o}),
    .b({\PWMF/n24 ,\PWMF/n24 }),
    .c({pnumcntF[1],pnumcntF[1]}),
    .clk(clk100m),
    .d({\PWMF/pnumr [1],\PWMF/pnumr [1]}),
    .mi({open_n25742,pwm_start_stop[31]}),
    .q({open_n25749,\PWMF/RemaTxNum[1]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg3_b10  (
    .a({_al_u2948_o,_al_u2948_o}),
    .b({\PWMF/n24 ,\PWMF/n24 }),
    .c({pnumcntF[10],pnumcntF[10]}),
    .clk(clk100m),
    .d({\PWMF/pnumr [10],\PWMF/pnumr [10]}),
    .mi({open_n25761,pwm_start_stop[31]}),
    .q({open_n25768,\PWMF/RemaTxNum[10]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg3_b13  (
    .a({_al_u2942_o,_al_u2942_o}),
    .b({\PWMF/n24 ,\PWMF/n24 }),
    .c({pnumcntF[13],pnumcntF[13]}),
    .clk(clk100m),
    .d({\PWMF/pnumr [13],\PWMF/pnumr [13]}),
    .mi({open_n25780,pwm_start_stop[31]}),
    .q({open_n25787,\PWMF/RemaTxNum[13]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg3_b14  (
    .a({_al_u2940_o,_al_u2940_o}),
    .b({\PWMF/n24 ,\PWMF/n24 }),
    .c({pnumcntF[14],pnumcntF[14]}),
    .clk(clk100m),
    .d({\PWMF/pnumr [14],\PWMF/pnumr [14]}),
    .mi({open_n25799,pwm_start_stop[31]}),
    .q({open_n25806,\PWMF/RemaTxNum[14]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg3_b17  (
    .a({_al_u2934_o,_al_u2934_o}),
    .b({\PWMF/n24 ,\PWMF/n24 }),
    .c({pnumcntF[17],pnumcntF[17]}),
    .clk(clk100m),
    .d({\PWMF/pnumr [17],\PWMF/pnumr [17]}),
    .mi({open_n25818,pwm_start_stop[31]}),
    .q({open_n25825,\PWMF/RemaTxNum[17]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg3_b18  (
    .a({_al_u2932_o,_al_u2932_o}),
    .b({\PWMF/n24 ,\PWMF/n24 }),
    .c({pnumcntF[18],pnumcntF[18]}),
    .clk(clk100m),
    .d({\PWMF/pnumr [18],\PWMF/pnumr [18]}),
    .mi({open_n25837,pwm_start_stop[31]}),
    .q({open_n25844,\PWMF/RemaTxNum[18]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg3_b20  (
    .a({_al_u2926_o,_al_u2926_o}),
    .b({\PWMF/n24 ,\PWMF/n24 }),
    .c({pnumcntF[20],pnumcntF[20]}),
    .clk(clk100m),
    .d({\PWMF/pnumr [20],\PWMF/pnumr [20]}),
    .mi({open_n25856,pwm_start_stop[31]}),
    .q({open_n25863,\PWMF/RemaTxNum[20]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg3_b21  (
    .a({_al_u2924_o,_al_u2924_o}),
    .b({\PWMF/n24 ,\PWMF/n24 }),
    .c({pnumcntF[21],pnumcntF[21]}),
    .clk(clk100m),
    .d({\PWMF/pnumr [21],\PWMF/pnumr [21]}),
    .mi({open_n25875,pwm_start_stop[31]}),
    .q({open_n25882,\PWMF/RemaTxNum[21]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg3_b3  (
    .a({_al_u2918_o,_al_u2918_o}),
    .b({\PWMF/n24 ,\PWMF/n24 }),
    .c({pnumcntF[3],pnumcntF[3]}),
    .clk(clk100m),
    .d({\PWMF/pnumr [3],\PWMF/pnumr [3]}),
    .mi({open_n25894,pwm_start_stop[31]}),
    .q({open_n25901,\PWMF/RemaTxNum[3]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg3_b4  (
    .a({_al_u2916_o,_al_u2916_o}),
    .b({\PWMF/n24 ,\PWMF/n24 }),
    .c({pnumcntF[4],pnumcntF[4]}),
    .clk(clk100m),
    .d({\PWMF/pnumr [4],\PWMF/pnumr [4]}),
    .mi({open_n25913,pwm_start_stop[31]}),
    .q({open_n25920,\PWMF/RemaTxNum[4]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg3_b7  (
    .a({_al_u2910_o,_al_u2910_o}),
    .b({\PWMF/n24 ,\PWMF/n24 }),
    .c({pnumcntF[7],pnumcntF[7]}),
    .clk(clk100m),
    .d({\PWMF/pnumr [7],\PWMF/pnumr [7]}),
    .mi({open_n25932,pwm_start_stop[31]}),
    .q({open_n25939,\PWMF/RemaTxNum[7]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUT1("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1011101010111010),
    .INIT_LUT1(16'b1111111100000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \PWMF/reg3_b8  (
    .a({_al_u2908_o,_al_u2908_o}),
    .b({\PWMF/n24 ,\PWMF/n24 }),
    .c({pnumcntF[8],pnumcntF[8]}),
    .clk(clk100m),
    .d({\PWMF/pnumr [8],\PWMF/pnumr [8]}),
    .mi({open_n25951,pwm_start_stop[31]}),
    .q({open_n25958,\PWMF/RemaTxNum[8]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.MACRO("PWMF/sub0/u0|PWMF/sub0/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("SUB_CARRY"),
    .INIT_LUT0(16'b0000000000000101),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMF/sub0/u0|PWMF/sub0/ucin  (
    .a({\PWMF/FreCnt [0],1'b0}),
    .b({1'b1,open_n25959}),
    .f({\PWMF/n12 [0],open_n25979}),
    .fco(\PWMF/sub0/c1 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMF/sub0/u0|PWMF/sub0/ucin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMF/sub0/u10|PWMF/sub0/u9  (
    .a(\PWMF/FreCnt [10:9]),
    .b(2'b00),
    .fci(\PWMF/sub0/c9 ),
    .f(\PWMF/n12 [10:9]),
    .fco(\PWMF/sub0/c11 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMF/sub0/u0|PWMF/sub0/ucin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMF/sub0/u12|PWMF/sub0/u11  (
    .a(\PWMF/FreCnt [12:11]),
    .b(2'b00),
    .fci(\PWMF/sub0/c11 ),
    .f(\PWMF/n12 [12:11]),
    .fco(\PWMF/sub0/c13 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMF/sub0/u0|PWMF/sub0/ucin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMF/sub0/u14|PWMF/sub0/u13  (
    .a(\PWMF/FreCnt [14:13]),
    .b(2'b00),
    .fci(\PWMF/sub0/c13 ),
    .f(\PWMF/n12 [14:13]),
    .fco(\PWMF/sub0/c15 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMF/sub0/u0|PWMF/sub0/ucin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMF/sub0/u16|PWMF/sub0/u15  (
    .a(\PWMF/FreCnt [16:15]),
    .b(2'b00),
    .fci(\PWMF/sub0/c15 ),
    .f(\PWMF/n12 [16:15]),
    .fco(\PWMF/sub0/c17 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMF/sub0/u0|PWMF/sub0/ucin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMF/sub0/u18|PWMF/sub0/u17  (
    .a(\PWMF/FreCnt [18:17]),
    .b(2'b00),
    .fci(\PWMF/sub0/c17 ),
    .f(\PWMF/n12 [18:17]),
    .fco(\PWMF/sub0/c19 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMF/sub0/u0|PWMF/sub0/ucin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMF/sub0/u20|PWMF/sub0/u19  (
    .a(\PWMF/FreCnt [20:19]),
    .b(2'b00),
    .fci(\PWMF/sub0/c19 ),
    .f(\PWMF/n12 [20:19]),
    .fco(\PWMF/sub0/c21 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMF/sub0/u0|PWMF/sub0/ucin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMF/sub0/u22|PWMF/sub0/u21  (
    .a(\PWMF/FreCnt [22:21]),
    .b(2'b00),
    .fci(\PWMF/sub0/c21 ),
    .f(\PWMF/n12 [22:21]),
    .fco(\PWMF/sub0/c23 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMF/sub0/u0|PWMF/sub0/ucin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMF/sub0/u24|PWMF/sub0/u23  (
    .a(\PWMF/FreCnt [24:23]),
    .b(2'b00),
    .fci(\PWMF/sub0/c23 ),
    .f(\PWMF/n12 [24:23]),
    .fco(\PWMF/sub0/c25 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMF/sub0/u0|PWMF/sub0/ucin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMF/sub0/u26|PWMF/sub0/u25  (
    .a(\PWMF/FreCnt [26:25]),
    .b(2'b00),
    .fci(\PWMF/sub0/c25 ),
    .f(\PWMF/n12 [26:25]));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMF/sub0/u0|PWMF/sub0/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMF/sub0/u2|PWMF/sub0/u1  (
    .a(\PWMF/FreCnt [2:1]),
    .b(2'b00),
    .fci(\PWMF/sub0/c1 ),
    .f(\PWMF/n12 [2:1]),
    .fco(\PWMF/sub0/c3 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMF/sub0/u0|PWMF/sub0/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMF/sub0/u4|PWMF/sub0/u3  (
    .a(\PWMF/FreCnt [4:3]),
    .b(2'b00),
    .fci(\PWMF/sub0/c3 ),
    .f(\PWMF/n12 [4:3]),
    .fco(\PWMF/sub0/c5 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMF/sub0/u0|PWMF/sub0/ucin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMF/sub0/u6|PWMF/sub0/u5  (
    .a(\PWMF/FreCnt [6:5]),
    .b(2'b00),
    .fci(\PWMF/sub0/c5 ),
    .f(\PWMF/n12 [6:5]),
    .fco(\PWMF/sub0/c7 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMF/sub0/u0|PWMF/sub0/ucin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMF/sub0/u8|PWMF/sub0/u7  (
    .a(\PWMF/FreCnt [8:7]),
    .b(2'b00),
    .fci(\PWMF/sub0/c7 ),
    .f(\PWMF/n12 [8:7]),
    .fco(\PWMF/sub0/c9 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMF/sub1/u0|PWMF/sub1/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("SUB_CARRY"),
    .INIT_LUT0(16'b0000000000000101),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMF/sub1/u0|PWMF/sub1/ucin  (
    .a({pnumcntF[0],1'b0}),
    .b({1'b1,open_n26271}),
    .f({\PWMF/n26 [0],open_n26291}),
    .fco(\PWMF/sub1/c1 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMF/sub1/u0|PWMF/sub1/ucin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMF/sub1/u10|PWMF/sub1/u9  (
    .a(pnumcntF[10:9]),
    .b(2'b00),
    .fci(\PWMF/sub1/c9 ),
    .f(\PWMF/n26 [10:9]),
    .fco(\PWMF/sub1/c11 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMF/sub1/u0|PWMF/sub1/ucin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMF/sub1/u12|PWMF/sub1/u11  (
    .a(pnumcntF[12:11]),
    .b(2'b00),
    .fci(\PWMF/sub1/c11 ),
    .f(\PWMF/n26 [12:11]),
    .fco(\PWMF/sub1/c13 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMF/sub1/u0|PWMF/sub1/ucin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMF/sub1/u14|PWMF/sub1/u13  (
    .a(pnumcntF[14:13]),
    .b(2'b00),
    .fci(\PWMF/sub1/c13 ),
    .f(\PWMF/n26 [14:13]),
    .fco(\PWMF/sub1/c15 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMF/sub1/u0|PWMF/sub1/ucin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMF/sub1/u16|PWMF/sub1/u15  (
    .a(pnumcntF[16:15]),
    .b(2'b00),
    .fci(\PWMF/sub1/c15 ),
    .f(\PWMF/n26 [16:15]),
    .fco(\PWMF/sub1/c17 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMF/sub1/u0|PWMF/sub1/ucin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMF/sub1/u18|PWMF/sub1/u17  (
    .a(pnumcntF[18:17]),
    .b(2'b00),
    .fci(\PWMF/sub1/c17 ),
    .f(\PWMF/n26 [18:17]),
    .fco(\PWMF/sub1/c19 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMF/sub1/u0|PWMF/sub1/ucin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMF/sub1/u20|PWMF/sub1/u19  (
    .a(pnumcntF[20:19]),
    .b(2'b00),
    .fci(\PWMF/sub1/c19 ),
    .f(\PWMF/n26 [20:19]),
    .fco(\PWMF/sub1/c21 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMF/sub1/u0|PWMF/sub1/ucin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMF/sub1/u22|PWMF/sub1/u21  (
    .a(pnumcntF[22:21]),
    .b(2'b00),
    .fci(\PWMF/sub1/c21 ),
    .f(\PWMF/n26 [22:21]),
    .fco(\PWMF/sub1/c23 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMF/sub1/u0|PWMF/sub1/ucin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMF/sub1/u23_al_u3483  (
    .a({open_n26450,pnumcntF[23]}),
    .b({open_n26451,1'b0}),
    .fci(\PWMF/sub1/c23 ),
    .f({open_n26470,\PWMF/n26 [23]}));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMF/sub1/u0|PWMF/sub1/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMF/sub1/u2|PWMF/sub1/u1  (
    .a(pnumcntF[2:1]),
    .b(2'b00),
    .fci(\PWMF/sub1/c1 ),
    .f(\PWMF/n26 [2:1]),
    .fco(\PWMF/sub1/c3 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMF/sub1/u0|PWMF/sub1/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMF/sub1/u4|PWMF/sub1/u3  (
    .a(pnumcntF[4:3]),
    .b(2'b00),
    .fci(\PWMF/sub1/c3 ),
    .f(\PWMF/n26 [4:3]),
    .fco(\PWMF/sub1/c5 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMF/sub1/u0|PWMF/sub1/ucin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMF/sub1/u6|PWMF/sub1/u5  (
    .a(pnumcntF[6:5]),
    .b(2'b00),
    .fci(\PWMF/sub1/c5 ),
    .f(\PWMF/n26 [6:5]),
    .fco(\PWMF/sub1/c7 ));
  EF2_PHY_MSLICE #(
    //.MACRO("PWMF/sub1/u0|PWMF/sub1/ucin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \PWMF/sub1/u8|PWMF/sub1/u7  (
    .a(pnumcntF[8:7]),
    .b(2'b00),
    .fci(\PWMF/sub1/c7 ),
    .f(\PWMF/n26 [8:7]),
    .fco(\PWMF/sub1/c9 ));
  EF2_PHY_MCU #(
    .GPIO_L0("ENABLE"),
    .GPIO_L1("ENABLE"),
    .GPIO_L10("DISABLE"),
    .GPIO_L11("DISABLE"),
    .GPIO_L12("DISABLE"),
    .GPIO_L13("DISABLE"),
    .GPIO_L14("DISABLE"),
    .GPIO_L15("DISABLE"),
    .GPIO_L2("DISABLE"),
    .GPIO_L3("DISABLE"),
    .GPIO_L4("DISABLE"),
    .GPIO_L5("DISABLE"),
    .GPIO_L6("DISABLE"),
    .GPIO_L7("DISABLE"),
    .GPIO_L8("ENABLE"),
    .GPIO_L9("ENABLE"))
    \U_AHB/M3WithAHB/mcu_inst  (
    .gpio_h_in(16'b0000000000000000),
    .h2h_hrdata(\U_AHB/h2h_hrdata ),
    .h2h_hreadyout(1'b1),
    .h2h_hresp(2'b00),
    .h2h_mclk(clk100m),
    .h2h_rstn(rstn),
    .ppm_clk(clk25m),
    .h2h_haddr({open_n26607,open_n26608,open_n26609,open_n26610,open_n26611,open_n26612,open_n26613,open_n26614,open_n26615,open_n26616,open_n26617,open_n26618,open_n26619,open_n26620,open_n26621,open_n26622,open_n26623,\U_AHB/h2h_haddrw [14:2],open_n26624,open_n26625}),
    .h2h_hwdata(\U_AHB/h2h_hwdata ),
    .h2h_hwrite(\U_AHB/h2h_hwritew ));  // al_ip/M3WithAHB.v(46)
  // src/AHB.v(25)
  // src/AHB.v(24)
  EF2_PHY_MSLICE #(
    //.LUT0("(D*C*B*A)"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/h2h_hwrite_reg|U_AHB/reg0_b1  (
    .a({\U_AHB/h2h_hwrite ,\U_AHB/h2h_hwrite }),
    .b({\U_AHB/h2h_haddr [13],\U_AHB/h2h_haddr [3]}),
    .c(\U_AHB/h2h_haddr [14:13]),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [4],\U_AHB/h2h_haddr [14]}),
    .mi({\U_AHB/h2h_hwritew ,\U_AHB/h2h_haddrw [3]}),
    .f({\U_AHB/n77 ,\U_AHB/n75 }),
    .q({\U_AHB/h2h_hwrite ,\U_AHB/h2h_haddr [3]}));  // src/AHB.v(25)
  // src/AHB.v(25)
  // src/AHB.v(25)
  EF2_PHY_MSLICE #(
    //.LUT0("(D*C*~B*A)"),
    //.LUT1("(D*~C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010000000000000),
    .INIT_LUT1(16'b0000100000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg0_b10|U_AHB/reg0_b2  (
    .a({\U_AHB/h2h_hwrite ,\U_AHB/h2h_hwrite }),
    .b({\U_AHB/h2h_haddr [12],\U_AHB/h2h_haddr [13]}),
    .c({\U_AHB/h2h_haddr [13],\U_AHB/h2h_haddr [14]}),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [14],\U_AHB/h2h_haddr [4]}),
    .mi({\U_AHB/h2h_haddrw [12],\U_AHB/h2h_haddrw [4]}),
    .f({\U_AHB/n71 ,\U_AHB/n55 }),
    .q({\U_AHB/h2h_haddr [12],\U_AHB/h2h_haddr [4]}));  // src/AHB.v(25)
  // src/AHB.v(25)
  // src/AHB.v(25)
  EF2_PHY_MSLICE #(
    //.LUT0("(D*C*B*A)"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg0_b12|U_AHB/reg0_b0  (
    .a({\U_AHB/h2h_hwrite ,\U_AHB/h2h_hwrite }),
    .b({\U_AHB/h2h_haddr [13],\U_AHB/h2h_haddr [2]}),
    .c(\U_AHB/h2h_haddr [14:13]),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [5],\U_AHB/h2h_haddr [14]}),
    .mi({\U_AHB/h2h_haddrw [14],\U_AHB/h2h_haddrw [2]}),
    .f({\U_AHB/n45 ,\U_AHB/n73 }),
    .q({\U_AHB/h2h_haddr [14],\U_AHB/h2h_haddr [2]}));  // src/AHB.v(25)
  // src/AHB.v(25)
  // src/AHB.v(25)
  EF2_PHY_MSLICE #(
    //.LUT0("(D*C*~B*A)"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010000000000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg0_b4|U_AHB/reg0_b3  (
    .a({\U_AHB/h2h_hwrite ,\U_AHB/h2h_hwrite }),
    .b({\U_AHB/h2h_haddr [13],\U_AHB/h2h_haddr [13]}),
    .c({\U_AHB/h2h_haddr [14],\U_AHB/h2h_haddr [14]}),
    .clk(clk100m),
    .d(\U_AHB/h2h_haddr [6:5]),
    .mi(\U_AHB/h2h_haddrw [6:5]),
    .f({\U_AHB/n47 ,\U_AHB/n57 }),
    .q(\U_AHB/h2h_haddr [6:5]));  // src/AHB.v(25)
  // src/AHB.v(25)
  // src/AHB.v(25)
  EF2_PHY_MSLICE #(
    //.LUT0("(D*C*B*A)"),
    //.LUT1("(D*C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b0010000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg0_b5|U_AHB/reg0_b11  (
    .a({\U_AHB/h2h_hwrite ,\U_AHB/h2h_hwrite }),
    .b({\U_AHB/h2h_haddr [13],\U_AHB/h2h_haddr [13]}),
    .c({\U_AHB/h2h_haddr [14],\U_AHB/h2h_haddr [14]}),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [7],\U_AHB/h2h_haddr [7]}),
    .mi({\U_AHB/h2h_haddrw [7],\U_AHB/h2h_haddrw [13]}),
    .f({\U_AHB/n61 ,\U_AHB/n79 }),
    .q({\U_AHB/h2h_haddr [7],\U_AHB/h2h_haddr [13]}));  // src/AHB.v(25)
  // src/AHB.v(25)
  // src/AHB.v(25)
  EF2_PHY_MSLICE #(
    //.LUT0("(D*C*~B*A)"),
    //.LUT1("(D*C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010000000000000),
    .INIT_LUT1(16'b0010000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg0_b6|U_AHB/reg0_b8  (
    .a({\U_AHB/h2h_hwrite ,\U_AHB/h2h_hwrite }),
    .b({\U_AHB/h2h_haddr [13],\U_AHB/h2h_haddr [13]}),
    .c({\U_AHB/h2h_haddr [14],\U_AHB/h2h_haddr [14]}),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [8],\U_AHB/h2h_haddr [10]}),
    .mi({\U_AHB/h2h_haddrw [8],\U_AHB/h2h_haddrw [10]}),
    .f({\U_AHB/n63 ,\U_AHB/n67 }),
    .q({\U_AHB/h2h_haddr [8],\U_AHB/h2h_haddr [10]}));  // src/AHB.v(25)
  // src/AHB.v(25)
  // src/AHB.v(25)
  EF2_PHY_MSLICE #(
    //.LUT0("(D*C*~B*A)"),
    //.LUT1("(D*C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0010000000000000),
    .INIT_LUT1(16'b0010000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg0_b7|U_AHB/reg0_b9  (
    .a({\U_AHB/h2h_hwrite ,\U_AHB/h2h_hwrite }),
    .b({\U_AHB/h2h_haddr [13],\U_AHB/h2h_haddr [13]}),
    .c({\U_AHB/h2h_haddr [14],\U_AHB/h2h_haddr [14]}),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [9],\U_AHB/h2h_haddr [11]}),
    .mi({\U_AHB/h2h_haddrw [9],\U_AHB/h2h_haddrw [11]}),
    .f({\U_AHB/n65 ,\U_AHB/n69 }),
    .q({\U_AHB/h2h_haddr [9],\U_AHB/h2h_haddr [11]}));  // src/AHB.v(25)
  // src/AHB.v(55)
  // src/AHB.v(55)
  EF2_PHY_LSLICE #(
    //.LUTF0("(0*~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C))"),
    //.LUTF1("(D*~C*~B*A)"),
    //.LUTG0("(1*~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C))"),
    //.LUTG1("(D*~C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000001000000000),
    .INIT_LUTG0(16'b0101001101011111),
    .INIT_LUTG1(16'b0000001000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg10_b0|U_AHB/reg10_b13  (
    .a({\U_AHB/h2h_hwrite ,pnumcntB[18]}),
    .b({\U_AHB/h2h_haddr [13],pnumcntC[18]}),
    .c({\U_AHB/h2h_haddr [14],\U_AHB/h2h_haddr [2]}),
    .ce(\U_AHB/n22 ),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [9],\U_AHB/h2h_haddr [3]}),
    .e({open_n26770,\U_AHB/h2h_haddr [13]}),
    .mi({\U_AHB/h2h_hwdata [0],\U_AHB/h2h_hwdata [13]}),
    .f({\U_AHB/n22 ,_al_u3238_o}),
    .q({freq9[0],freq9[13]}));  // src/AHB.v(55)
  // src/AHB.v(55)
  // src/AHB.v(55)
  EF2_PHY_MSLICE #(
    //.LUT0("(~C*~B*~D)"),
    //.LUT1("(~C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000011),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg10_b10|U_AHB/reg10_b1  (
    .b({open_n26789,\U_AHB/h2h_haddr [13]}),
    .c({\U_AHB/h2h_haddr [14],\U_AHB/h2h_haddr [14]}),
    .ce(\U_AHB/n22 ),
    .clk(clk100m),
    .d({\U_AHB/h2h_hwrite ,\U_AHB/h2h_hwrite }),
    .mi({\U_AHB/h2h_hwdata [10],\U_AHB/h2h_hwdata [1]}),
    .f({_al_u3061_o,\U_AHB/n82 }),
    .q({freq9[10],freq9[1]}));  // src/AHB.v(55)
  // src/AHB.v(55)
  // src/AHB.v(55)
  EF2_PHY_MSLICE #(
    //.LUT0("(D*~C*B*A)"),
    //.LUT1("(~D*~C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100000000000),
    .INIT_LUT1(16'b0000000000000010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg10_b14|U_AHB/reg10_b11  (
    .a({\U_AHB/n95_lutinv ,\U_AHB/h2h_hwrite }),
    .b({\U_AHB/h2h_haddr [7],\U_AHB/h2h_haddr [13]}),
    .c({\U_AHB/h2h_haddr [8],\U_AHB/h2h_haddr [14]}),
    .ce(\U_AHB/n22 ),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [9],\U_AHB/h2h_haddr [7]}),
    .mi({\U_AHB/h2h_hwdata [14],\U_AHB/h2h_hwdata [11]}),
    .f({\U_AHB/n104_lutinv ,\U_AHB/n36 }),
    .q({freq9[14],freq9[11]}));  // src/AHB.v(55)
  // src/AHB.v(55)
  // src/AHB.v(55)
  EF2_PHY_MSLICE #(
    //.LUT0("(D*~C*B*A)"),
    //.LUT1("(D*~C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100000000000),
    .INIT_LUT1(16'b0000001000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg10_b15|U_AHB/reg10_b12  (
    .a({\U_AHB/n95_lutinv ,\U_AHB/h2h_hwrite }),
    .b({\U_AHB/h2h_haddr [7],\U_AHB/h2h_haddr [13]}),
    .c({\U_AHB/h2h_haddr [8],\U_AHB/h2h_haddr [14]}),
    .ce(\U_AHB/n22 ),
    .clk(clk100m),
    .d(\U_AHB/h2h_haddr [9:8]),
    .mi({\U_AHB/h2h_hwdata [15],\U_AHB/h2h_hwdata [12]}),
    .f({\U_AHB/n102 ,\U_AHB/n38 }),
    .q({freq9[15],freq9[12]}));  // src/AHB.v(55)
  // src/AHB.v(55)
  // src/AHB.v(55)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg10_b17|U_AHB/reg10_b16  (
    .a({_al_u3171_o,_al_u3175_o}),
    .b({\U_AHB/n113_lutinv ,\U_AHB/n104_lutinv }),
    .c({\U_AHB/n111 ,\U_AHB/n102 }),
    .ce(\U_AHB/n22 ),
    .clk(clk100m),
    .d({pnumcntA[23],\U_AHB/h2h_hrdata [23]}),
    .e({\U_AHB/h2h_hrdata [23],limit_l_pad[7]}),
    .mi(\U_AHB/h2h_hwdata [17:16]),
    .f({_al_u3172_o,_al_u3176_o}),
    .q(freq9[17:16]));  // src/AHB.v(55)
  // src/AHB.v(55)
  // src/AHB.v(55)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg10_b19|U_AHB/reg10_b18  (
    .a({_al_u3182_o,_al_u3186_o}),
    .b({\U_AHB/n113_lutinv ,\U_AHB/n104_lutinv }),
    .c({\U_AHB/n111 ,\U_AHB/n102 }),
    .ce(\U_AHB/n22 ),
    .clk(clk100m),
    .d({pnumcntA[22],\U_AHB/h2h_hrdata [22]}),
    .e({\U_AHB/h2h_hrdata [22],limit_l_pad[6]}),
    .mi(\U_AHB/h2h_hwdata [19:18]),
    .f({_al_u3183_o,_al_u3187_o}),
    .q(freq9[19:18]));  // src/AHB.v(55)
  // src/AHB.v(55)
  // src/AHB.v(55)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg10_b20|U_AHB/reg10_b2  (
    .a({_al_u3193_o,_al_u3197_o}),
    .b({\U_AHB/n113_lutinv ,\U_AHB/n104_lutinv }),
    .c({\U_AHB/n111 ,\U_AHB/n102 }),
    .ce(\U_AHB/n22 ),
    .clk(clk100m),
    .d({pnumcntA[21],\U_AHB/h2h_hrdata [21]}),
    .e({\U_AHB/h2h_hrdata [21],limit_l_pad[5]}),
    .mi({\U_AHB/h2h_hwdata [20],\U_AHB/h2h_hwdata [2]}),
    .f({_al_u3194_o,_al_u3198_o}),
    .q({freq9[20],freq9[2]}));  // src/AHB.v(55)
  // src/AHB.v(55)
  // src/AHB.v(55)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg10_b22|U_AHB/reg10_b21  (
    .a({_al_u3204_o,_al_u3208_o}),
    .b({\U_AHB/n113_lutinv ,\U_AHB/n104_lutinv }),
    .c({\U_AHB/n111 ,\U_AHB/n102 }),
    .ce(\U_AHB/n22 ),
    .clk(clk100m),
    .d({pnumcntA[20],\U_AHB/h2h_hrdata [20]}),
    .e({\U_AHB/h2h_hrdata [20],limit_l_pad[4]}),
    .mi(\U_AHB/h2h_hwdata [22:21]),
    .f({_al_u3205_o,_al_u3209_o}),
    .q(freq9[22:21]));  // src/AHB.v(55)
  // src/AHB.v(55)
  // src/AHB.v(55)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg10_b24|U_AHB/reg10_b23  (
    .a({_al_u3226_o,_al_u3230_o}),
    .b({\U_AHB/n113_lutinv ,\U_AHB/n104_lutinv }),
    .c({\U_AHB/n111 ,\U_AHB/n102 }),
    .ce(\U_AHB/n22 ),
    .clk(clk100m),
    .d({pnumcntA[19],\U_AHB/h2h_hrdata [19]}),
    .e({\U_AHB/h2h_hrdata [19],limit_l_pad[3]}),
    .mi(\U_AHB/h2h_hwdata [24:23]),
    .f({_al_u3227_o,_al_u3231_o}),
    .q(freq9[24:23]));  // src/AHB.v(55)
  // src/AHB.v(55)
  // src/AHB.v(55)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg10_b3|U_AHB/reg10_b26  (
    .a({_al_u3248_o,_al_u3252_o}),
    .b({\U_AHB/n113_lutinv ,\U_AHB/n104_lutinv }),
    .c({\U_AHB/n111 ,\U_AHB/n102 }),
    .ce(\U_AHB/n22 ),
    .clk(clk100m),
    .d({pnumcntA[17],\U_AHB/h2h_hrdata [17]}),
    .e({\U_AHB/h2h_hrdata [17],limit_l_pad[1]}),
    .mi({\U_AHB/h2h_hwdata [3],\U_AHB/h2h_hwdata [26]}),
    .f({_al_u3249_o,_al_u3253_o}),
    .q({freq9[3],freq9[26]}));  // src/AHB.v(55)
  // src/AHB.v(55)
  // src/AHB.v(55)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg10_b5|U_AHB/reg10_b4  (
    .a({_al_u3259_o,_al_u3263_o}),
    .b({\U_AHB/n113_lutinv ,\U_AHB/n104_lutinv }),
    .c({\U_AHB/n111 ,\U_AHB/n102 }),
    .ce(\U_AHB/n22 ),
    .clk(clk100m),
    .d({pnumcntA[16],\U_AHB/h2h_hrdata [16]}),
    .e({\U_AHB/h2h_hrdata [16],limit_l_pad[0]}),
    .mi(\U_AHB/h2h_hwdata [5:4]),
    .f({_al_u3260_o,_al_u3264_o}),
    .q(freq9[5:4]));  // src/AHB.v(55)
  // src/AHB.v(55)
  // src/AHB.v(55)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg10_b7|U_AHB/reg10_b6  (
    .a({_al_u3270_o,_al_u3274_o}),
    .b({\U_AHB/n113_lutinv ,\U_AHB/n104_lutinv }),
    .c({\U_AHB/n111 ,\U_AHB/n102 }),
    .ce(\U_AHB/n22 ),
    .clk(clk100m),
    .d({pnumcntA[15],\U_AHB/h2h_hrdata [15]}),
    .e({\U_AHB/h2h_hrdata [15],limit_r_pad[15]}),
    .mi(\U_AHB/h2h_hwdata [7:6]),
    .f({_al_u3271_o,_al_u3275_o}),
    .q(freq9[7:6]));  // src/AHB.v(55)
  // src/AHB.v(55)
  // src/AHB.v(55)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg10_b9|U_AHB/reg10_b8  (
    .a({_al_u3281_o,_al_u3285_o}),
    .b({\U_AHB/n113_lutinv ,\U_AHB/n104_lutinv }),
    .c({\U_AHB/n111 ,\U_AHB/n102 }),
    .ce(\U_AHB/n22 ),
    .clk(clk100m),
    .d({pnumcntA[14],\U_AHB/h2h_hrdata [14]}),
    .e({\U_AHB/h2h_hrdata [14],limit_r_pad[14]}),
    .mi(\U_AHB/h2h_hwdata [9:8]),
    .f({_al_u3282_o,_al_u3286_o}),
    .q(freq9[9:8]));  // src/AHB.v(55)
  // src/AHB.v(56)
  // src/AHB.v(56)
  EF2_PHY_MSLICE #(
    //.LUT0("(D*~C*~B*A)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000000000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg11_b10|U_AHB/reg11_b0  (
    .a({open_n26976,\U_AHB/h2h_hwrite }),
    .b({open_n26977,\U_AHB/h2h_haddr [13]}),
    .c({\U_AHB/h2h_haddr [10],\U_AHB/h2h_haddr [14]}),
    .ce(\U_AHB/n24 ),
    .clk(clk100m),
    .d({\U_AHB/n104_lutinv ,\U_AHB/h2h_haddr [10]}),
    .mi({\U_AHB/h2h_hwdata [10],\U_AHB/h2h_hwdata [0]}),
    .f({\U_AHB/n105 ,\U_AHB/n24 }),
    .q({freqA[10],freqA[0]}));  // src/AHB.v(56)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*~B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg11_b11  (
    .b({open_n26994,\U_AHB/h2h_haddr [10]}),
    .c({open_n26995,\U_AHB/h2h_haddr [11]}),
    .ce(\U_AHB/n24 ),
    .clk(clk100m),
    .d({open_n26996,\U_AHB/n104_lutinv }),
    .mi({open_n27007,\U_AHB/h2h_hwdata [11]}),
    .f({open_n27009,\U_AHB/n108 }),
    .q({open_n27013,freqA[11]}));  // src/AHB.v(56)
  // src/AHB.v(56)
  // src/AHB.v(56)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg11_b14|U_AHB/reg11_b13  (
    .a({_al_u3292_o,_al_u3296_o}),
    .b({\U_AHB/n113_lutinv ,\U_AHB/n104_lutinv }),
    .c({\U_AHB/n111 ,\U_AHB/n102 }),
    .ce(\U_AHB/n24 ),
    .clk(clk100m),
    .d({pnumcntA[13],\U_AHB/h2h_hrdata [13]}),
    .e({\U_AHB/h2h_hrdata [13],limit_r_pad[13]}),
    .mi(\U_AHB/h2h_hwdata [14:13]),
    .f({_al_u3293_o,_al_u3297_o}),
    .q(freqA[14:13]));  // src/AHB.v(56)
  // src/AHB.v(56)
  // src/AHB.v(56)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg11_b16|U_AHB/reg11_b15  (
    .a({_al_u3303_o,_al_u3307_o}),
    .b({\U_AHB/n113_lutinv ,\U_AHB/n104_lutinv }),
    .c({\U_AHB/n111 ,\U_AHB/n102 }),
    .ce(\U_AHB/n24 ),
    .clk(clk100m),
    .d({pnumcntA[12],\U_AHB/h2h_hrdata [12]}),
    .e({\U_AHB/h2h_hrdata [12],limit_r_pad[12]}),
    .mi(\U_AHB/h2h_hwdata [16:15]),
    .f({_al_u3304_o,_al_u3308_o}),
    .q(freqA[16:15]));  // src/AHB.v(56)
  // src/AHB.v(56)
  // src/AHB.v(56)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg11_b18|U_AHB/reg11_b17  (
    .a({_al_u3314_o,_al_u3318_o}),
    .b({\U_AHB/n113_lutinv ,\U_AHB/n104_lutinv }),
    .c({\U_AHB/n111 ,\U_AHB/n102 }),
    .ce(\U_AHB/n24 ),
    .clk(clk100m),
    .d({pnumcntA[11],\U_AHB/h2h_hrdata [11]}),
    .e({\U_AHB/h2h_hrdata [11],limit_r_pad[11]}),
    .mi(\U_AHB/h2h_hwdata [18:17]),
    .f({_al_u3315_o,_al_u3319_o}),
    .q(freqA[18:17]));  // src/AHB.v(56)
  // src/AHB.v(56)
  // src/AHB.v(56)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~D*~C*~B*A)"),
    //.LUTF1("(~D*~C*B*A)"),
    //.LUTG0("(~D*~C*~B*A)"),
    //.LUTG1("(~D*~C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000001000),
    .INIT_LUTG0(16'b0000000000000010),
    .INIT_LUTG1(16'b0000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg11_b1|U_AHB/reg11_b12  (
    .a({\U_AHB/n104_lutinv ,\U_AHB/n104_lutinv }),
    .b({\U_AHB/h2h_haddr [12],\U_AHB/h2h_haddr [12]}),
    .c({\U_AHB/h2h_haddr [10],\U_AHB/h2h_haddr [10]}),
    .ce(\U_AHB/n24 ),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [11],\U_AHB/h2h_haddr [11]}),
    .mi({\U_AHB/h2h_hwdata [1],\U_AHB/h2h_hwdata [12]}),
    .f({\U_AHB/n111 ,\U_AHB/n113_lutinv }),
    .q({freqA[1],freqA[12]}));  // src/AHB.v(56)
  // src/AHB.v(56)
  // src/AHB.v(56)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg11_b21|U_AHB/reg11_b20  (
    .a({_al_u3092_o,_al_u3097_o}),
    .b({\U_AHB/n113_lutinv ,\U_AHB/n104_lutinv }),
    .c({\U_AHB/n111 ,\U_AHB/n102 }),
    .ce(\U_AHB/n24 ),
    .clk(clk100m),
    .d({pnumcntA[9],\U_AHB/h2h_hrdata [9]}),
    .e({\U_AHB/h2h_hrdata [9],limit_r_pad[9]}),
    .mi(\U_AHB/h2h_hwdata [21:20]),
    .f({_al_u3094_o,_al_u3098_o}),
    .q(freqA[21:20]));  // src/AHB.v(56)
  // src/AHB.v(56)
  // src/AHB.v(56)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg11_b23|U_AHB/reg11_b22  (
    .a({_al_u3104_o,_al_u3108_o}),
    .b({\U_AHB/n113_lutinv ,\U_AHB/n104_lutinv }),
    .c({\U_AHB/n111 ,\U_AHB/n102 }),
    .ce(\U_AHB/n24 ),
    .clk(clk100m),
    .d({pnumcntA[8],\U_AHB/h2h_hrdata [8]}),
    .e({\U_AHB/h2h_hrdata [8],limit_r_pad[8]}),
    .mi(\U_AHB/h2h_hwdata [23:22]),
    .f({_al_u3105_o,_al_u3109_o}),
    .q(freqA[23:22]));  // src/AHB.v(56)
  // src/AHB.v(56)
  // src/AHB.v(56)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg11_b25|U_AHB/reg11_b24  (
    .a({_al_u3115_o,_al_u3119_o}),
    .b({\U_AHB/n113_lutinv ,\U_AHB/n104_lutinv }),
    .c({\U_AHB/n111 ,\U_AHB/n102 }),
    .ce(\U_AHB/n24 ),
    .clk(clk100m),
    .d({pnumcntA[7],\U_AHB/h2h_hrdata [7]}),
    .e({\U_AHB/h2h_hrdata [7],limit_r_pad[7]}),
    .mi(\U_AHB/h2h_hwdata [25:24]),
    .f({_al_u3116_o,_al_u3120_o}),
    .q(freqA[25:24]));  // src/AHB.v(56)
  // src/AHB.v(56)
  // src/AHB.v(56)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg11_b2|U_AHB/reg11_b19  (
    .a({_al_u3325_o,_al_u3329_o}),
    .b({\U_AHB/n113_lutinv ,\U_AHB/n104_lutinv }),
    .c({\U_AHB/n111 ,\U_AHB/n102 }),
    .ce(\U_AHB/n24 ),
    .clk(clk100m),
    .d({pnumcntA[10],\U_AHB/h2h_hrdata [10]}),
    .e({\U_AHB/h2h_hrdata [10],limit_r_pad[10]}),
    .mi({\U_AHB/h2h_hwdata [2],\U_AHB/h2h_hwdata [19]}),
    .f({_al_u3326_o,_al_u3330_o}),
    .q({freqA[2],freqA[19]}));  // src/AHB.v(56)
  // src/AHB.v(56)
  // src/AHB.v(56)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg11_b3|U_AHB/reg11_b26  (
    .a({_al_u3126_o,_al_u3130_o}),
    .b({\U_AHB/n113_lutinv ,\U_AHB/n104_lutinv }),
    .c({\U_AHB/n111 ,\U_AHB/n102 }),
    .ce(\U_AHB/n24 ),
    .clk(clk100m),
    .d({pnumcntA[6],\U_AHB/h2h_hrdata [6]}),
    .e({\U_AHB/h2h_hrdata [6],limit_r_pad[6]}),
    .mi({\U_AHB/h2h_hwdata [3],\U_AHB/h2h_hwdata [26]}),
    .f({_al_u3127_o,_al_u3131_o}),
    .q({freqA[3],freqA[26]}));  // src/AHB.v(56)
  // src/AHB.v(56)
  // src/AHB.v(56)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg11_b5|U_AHB/reg11_b4  (
    .a({_al_u3137_o,_al_u3142_o}),
    .b({\U_AHB/n113_lutinv ,\U_AHB/n104_lutinv }),
    .c({\U_AHB/n111 ,\U_AHB/n102 }),
    .ce(\U_AHB/n24 ),
    .clk(clk100m),
    .d({pnumcntA[5],\U_AHB/h2h_hrdata [5]}),
    .e({\U_AHB/h2h_hrdata [5],limit_r_pad[5]}),
    .mi(\U_AHB/h2h_hwdata [5:4]),
    .f({_al_u3138_o,_al_u3143_o}),
    .q(freqA[5:4]));  // src/AHB.v(56)
  // src/AHB.v(56)
  // src/AHB.v(56)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg11_b7|U_AHB/reg11_b6  (
    .a({_al_u3149_o,_al_u3153_o}),
    .b({\U_AHB/n113_lutinv ,\U_AHB/n104_lutinv }),
    .c({\U_AHB/n111 ,\U_AHB/n102 }),
    .ce(\U_AHB/n24 ),
    .clk(clk100m),
    .d({pnumcntA[4],\U_AHB/h2h_hrdata [4]}),
    .e({\U_AHB/h2h_hrdata [4],limit_r_pad[4]}),
    .mi(\U_AHB/h2h_hwdata [7:6]),
    .f({_al_u3150_o,_al_u3154_o}),
    .q(freqA[7:6]));  // src/AHB.v(56)
  // src/AHB.v(56)
  // src/AHB.v(56)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg11_b9|U_AHB/reg11_b8  (
    .a({_al_u3160_o,_al_u3164_o}),
    .b({\U_AHB/n113_lutinv ,\U_AHB/n104_lutinv }),
    .c({\U_AHB/n111 ,\U_AHB/n102 }),
    .ce(\U_AHB/n24 ),
    .clk(clk100m),
    .d({pnumcntA[3],\U_AHB/h2h_hrdata [3]}),
    .e({\U_AHB/h2h_hrdata [3],limit_r_pad[3]}),
    .mi(\U_AHB/h2h_hwdata [9:8]),
    .f({_al_u3161_o,_al_u3165_o}),
    .q(freqA[9:8]));  // src/AHB.v(56)
  // src/AHB.v(57)
  // src/AHB.v(57)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg12_b10|U_AHB/reg12_b1  (
    .a({_al_u3215_o,_al_u3219_o}),
    .b({\U_AHB/n113_lutinv ,\U_AHB/n104_lutinv }),
    .c({\U_AHB/n111 ,\U_AHB/n102 }),
    .ce(\U_AHB/n26 ),
    .clk(clk100m),
    .d({pnumcntA[2],\U_AHB/h2h_hrdata [2]}),
    .e({\U_AHB/h2h_hrdata [2],limit_r_pad[2]}),
    .mi({\U_AHB/h2h_hwdata [10],\U_AHB/h2h_hwdata [1]}),
    .f({_al_u3216_o,_al_u3220_o}),
    .q({freqB[10],freqB[1]}));  // src/AHB.v(57)
  // src/AHB.v(57)
  // src/AHB.v(57)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg12_b12|U_AHB/reg12_b11  (
    .a({_al_u3336_o,_al_u3340_o}),
    .b({\U_AHB/n113_lutinv ,\U_AHB/n104_lutinv }),
    .c({\U_AHB/n111 ,\U_AHB/n102 }),
    .ce(\U_AHB/n26 ),
    .clk(clk100m),
    .d({pnumcntA[1],\U_AHB/h2h_hrdata [1]}),
    .e({\U_AHB/h2h_hrdata [1],limit_r_pad[1]}),
    .mi(\U_AHB/h2h_hwdata [12:11]),
    .f({_al_u3337_o,_al_u3341_o}),
    .q(freqB[12:11]));  // src/AHB.v(57)
  // src/AHB.v(57)
  // src/AHB.v(57)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*C)*~(D*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(1*C)*~(D*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000001010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg12_b14|U_AHB/reg12_b13  (
    .a({_al_u3347_o,_al_u3351_o}),
    .b({\U_AHB/n113_lutinv ,\U_AHB/n104_lutinv }),
    .c({\U_AHB/n111 ,\U_AHB/n102 }),
    .ce(\U_AHB/n26 ),
    .clk(clk100m),
    .d({pnumcntA[0],\U_AHB/h2h_hrdata [0]}),
    .e({\U_AHB/h2h_hrdata [0],limit_r_pad[0]}),
    .mi(\U_AHB/h2h_hwdata [14:13]),
    .f({_al_u3348_o,_al_u3352_o}),
    .q(freqB[14:13]));  // src/AHB.v(57)
  // src/AHB.v(57)
  // src/AHB.v(57)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*B*A*~(0@D))"),
    //.LUTF1("(~(~D*B)*~(~C*A))"),
    //.LUTG0("(C*B*A*~(1@D))"),
    //.LUTG1("(~(~D*B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b1111010100110001),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b1111010100110001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg12_b15|U_AHB/reg12_b21  (
    .a({\PWMB/FreCnt [12],_al_u1558_o}),
    .b({\PWMB/FreCnt [15],_al_u1560_o}),
    .c({\PWMB/FreCntr [12],_al_u1561_o}),
    .ce(\U_AHB/n26 ),
    .clk(clk100m),
    .d({\PWMB/FreCntr [15],\PWMB/FreCnt [21]}),
    .e({open_n27256,\PWMB/FreCntr [21]}),
    .mi({\U_AHB/h2h_hwdata [15],\U_AHB/h2h_hwdata [21]}),
    .f({_al_u1561_o,_al_u1562_o}),
    .q({freqB[15],freqB[21]}));  // src/AHB.v(57)
  // src/AHB.v(57)
  // src/AHB.v(57)
  EF2_PHY_MSLICE #(
    //.LUT0("(D*~C*~B*A)"),
    //.LUT1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000000000),
    .INIT_LUT1(16'b1000010000100001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg12_b16|U_AHB/reg12_b0  (
    .a({\PWMB/FreCnt [16],\U_AHB/h2h_hwrite }),
    .b({\PWMB/FreCnt [3],\U_AHB/h2h_haddr [13]}),
    .c({\PWMB/FreCntr [16],\U_AHB/h2h_haddr [14]}),
    .ce(\U_AHB/n26 ),
    .clk(clk100m),
    .d({\PWMB/FreCntr [3],\U_AHB/h2h_haddr [11]}),
    .mi({\U_AHB/h2h_hwdata [16],\U_AHB/h2h_hwdata [0]}),
    .f({_al_u1551_o,\U_AHB/n26 }),
    .q({freqB[16],freqB[0]}));  // src/AHB.v(57)
  // src/AHB.v(57)
  // src/AHB.v(57)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg12_b17|U_AHB/reg12_b22  (
    .a({open_n27287,_al_u1146_o}),
    .b({_al_u1145_o,\PWMB/FreCnt [2]}),
    .c({_al_u1147_o,\PWMB/FreCnt [20]}),
    .ce(\U_AHB/n26 ),
    .clk(clk100m),
    .d({_al_u1143_o,\PWMB/FreCnt [21]}),
    .e({open_n27288,\PWMB/FreCnt [22]}),
    .mi({\U_AHB/h2h_hwdata [17],\U_AHB/h2h_hwdata [22]}),
    .f({\PWMB/n0_lutinv ,_al_u1147_o}),
    .q({freqB[17],freqB[22]}));  // src/AHB.v(57)
  // src/AHB.v(57)
  // src/AHB.v(57)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg12_b19|U_AHB/reg12_b18  (
    .b({limit_l_pad[11],open_n27307}),
    .c({limit_r_pad[11],pwm_state_read[11]}),
    .ce(\U_AHB/n26 ),
    .clk(clk100m),
    .d({\PWMB/n11 ,\PWMB/n0_lutinv }),
    .mi(\U_AHB/h2h_hwdata [19:18]),
    .f({_al_u3041_o,\PWMB/n24 }),
    .q(freqB[19:18]));  // src/AHB.v(57)
  // src/AHB.v(57)
  // src/AHB.v(57)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~D*~C*~B*A)"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(~D*~C*~B*A)"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b0000000000000010),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg12_b20|U_AHB/reg12_b7  (
    .a({\PWMB/FreCnt [20],_al_u1142_o}),
    .b({\PWMB/FreCnt [26],\PWMB/FreCnt [7]}),
    .c({\PWMB/FreCntr [20],\PWMB/FreCnt [8]}),
    .ce(\U_AHB/n26 ),
    .clk(clk100m),
    .d({\PWMB/FreCntr [26],\PWMB/FreCnt [9]}),
    .mi({\U_AHB/h2h_hwdata [20],\U_AHB/h2h_hwdata [7]}),
    .f({_al_u1555_o,_al_u1143_o}),
    .q({freqB[20],freqB[7]}));  // src/AHB.v(57)
  // src/AHB.v(57)
  // src/AHB.v(57)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg12_b23|U_AHB/reg12_b3  (
    .a({\PWMB/FreCnt [23],_al_u1141_o}),
    .b({\PWMB/FreCnt [24],\PWMB/FreCnt [3]}),
    .c({\PWMB/FreCnt [25],\PWMB/FreCnt [4]}),
    .ce(\U_AHB/n26 ),
    .clk(clk100m),
    .d({\PWMB/FreCnt [26],\PWMB/FreCnt [5]}),
    .e({open_n27344,\PWMB/FreCnt [6]}),
    .mi({\U_AHB/h2h_hwdata [23],\U_AHB/h2h_hwdata [3]}),
    .f({_al_u1141_o,_al_u1142_o}),
    .q({freqB[23],freqB[3]}));  // src/AHB.v(57)
  // src/AHB.v(57)
  // src/AHB.v(57)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(D*~B)*~(~C*A))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(~(D*~B)*~(~C*A))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100010011110101),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1100010011110101),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg12_b24|U_AHB/reg12_b2  (
    .a({\PWMB/FreCnt [0],\PWMB/FreCnt [1]}),
    .b(\PWMB/FreCnt [24:23]),
    .c({\PWMB/FreCntr [0],\PWMB/FreCntr [2]}),
    .ce(\U_AHB/n26 ),
    .clk(clk100m),
    .d({\PWMB/FreCntr [24],\PWMB/FreCntr [24]}),
    .mi({\U_AHB/h2h_hwdata [24],\U_AHB/h2h_hwdata [2]}),
    .f({_al_u1559_o,_al_u2640_o}),
    .q({freqB[24],freqB[2]}));  // src/AHB.v(57)
  // src/AHB.v(57)
  // src/AHB.v(57)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C*D))"),
    //.LUT1("(C*~(A*~(D*B)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000110011001100),
    .INIT_LUT1(16'b1101000001010000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg12_b26|U_AHB/reg12_b5  (
    .a({_al_u3240_o,open_n27379}),
    .b({\U_AHB/n102 ,_al_u3061_o}),
    .c({_al_u3061_o,pwm_state_read[5]}),
    .ce(\U_AHB/n26 ),
    .clk(clk100m),
    .d({limit_l_pad[2],\U_AHB/n96 }),
    .mi({\U_AHB/h2h_hwdata [26],\U_AHB/h2h_hwdata [5]}),
    .f({_al_u3241_o,_al_u3139_o}),
    .q({freqB[26],freqB[5]}));  // src/AHB.v(57)
  // src/AHB.v(57)
  // src/AHB.v(57)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*~(~(0*B)*~(D*A)))"),
    //.LUTF1("(C*~(~(0*B)*~(D*A)))"),
    //.LUTG0("(C*~(~(1*B)*~(D*A)))"),
    //.LUTG1("(C*~(~(1*B)*~(D*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010000000000000),
    .INIT_LUTF1(16'b1010000000000000),
    .INIT_LUTG0(16'b1110000011000000),
    .INIT_LUTG1(16'b1110000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg12_b8|U_AHB/reg12_b9  (
    .a({\U_AHB/n96 ,\U_AHB/n96 }),
    .b({\U_AHB/n102 ,\U_AHB/n102 }),
    .c({_al_u3061_o,_al_u3061_o}),
    .ce(\U_AHB/n26 ),
    .clk(clk100m),
    .d({pwm_state_read[8],pwm_state_read[9]}),
    .e({limit_l_pad[8],limit_l_pad[9]}),
    .mi({\U_AHB/h2h_hwdata [8],\U_AHB/h2h_hwdata [9]}),
    .f({_al_u3080_o,_al_u3078_o}),
    .q({freqB[8],freqB[9]}));  // src/AHB.v(57)
  // src/AHB.v(58)
  // src/AHB.v(58)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg13_b10|U_AHB/reg13_b13  (
    .a({\PWMC/FreCnt [0],_al_u1576_o}),
    .b({\PWMC/FreCnt [10],\PWMC/FreCnt [13]}),
    .c({\PWMC/FreCntr [0],\PWMC/FreCnt [19]}),
    .ce(\U_AHB/n28 ),
    .clk(clk100m),
    .d({\PWMC/FreCntr [10],\PWMC/FreCntr [13]}),
    .e({open_n27410,\PWMC/FreCntr [19]}),
    .mi({\U_AHB/h2h_hwdata [10],\U_AHB/h2h_hwdata [13]}),
    .f({_al_u1576_o,_al_u1577_o}),
    .q({freqC[10],freqC[13]}));  // src/AHB.v(58)
  // src/AHB.v(58)
  // src/AHB.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~D*~C*B*A)"),
    //.LUT1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001000),
    .INIT_LUT1(16'b1000010000100001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg13_b11|U_AHB/reg13_b0  (
    .a({\PWMC/FreCnt [11],\U_AHB/h2h_hwrite }),
    .b({\PWMC/FreCnt [25],\U_AHB/h2h_haddr [12]}),
    .c({\PWMC/FreCntr [11],\U_AHB/h2h_haddr [13]}),
    .ce(\U_AHB/n28 ),
    .clk(clk100m),
    .d({\PWMC/FreCntr [25],\U_AHB/h2h_haddr [14]}),
    .mi({\U_AHB/h2h_hwdata [11],\U_AHB/h2h_hwdata [0]}),
    .f({_al_u1582_o,\U_AHB/n28 }),
    .q({freqC[11],freqC[0]}));  // src/AHB.v(58)
  // src/AHB.v(58)
  // src/AHB.v(58)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*B*A*~(0@D))"),
    //.LUTF1("(~(~D*B)*~(C*~A))"),
    //.LUTG0("(C*B*A*~(1@D))"),
    //.LUTG1("(~(~D*B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b1010111100100011),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b1010111100100011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg13_b15|U_AHB/reg13_b12  (
    .a({\PWMC/FreCnt [15],_al_u1575_o}),
    .b({\PWMC/FreCnt [21],_al_u1577_o}),
    .c({\PWMC/FreCntr [15],_al_u1578_o}),
    .ce(\U_AHB/n28 ),
    .clk(clk100m),
    .d({\PWMC/FreCntr [21],\PWMC/FreCnt [12]}),
    .e({open_n27441,\PWMC/FreCntr [12]}),
    .mi({\U_AHB/h2h_hwdata [15],\U_AHB/h2h_hwdata [12]}),
    .f({_al_u1578_o,_al_u1579_o}),
    .q({freqC[15],freqC[12]}));  // src/AHB.v(58)
  // src/AHB.v(58)
  // src/AHB.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b1000010000100001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg13_b17|U_AHB/reg13_b9  (
    .a({\PWMC/FreCnt [17],open_n27458}),
    .b({\PWMC/FreCnt [6],open_n27459}),
    .c({\PWMC/FreCntr [17],_al_u3061_o}),
    .ce(\U_AHB/n28 ),
    .clk(clk100m),
    .d({\PWMC/FreCntr [6],\U_AHB/n104_lutinv }),
    .mi({\U_AHB/h2h_hwdata [17],\U_AHB/h2h_hwdata [9]}),
    .f({_al_u1580_o,_al_u3065_o}),
    .q({freqC[17],freqC[9]}));  // src/AHB.v(58)
  // src/AHB.v(58)
  // src/AHB.v(58)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*~(~(0*B)*~(D*A)))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(C*~(~(1*B)*~(D*A)))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010000000000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b1110000011000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg13_b18|U_AHB/reg13_b5  (
    .a({open_n27474,\U_AHB/n96 }),
    .b({limit_l_pad[12],\U_AHB/n102 }),
    .c({limit_r_pad[12],_al_u3061_o}),
    .ce(\U_AHB/n28 ),
    .clk(clk100m),
    .d({\PWMC/n11 ,pwm_state_read[12]}),
    .e({open_n27475,limit_l_pad[12]}),
    .mi({\U_AHB/h2h_hwdata [18],\U_AHB/h2h_hwdata [5]}),
    .f({_al_u3044_o,_al_u3072_o}),
    .q({freqC[18],freqC[5]}));  // src/AHB.v(58)
  // src/AHB.v(58)
  // src/AHB.v(58)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg13_b19|U_AHB/reg13_b22  (
    .a({\PWMC/FreCnt [16],_al_u1183_o}),
    .b({\PWMC/FreCnt [17],\PWMC/FreCnt [2]}),
    .c({\PWMC/FreCnt [18],\PWMC/FreCnt [20]}),
    .ce(\U_AHB/n28 ),
    .clk(clk100m),
    .d({\PWMC/FreCnt [19],\PWMC/FreCnt [21]}),
    .e({open_n27492,\PWMC/FreCnt [22]}),
    .mi({\U_AHB/h2h_hwdata [19],\U_AHB/h2h_hwdata [22]}),
    .f({_al_u1183_o,_al_u1184_o}),
    .q({freqC[19],freqC[22]}));  // src/AHB.v(58)
  // src/AHB.v(58)
  // src/AHB.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(D*~B)*~(~C*A))"),
    //.LUT1("(D*~(C@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100010011110101),
    .INIT_LUT1(16'b1100001100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg13_b1|U_AHB/reg13_b21  (
    .a({open_n27509,\PWMC/FreCnt [15]}),
    .b({\PWMC/FreCnt [1],\PWMC/FreCnt [21]}),
    .c({\PWMC/FreCntr [1],\PWMC/FreCntr [15]}),
    .ce(\U_AHB/n28 ),
    .clk(clk100m),
    .d({_al_u1574_o,\PWMC/FreCntr [21]}),
    .mi({\U_AHB/h2h_hwdata [1],\U_AHB/h2h_hwdata [21]}),
    .f({_al_u1575_o,_al_u1574_o}),
    .q({freqC[1],freqC[21]}));  // src/AHB.v(58)
  // src/AHB.v(58)
  // src/AHB.v(58)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(~0*C)*~(D*~B))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(A*~(~1*C)*~(D*~B))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000001010),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000100010101010),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg13_b20|U_AHB/reg13_b16  (
    .a({\PWMC/FreCnt [20],_al_u2720_o}),
    .b({\PWMC/FreCnt [26],\PWMC/FreCnt [15]}),
    .c({\PWMC/FreCntr [20],\PWMC/FreCnt [19]}),
    .ce(\U_AHB/n28 ),
    .clk(clk100m),
    .d({\PWMC/FreCntr [26],\PWMC/FreCntr [16]}),
    .e({open_n27524,\PWMC/FreCntr [20]}),
    .mi({\U_AHB/h2h_hwdata [20],\U_AHB/h2h_hwdata [16]}),
    .f({_al_u1572_o,_al_u2721_o}),
    .q({freqC[20],freqC[16]}));  // src/AHB.v(58)
  // src/AHB.v(58)
  // src/AHB.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~D*~C*~B*A)"),
    //.LUT1("(B*A*~(D*~C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000010),
    .INIT_LUT1(16'b1000000010001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg13_b23|U_AHB/reg13_b7  (
    .a({_al_u2717_o,_al_u1179_o}),
    .b({_al_u2718_o,\PWMC/FreCnt [7]}),
    .c({\PWMC/FreCnt [23],\PWMC/FreCnt [8]}),
    .ce(\U_AHB/n28 ),
    .clk(clk100m),
    .d({\PWMC/FreCntr [24],\PWMC/FreCnt [9]}),
    .mi({\U_AHB/h2h_hwdata [23],\U_AHB/h2h_hwdata [7]}),
    .f({_al_u2719_o,_al_u1180_o}),
    .q({freqC[23],freqC[7]}));  // src/AHB.v(58)
  // src/AHB.v(58)
  // src/AHB.v(58)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg13_b24|U_AHB/reg13_b3  (
    .a({\PWMC/FreCnt [23],_al_u1178_o}),
    .b({\PWMC/FreCnt [24],\PWMC/FreCnt [3]}),
    .c({\PWMC/FreCnt [25],\PWMC/FreCnt [4]}),
    .ce(\U_AHB/n28 ),
    .clk(clk100m),
    .d({\PWMC/FreCnt [26],\PWMC/FreCnt [5]}),
    .e({open_n27555,\PWMC/FreCnt [6]}),
    .mi({\U_AHB/h2h_hwdata [24],\U_AHB/h2h_hwdata [3]}),
    .f({_al_u1178_o,_al_u1179_o}),
    .q({freqC[24],freqC[3]}));  // src/AHB.v(58)
  // src/AHB.v(58)
  // src/AHB.v(58)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*~(~(0*B)*~(D*A)))"),
    //.LUTF1("(C*~(~(0*B)*~(D*A)))"),
    //.LUTG0("(C*~(~(1*B)*~(D*A)))"),
    //.LUTG1("(C*~(~(1*B)*~(D*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010000000000000),
    .INIT_LUTF1(16'b1010000000000000),
    .INIT_LUTG0(16'b1110000011000000),
    .INIT_LUTG1(16'b1110000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg13_b26|U_AHB/reg13_b8  (
    .a({\U_AHB/n96 ,\U_AHB/n96 }),
    .b({\U_AHB/n102 ,\U_AHB/n102 }),
    .c({_al_u3061_o,_al_u3061_o}),
    .ce(\U_AHB/n28 ),
    .clk(clk100m),
    .d({pwm_state_read[10],pwm_state_read[14]}),
    .e({limit_l_pad[10],limit_l_pad[14]}),
    .mi({\U_AHB/h2h_hwdata [26],\U_AHB/h2h_hwdata [8]}),
    .f({_al_u3076_o,_al_u3068_o}),
    .q({freqC[26],freqC[8]}));  // src/AHB.v(58)
  // src/AHB.v(58)
  // src/AHB.v(58)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*~(~(0*B)*~(D*A)))"),
    //.LUTF1("(C*~(~(0*B)*~(D*A)))"),
    //.LUTG0("(C*~(~(1*B)*~(D*A)))"),
    //.LUTG1("(C*~(~(1*B)*~(D*A)))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010000000000000),
    .INIT_LUTF1(16'b1010000000000000),
    .INIT_LUTG0(16'b1110000011000000),
    .INIT_LUTG1(16'b1110000011000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg13_b4|U_AHB/reg13_b6  (
    .a({\U_AHB/n96 ,\U_AHB/n96 }),
    .b({\U_AHB/n102 ,\U_AHB/n102 }),
    .c({_al_u3061_o,_al_u3061_o}),
    .ce(\U_AHB/n28 ),
    .clk(clk100m),
    .d({pwm_state_read[11],pwm_state_read[13]}),
    .e({limit_l_pad[11],limit_l_pad[13]}),
    .mi({\U_AHB/h2h_hwdata [4],\U_AHB/h2h_hwdata [6]}),
    .f({_al_u3074_o,_al_u3070_o}),
    .q({freqC[4],freqC[6]}));  // src/AHB.v(58)
  // src/AHB.v(60)
  // src/AHB.v(60)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~((0*C)*~(B)*~(D)+(0*C)*B*~(D)+~((0*C))*B*D+(0*C)*B*D))"),
    //.LUTF1("(~D*C*B*A)"),
    //.LUTG0("(A*~((1*C)*~(B)*~(D)+(1*C)*B*~(D)+~((1*C))*B*D+(1*C)*B*D))"),
    //.LUTG1("(~D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b0010001000001010),
    .INIT_LUTG1(16'b0000000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg14_b0|U_AHB/reg14_b1  (
    .a({\U_AHB/h2h_hwrite ,_al_u3061_o}),
    .b({\U_AHB/h2h_haddr [2],pnumcntB[0]}),
    .c({\U_AHB/h2h_haddr [13],pnumcntC[0]}),
    .ce(\U_AHB/n30 ),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [14],\U_AHB/h2h_haddr [2]}),
    .e({open_n27604,\U_AHB/h2h_haddr [3]}),
    .mi({\U_AHB/h2h_hwdata [0],\U_AHB/h2h_hwdata [1]}),
    .f({\U_AHB/n30 ,_al_u3349_o}),
    .q({freqD[0],freqD[1]}));  // src/AHB.v(60)
  // src/AHB.v(60)
  // src/AHB.v(60)
  EF2_PHY_MSLICE #(
    //.LUT0("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    //.LUT1("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101001101011111),
    .INIT_LUT1(16'b0101001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg14_b12|U_AHB/reg14_b10  (
    .a(pnumcnt0[1:0]),
    .b(pnumcnt1[1:0]),
    .c({\U_AHB/h2h_haddr [2],\U_AHB/h2h_haddr [2]}),
    .ce(\U_AHB/n30 ),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [3],\U_AHB/h2h_haddr [3]}),
    .mi({\U_AHB/h2h_hwdata [12],\U_AHB/h2h_hwdata [10]}),
    .f({_al_u3332_o,_al_u3343_o}),
    .q({freqD[12],freqD[10]}));  // src/AHB.v(60)
  // src/AHB.v(60)
  // src/AHB.v(60)
  EF2_PHY_MSLICE #(
    //.LUT0("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    //.LUT1("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101001101011111),
    .INIT_LUT1(16'b0101001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg14_b14|U_AHB/reg14_b8  (
    .a({pnumcnt0[10],pnumcnt0[2]}),
    .b({pnumcnt1[10],pnumcnt1[2]}),
    .c({\U_AHB/h2h_haddr [2],\U_AHB/h2h_haddr [2]}),
    .ce(\U_AHB/n30 ),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [3],\U_AHB/h2h_haddr [3]}),
    .mi({\U_AHB/h2h_hwdata [14],\U_AHB/h2h_hwdata [8]}),
    .f({_al_u3321_o,_al_u3211_o}),
    .q({freqD[14],freqD[8]}));  // src/AHB.v(60)
  // src/AHB.v(60)
  // src/AHB.v(60)
  EF2_PHY_MSLICE #(
    //.LUT0("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    //.LUT1("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101001101011111),
    .INIT_LUT1(16'b0101001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg14_b16|U_AHB/reg14_b3  (
    .a({pnumcnt0[11],pnumcnt0[17]}),
    .b({pnumcnt1[11],pnumcnt1[17]}),
    .c({\U_AHB/h2h_haddr [2],\U_AHB/h2h_haddr [2]}),
    .ce(\U_AHB/n30 ),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [3],\U_AHB/h2h_haddr [3]}),
    .mi({\U_AHB/h2h_hwdata [16],\U_AHB/h2h_hwdata [3]}),
    .f({_al_u3310_o,_al_u3244_o}),
    .q({freqD[16],freqD[3]}));  // src/AHB.v(60)
  // src/AHB.v(60)
  // src/AHB.v(60)
  EF2_PHY_MSLICE #(
    //.LUT0("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    //.LUT1("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101001101011111),
    .INIT_LUT1(16'b0101001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg14_b18|U_AHB/reg14_b25  (
    .a({pnumcnt0[12],pnumcnt0[16]}),
    .b({pnumcnt1[12],pnumcnt1[16]}),
    .c({\U_AHB/h2h_haddr [2],\U_AHB/h2h_haddr [2]}),
    .ce(\U_AHB/n30 ),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [3],\U_AHB/h2h_haddr [3]}),
    .mi({\U_AHB/h2h_hwdata [18],\U_AHB/h2h_hwdata [25]}),
    .f({_al_u3299_o,_al_u3255_o}),
    .q({freqD[18],freqD[25]}));  // src/AHB.v(60)
  // src/AHB.v(60)
  // src/AHB.v(60)
  EF2_PHY_MSLICE #(
    //.LUT0("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    //.LUT1("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101001101011111),
    .INIT_LUT1(16'b0101001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg14_b21|U_AHB/reg14_b23  (
    .a({pnumcnt0[14],pnumcnt0[15]}),
    .b({pnumcnt1[14],pnumcnt1[15]}),
    .c({\U_AHB/h2h_haddr [2],\U_AHB/h2h_haddr [2]}),
    .ce(\U_AHB/n30 ),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [3],\U_AHB/h2h_haddr [3]}),
    .mi({\U_AHB/h2h_hwdata [21],\U_AHB/h2h_hwdata [23]}),
    .f({_al_u3277_o,_al_u3266_o}),
    .q({freqD[21],freqD[23]}));  // src/AHB.v(60)
  // src/AHB.v(61)
  // src/AHB.v(61)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~((0*C)*~(B)*~(D)+(0*C)*B*~(D)+~((0*C))*B*D+(0*C)*B*D))"),
    //.LUTF1("(~D*C*B*A)"),
    //.LUTG0("(A*~((1*C)*~(B)*~(D)+(1*C)*B*~(D)+~((1*C))*B*D+(1*C)*B*D))"),
    //.LUTG1("(~D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b0010001000001010),
    .INIT_LUTG1(16'b0000000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg15_b0|U_AHB/reg15_b3  (
    .a({\U_AHB/h2h_hwrite ,_al_u3061_o}),
    .b({\U_AHB/h2h_haddr [3],pnumcntB[9]}),
    .c({\U_AHB/h2h_haddr [13],pnumcntC[9]}),
    .ce(\U_AHB/n32 ),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [14],\U_AHB/h2h_haddr [2]}),
    .e({open_n27691,\U_AHB/h2h_haddr [3]}),
    .mi({\U_AHB/h2h_hwdata [0],\U_AHB/h2h_hwdata [3]}),
    .f({\U_AHB/n32 ,_al_u3095_o}),
    .q({freqE[0],freqE[3]}));  // src/AHB.v(61)
  // src/AHB.v(61)
  // src/AHB.v(61)
  EF2_PHY_MSLICE #(
    //.LUT0("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    //.LUT1("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101001101011111),
    .INIT_LUT1(16'b0101001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg15_b10|U_AHB/reg15_b7  (
    .a({pnumcntB[21],pnumcnt0[9]}),
    .b({pnumcntC[21],pnumcnt1[9]}),
    .c({\U_AHB/h2h_haddr [2],\U_AHB/h2h_haddr [2]}),
    .ce(\U_AHB/n32 ),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [3],\U_AHB/h2h_haddr [3]}),
    .mi({\U_AHB/h2h_hwdata [10],\U_AHB/h2h_hwdata [7]}),
    .f({_al_u3195_o,_al_u3082_o}),
    .q({freqE[10],freqE[7]}));  // src/AHB.v(61)
  // src/AHB.v(61)
  // src/AHB.v(61)
  EF2_PHY_MSLICE #(
    //.LUT0("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    //.LUT1("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101001101011111),
    .INIT_LUT1(16'b0101001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg15_b11|U_AHB/reg15_b26  (
    .a({pnumcnt0[21],pnumcnt0[8]}),
    .b({pnumcnt1[21],pnumcnt1[8]}),
    .c({\U_AHB/h2h_haddr [2],\U_AHB/h2h_haddr [2]}),
    .ce(\U_AHB/n32 ),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [3],\U_AHB/h2h_haddr [3]}),
    .mi({\U_AHB/h2h_hwdata [11],\U_AHB/h2h_hwdata [26]}),
    .f({_al_u3189_o,_al_u3100_o}),
    .q({freqE[11],freqE[26]}));  // src/AHB.v(61)
  // src/AHB.v(61)
  // src/AHB.v(61)
  EF2_PHY_MSLICE #(
    //.LUT0("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    //.LUT1("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101001101011111),
    .INIT_LUT1(16'b0101001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg15_b13|U_AHB/reg15_b24  (
    .a({pnumcnt0[22],pnumcnt0[7]}),
    .b({pnumcnt1[22],pnumcnt1[7]}),
    .c({\U_AHB/h2h_haddr [2],\U_AHB/h2h_haddr [2]}),
    .ce(\U_AHB/n32 ),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [3],\U_AHB/h2h_haddr [3]}),
    .mi({\U_AHB/h2h_hwdata [13],\U_AHB/h2h_hwdata [24]}),
    .f({_al_u3178_o,_al_u3111_o}),
    .q({freqE[13],freqE[24]}));  // src/AHB.v(61)
  // src/AHB.v(61)
  // src/AHB.v(61)
  EF2_PHY_MSLICE #(
    //.LUT0("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    //.LUT1("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101001101011111),
    .INIT_LUT1(16'b0101001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg15_b15|U_AHB/reg15_b22  (
    .a({pnumcnt0[23],pnumcnt0[6]}),
    .b({pnumcnt1[23],pnumcnt1[6]}),
    .c({\U_AHB/h2h_haddr [2],\U_AHB/h2h_haddr [2]}),
    .ce(\U_AHB/n32 ),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [3],\U_AHB/h2h_haddr [3]}),
    .mi({\U_AHB/h2h_hwdata [15],\U_AHB/h2h_hwdata [22]}),
    .f({_al_u3167_o,_al_u3122_o}),
    .q({freqE[15],freqE[22]}));  // src/AHB.v(61)
  // src/AHB.v(61)
  // src/AHB.v(61)
  EF2_PHY_MSLICE #(
    //.LUT0("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    //.LUT1("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101001101011111),
    .INIT_LUT1(16'b0101001101011111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg15_b1|U_AHB/reg15_b17  (
    .a({pnumcnt0[20],pnumcnt0[3]}),
    .b({pnumcnt1[20],pnumcnt1[3]}),
    .c({\U_AHB/h2h_haddr [2],\U_AHB/h2h_haddr [2]}),
    .ce(\U_AHB/n32 ),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [3],\U_AHB/h2h_haddr [3]}),
    .mi({\U_AHB/h2h_hwdata [1],\U_AHB/h2h_hwdata [17]}),
    .f({_al_u3200_o,_al_u3156_o}),
    .q({freqE[1],freqE[17]}));  // src/AHB.v(61)
  // src/AHB.v(61)
  // src/AHB.v(61)
  EF2_PHY_MSLICE #(
    //.LUT0("(D*~C*~B*~A)"),
    //.LUT1("(C*~B*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000100000000),
    .INIT_LUT1(16'b0000000000110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg15_b5|U_AHB/reg15_b6  (
    .a({open_n27778,\U_AHB/h2h_haddr [2]}),
    .b({\U_AHB/h2h_haddr [3],\U_AHB/h2h_haddr [3]}),
    .c({\U_AHB/h2h_haddr [4],\U_AHB/h2h_haddr [4]}),
    .ce(\U_AHB/n32 ),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [2],\U_AHB/h2h_haddr [5]}),
    .mi({\U_AHB/h2h_hwdata [5],\U_AHB/h2h_hwdata [6]}),
    .f({\U_AHB/n87 ,\U_AHB/n90 }),
    .q({freqE[5],freqE[6]}));  // src/AHB.v(61)
  // src/AHB.v(61)
  // src/AHB.v(61)
  EF2_PHY_LSLICE #(
    //.LUTF0("(0*~D*~C*~B*~A)"),
    //.LUTF1("(~0*~D*~C*~B*~A)"),
    //.LUTG0("(1*~D*~C*~B*~A)"),
    //.LUTG1("(~1*~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000000000000001),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg15_b8|U_AHB/reg15_b4  (
    .a({\U_AHB/h2h_haddr [2],\U_AHB/h2h_haddr [2]}),
    .b({\U_AHB/h2h_haddr [3],\U_AHB/h2h_haddr [3]}),
    .c({\U_AHB/h2h_haddr [4],\U_AHB/h2h_haddr [4]}),
    .ce(\U_AHB/n32 ),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [5],\U_AHB/h2h_haddr [5]}),
    .e({\U_AHB/h2h_haddr [6],\U_AHB/h2h_haddr [6]}),
    .mi({\U_AHB/h2h_hwdata [8],\U_AHB/h2h_hwdata [4]}),
    .f({\U_AHB/n95_lutinv ,\U_AHB/n93 }),
    .q({freqE[8],freqE[4]}));  // src/AHB.v(61)
  // src/AHB.v(62)
  // src/AHB.v(62)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(D*~C*B*A)"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(D*~C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b0000100000000000),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b0000100000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg16_b0|U_AHB/reg16_b17  (
    .a({\U_AHB/h2h_hwrite ,_al_u1620_o}),
    .b({\U_AHB/h2h_haddr [13],\PWMF/FreCnt [17]}),
    .c({\U_AHB/h2h_haddr [14],\PWMF/FreCnt [8]}),
    .ce(\U_AHB/n34 ),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [4],\PWMF/FreCntr [17]}),
    .e({open_n27809,\PWMF/FreCntr [8]}),
    .mi({\U_AHB/h2h_hwdata [0],\U_AHB/h2h_hwdata [17]}),
    .f({\U_AHB/n34 ,_al_u1621_o}),
    .q({freqF[0],freqF[17]}));  // src/AHB.v(62)
  // src/AHB.v(62)
  // src/AHB.v(62)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1000010000100001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg16_b10|U_AHB/reg16_b19  (
    .a({\PWMF/FreCnt [10],open_n27826}),
    .b({\PWMF/FreCnt [2],open_n27827}),
    .c({\PWMF/FreCntr [10],pwm_state_read[15]}),
    .ce(\U_AHB/n34 ),
    .clk(clk100m),
    .d({\PWMF/FreCntr [2],\PWMF/n0_lutinv }),
    .mi({\U_AHB/h2h_hwdata [10],\U_AHB/h2h_hwdata [19]}),
    .f({_al_u1627_o,\PWMF/n24 }),
    .q({freqF[10],freqF[19]}));  // src/AHB.v(62)
  // src/AHB.v(62)
  // src/AHB.v(62)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(D*~B)*~(C*~A))"),
    //.LUT1("(~(~D*B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000110010101111),
    .INIT_LUT1(16'b1111010100110001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg16_b14|U_AHB/reg16_b15  (
    .a(\PWMF/FreCnt [13:12]),
    .b({\PWMF/FreCnt [23],\PWMF/FreCnt [15]}),
    .c({\PWMF/FreCntr [14],\PWMF/FreCntr [12]}),
    .ce(\U_AHB/n34 ),
    .clk(clk100m),
    .d({\PWMF/FreCntr [24],\PWMF/FreCntr [15]}),
    .mi({\U_AHB/h2h_hwdata [14],\U_AHB/h2h_hwdata [15]}),
    .f({_al_u2967_o,_al_u1626_o}),
    .q({freqF[14],freqF[15]}));  // src/AHB.v(62)
  // src/AHB.v(62)
  // src/AHB.v(62)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg16_b16|U_AHB/reg16_b13  (
    .a({\PWMF/FreCnt [16],_al_u1635_o}),
    .b({\PWMF/FreCnt [26],\PWMF/FreCnt [13]}),
    .c({\PWMF/FreCntr [16],\PWMF/FreCnt [19]}),
    .ce(\U_AHB/n34 ),
    .clk(clk100m),
    .d({\PWMF/FreCntr [26],\PWMF/FreCntr [13]}),
    .e({open_n27856,\PWMF/FreCntr [19]}),
    .mi({\U_AHB/h2h_hwdata [16],\U_AHB/h2h_hwdata [13]}),
    .f({_al_u1635_o,_al_u1636_o}),
    .q({freqF[16],freqF[13]}));  // src/AHB.v(62)
  // src/AHB.v(62)
  // src/AHB.v(62)
  EF2_PHY_MSLICE #(
    //.LUT0("(~D*~C*~B*~A)"),
    //.LUT1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000001),
    .INIT_LUT1(16'b1000010000100001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg16_b18|U_AHB/reg16_b26  (
    .a({\PWMF/FreCnt [18],pnumcntC[18]}),
    .b({\PWMF/FreCnt [5],pnumcntC[19]}),
    .c({\PWMF/FreCntr [18],pnumcntC[1]}),
    .ce(\U_AHB/n34 ),
    .clk(clk100m),
    .d({\PWMF/FreCntr [5],pnumcntC[20]}),
    .mi({\U_AHB/h2h_hwdata [18],\U_AHB/h2h_hwdata [26]}),
    .f({_al_u1624_o,_al_u2661_o}),
    .q({freqF[18],freqF[26]}));  // src/AHB.v(62)
  // src/AHB.v(62)
  // src/AHB.v(62)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg16_b23|U_AHB/reg16_b3  (
    .a({\PWMF/FreCnt [23],_al_u1289_o}),
    .b({\PWMF/FreCnt [24],\PWMF/FreCnt [3]}),
    .c({\PWMF/FreCnt [25],\PWMF/FreCnt [4]}),
    .ce(\U_AHB/n34 ),
    .clk(clk100m),
    .d({\PWMF/FreCnt [26],\PWMF/FreCnt [5]}),
    .e({open_n27887,\PWMF/FreCnt [6]}),
    .mi({\U_AHB/h2h_hwdata [23],\U_AHB/h2h_hwdata [3]}),
    .f({_al_u1289_o,_al_u1290_o}),
    .q({freqF[23],freqF[3]}));  // src/AHB.v(62)
  // src/AHB.v(62)
  // src/AHB.v(62)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg16_b25|U_AHB/reg16_b20  (
    .a({\PWMF/FreCnt [11],_al_u1633_o}),
    .b({\PWMF/FreCnt [25],\PWMF/FreCnt [14]}),
    .c({\PWMF/FreCntr [11],\PWMF/FreCnt [20]}),
    .ce(\U_AHB/n34 ),
    .clk(clk100m),
    .d({\PWMF/FreCntr [25],\PWMF/FreCntr [14]}),
    .e({open_n27904,\PWMF/FreCntr [20]}),
    .mi({\U_AHB/h2h_hwdata [25],\U_AHB/h2h_hwdata [20]}),
    .f({_al_u1633_o,_al_u1634_o}),
    .q({freqF[25],freqF[20]}));  // src/AHB.v(62)
  // src/AHB.v(62)
  // src/AHB.v(62)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*~(~(0*B)*~(D*A)))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(C*~(~(1*B)*~(D*A)))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010000000000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b1110000011000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg16_b2|U_AHB/reg16_b22  (
    .a({open_n27921,\U_AHB/n96 }),
    .b({limit_l_pad[15],\U_AHB/n102 }),
    .c({limit_r_pad[15],_al_u3061_o}),
    .ce(\U_AHB/n34 ),
    .clk(clk100m),
    .d({\PWMF/n11 ,pwm_state_read[15]}),
    .e({open_n27922,limit_l_pad[15]}),
    .mi({\U_AHB/h2h_hwdata [2],\U_AHB/h2h_hwdata [22]}),
    .f({_al_u3053_o,_al_u3062_o}),
    .q({freqF[2],freqF[22]}));  // src/AHB.v(62)
  // src/AHB.v(62)
  // src/AHB.v(62)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(~D*~C*~B*A)"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(~D*~C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b0000000000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg16_b7|U_AHB/reg16_b4  (
    .a({_al_u1290_o,_al_u1622_o}),
    .b({\PWMF/FreCnt [7],\PWMF/FreCnt [4]}),
    .c({\PWMF/FreCnt [8],\PWMF/FreCnt [9]}),
    .ce(\U_AHB/n34 ),
    .clk(clk100m),
    .d({\PWMF/FreCnt [9],\PWMF/FreCntr [4]}),
    .e({open_n27939,\PWMF/FreCntr [9]}),
    .mi({\U_AHB/h2h_hwdata [7],\U_AHB/h2h_hwdata [4]}),
    .f({_al_u1291_o,_al_u1623_o}),
    .q({freqF[7],freqF[4]}));  // src/AHB.v(62)
  // src/AHB.v(64)
  // src/AHB.v(64)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUT1("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1101110011110000),
    .INIT_LUT1(16'b1101110011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg17_b0|U_AHB/reg17_b9  (
    .a({\U_AHB/n38 ,\U_AHB/n38 }),
    .b({\U_AHB/n36 ,\U_AHB/n36 }),
    .c({gpio_out_pad[0],gpio_out_pad[9]}),
    .clk(clk100m),
    .d({\U_AHB/h2h_hwdata [0],\U_AHB/h2h_hwdata [9]}),
    .q({gpio_out_pad[0],gpio_out_pad[9]}));  // src/AHB.v(64)
  // src/AHB.v(64)
  // src/AHB.v(64)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUT1("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1101110011110000),
    .INIT_LUT1(16'b1101110011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg17_b10|U_AHB/reg17_b8  (
    .a({\U_AHB/n38 ,\U_AHB/n38 }),
    .b({\U_AHB/n36 ,\U_AHB/n36 }),
    .c({gpio_out_pad[10],gpio_out_pad[8]}),
    .clk(clk100m),
    .d({\U_AHB/h2h_hwdata [10],\U_AHB/h2h_hwdata [8]}),
    .q({gpio_out_pad[10],gpio_out_pad[8]}));  // src/AHB.v(64)
  // src/AHB.v(64)
  // src/AHB.v(64)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTF1("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG0("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG1("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101110011110000),
    .INIT_LUTF1(16'b1101110011110000),
    .INIT_LUTG0(16'b1101110011110000),
    .INIT_LUTG1(16'b1101110011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg17_b11|U_AHB/reg17_b7  (
    .a({\U_AHB/n38 ,\U_AHB/n38 }),
    .b({\U_AHB/n36 ,\U_AHB/n36 }),
    .c({gpio_out_pad[11],gpio_out_pad[7]}),
    .clk(clk100m),
    .d({\U_AHB/h2h_hwdata [11],\U_AHB/h2h_hwdata [7]}),
    .q({gpio_out_pad[11],gpio_out_pad[7]}));  // src/AHB.v(64)
  // src/AHB.v(64)
  // src/AHB.v(64)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTF1("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG0("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG1("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101110011110000),
    .INIT_LUTF1(16'b1101110011110000),
    .INIT_LUTG0(16'b1101110011110000),
    .INIT_LUTG1(16'b1101110011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg17_b12|U_AHB/reg17_b6  (
    .a({\U_AHB/n38 ,\U_AHB/n38 }),
    .b({\U_AHB/n36 ,\U_AHB/n36 }),
    .c({gpio_out_pad[12],gpio_out_pad[6]}),
    .clk(clk100m),
    .d({\U_AHB/h2h_hwdata [12],\U_AHB/h2h_hwdata [6]}),
    .q({gpio_out_pad[12],gpio_out_pad[6]}));  // src/AHB.v(64)
  // src/AHB.v(64)
  // src/AHB.v(64)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUT1("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1101110011110000),
    .INIT_LUT1(16'b1101110011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg17_b13|U_AHB/reg17_b5  (
    .a({\U_AHB/n38 ,\U_AHB/n38 }),
    .b({\U_AHB/n36 ,\U_AHB/n36 }),
    .c({gpio_out_pad[13],gpio_out_pad[5]}),
    .clk(clk100m),
    .d({\U_AHB/h2h_hwdata [13],\U_AHB/h2h_hwdata [5]}),
    .q({gpio_out_pad[13],gpio_out_pad[5]}));  // src/AHB.v(64)
  // src/AHB.v(64)
  // src/AHB.v(64)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUT1("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1101110011110000),
    .INIT_LUT1(16'b1101110011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg17_b14|U_AHB/reg17_b4  (
    .a({\U_AHB/n38 ,\U_AHB/n38 }),
    .b({\U_AHB/n36 ,\U_AHB/n36 }),
    .c({gpio_out_pad[14],gpio_out_pad[4]}),
    .clk(clk100m),
    .d({\U_AHB/h2h_hwdata [14],\U_AHB/h2h_hwdata [4]}),
    .q({gpio_out_pad[14],gpio_out_pad[4]}));  // src/AHB.v(64)
  // src/AHB.v(64)
  // src/AHB.v(64)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTF1("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG0("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG1("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101110011110000),
    .INIT_LUTF1(16'b1101110011110000),
    .INIT_LUTG0(16'b1101110011110000),
    .INIT_LUTG1(16'b1101110011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg17_b15|U_AHB/reg17_b3  (
    .a({\U_AHB/n38 ,\U_AHB/n38 }),
    .b({\U_AHB/n36 ,\U_AHB/n36 }),
    .c({gpio_out_pad[15],gpio_out_pad[3]}),
    .clk(clk100m),
    .d({\U_AHB/h2h_hwdata [15],\U_AHB/h2h_hwdata [3]}),
    .q({gpio_out_pad[15],gpio_out_pad[3]}));  // src/AHB.v(64)
  // src/AHB.v(64)
  // src/AHB.v(64)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTF1("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG0("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG1("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101110011110000),
    .INIT_LUTF1(16'b1101110011110000),
    .INIT_LUTG0(16'b1101110011110000),
    .INIT_LUTG1(16'b1101110011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg17_b16|U_AHB/reg17_b26  (
    .a({\U_AHB/n38 ,\U_AHB/n38 }),
    .b({\U_AHB/n36 ,\U_AHB/n36 }),
    .c({gpio_out_pad[16],gpio_out_pad[26]}),
    .clk(clk100m),
    .d({\U_AHB/h2h_hwdata [16],\U_AHB/h2h_hwdata [26]}),
    .q({gpio_out_pad[16],gpio_out_pad[26]}));  // src/AHB.v(64)
  // src/AHB.v(64)
  // src/AHB.v(64)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUT1("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1101110011110000),
    .INIT_LUT1(16'b1101110011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg17_b17|U_AHB/reg17_b25  (
    .a({\U_AHB/n38 ,\U_AHB/n38 }),
    .b({\U_AHB/n36 ,\U_AHB/n36 }),
    .c({gpio_out_pad[17],gpio_out_pad[25]}),
    .clk(clk100m),
    .d({\U_AHB/h2h_hwdata [17],\U_AHB/h2h_hwdata [25]}),
    .q({gpio_out_pad[17],gpio_out_pad[25]}));  // src/AHB.v(64)
  // src/AHB.v(64)
  // src/AHB.v(64)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUT1("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1101110011110000),
    .INIT_LUT1(16'b1101110011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg17_b18|U_AHB/reg17_b24  (
    .a({\U_AHB/n38 ,\U_AHB/n38 }),
    .b({\U_AHB/n36 ,\U_AHB/n36 }),
    .c({gpio_out_pad[18],gpio_out_pad[24]}),
    .clk(clk100m),
    .d({\U_AHB/h2h_hwdata [18],\U_AHB/h2h_hwdata [24]}),
    .q({gpio_out_pad[18],gpio_out_pad[24]}));  // src/AHB.v(64)
  // src/AHB.v(64)
  // src/AHB.v(64)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTF1("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG0("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG1("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101110011110000),
    .INIT_LUTF1(16'b1101110011110000),
    .INIT_LUTG0(16'b1101110011110000),
    .INIT_LUTG1(16'b1101110011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg17_b19|U_AHB/reg17_b23  (
    .a({\U_AHB/n38 ,\U_AHB/n38 }),
    .b({\U_AHB/n36 ,\U_AHB/n36 }),
    .c({gpio_out_pad[19],gpio_out_pad[23]}),
    .clk(clk100m),
    .d({\U_AHB/h2h_hwdata [19],\U_AHB/h2h_hwdata [23]}),
    .q({gpio_out_pad[19],gpio_out_pad[23]}));  // src/AHB.v(64)
  // src/AHB.v(64)
  // src/AHB.v(64)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTF1("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG0("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG1("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101110011110000),
    .INIT_LUTF1(16'b1101110011110000),
    .INIT_LUTG0(16'b1101110011110000),
    .INIT_LUTG1(16'b1101110011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg17_b1|U_AHB/reg17_b22  (
    .a({\U_AHB/n38 ,\U_AHB/n38 }),
    .b({\U_AHB/n36 ,\U_AHB/n36 }),
    .c({gpio_out_pad[1],gpio_out_pad[22]}),
    .clk(clk100m),
    .d({\U_AHB/h2h_hwdata [1],\U_AHB/h2h_hwdata [22]}),
    .q({gpio_out_pad[1],gpio_out_pad[22]}));  // src/AHB.v(64)
  // src/AHB.v(64)
  // src/AHB.v(64)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUT1("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1101110011110000),
    .INIT_LUT1(16'b1101110011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg17_b20|U_AHB/reg17_b21  (
    .a({\U_AHB/n38 ,\U_AHB/n38 }),
    .b({\U_AHB/n36 ,\U_AHB/n36 }),
    .c({gpio_out_pad[20],gpio_out_pad[21]}),
    .clk(clk100m),
    .d({\U_AHB/h2h_hwdata [20],\U_AHB/h2h_hwdata [21]}),
    .q({gpio_out_pad[20],gpio_out_pad[21]}));  // src/AHB.v(64)
  // src/AHB.v(64)
  // src/AHB.v(64)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUT1("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1101110011110000),
    .INIT_LUT1(16'b1101110011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg17_b27|U_AHB/reg17_b2  (
    .a({\U_AHB/n38 ,\U_AHB/n38 }),
    .b({\U_AHB/n36 ,\U_AHB/n36 }),
    .c({gpio_out_pad[27],gpio_out_pad[2]}),
    .clk(clk100m),
    .d({\U_AHB/h2h_hwdata [27],\U_AHB/h2h_hwdata [2]}),
    .q({gpio_out_pad[27],gpio_out_pad[2]}));  // src/AHB.v(64)
  // src/AHB.v(64)
  // src/AHB.v(64)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTF1("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG0("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG1("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1101110011110000),
    .INIT_LUTF1(16'b1101110011110000),
    .INIT_LUTG0(16'b1101110011110000),
    .INIT_LUTG1(16'b1101110011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg17_b28|U_AHB/reg17_b31  (
    .a({\U_AHB/n38 ,\U_AHB/n38 }),
    .b({\U_AHB/n36 ,\U_AHB/n36 }),
    .c({gpio_out_pad[28],gpio_out_pad[31]}),
    .clk(clk100m),
    .d({\U_AHB/h2h_hwdata [28],\U_AHB/h2h_hwdata [31]}),
    .q({gpio_out_pad[28],gpio_out_pad[31]}));  // src/AHB.v(64)
  // src/OnePWM.v(48)
  // src/AHB.v(64)
  EF2_PHY_LSLICE #(
    //.LUTF0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTF1("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUTG0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUTG1("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000011001010),
    .INIT_LUTF1(16'b1101110011110000),
    .INIT_LUTG0(16'b1100000011001010),
    .INIT_LUTG1(16'b1101110011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg17_b30|PWM6/reg2_b27  (
    .a({\U_AHB/n38 ,\PWM6/pnumr [27]}),
    .b({\U_AHB/n36 ,pnum6[27]}),
    .c({gpio_out_pad[30],pnum6[32]}),
    .clk(clk100m),
    .d({\U_AHB/h2h_hwdata [30],pwm_start_stop[22]}),
    .q({gpio_out_pad[30],\PWM6/pnumr[27]_keep }));  // src/OnePWM.v(48)
  // src/AHB.v(67)
  // src/AHB.v(67)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b1010100000100000),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b1010100000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg18_b0|U_AHB/reg18_b28  (
    .a({\PWM0/n24 ,_al_u3312_o}),
    .b({\PWM0/n25_neg_lutinv ,\U_AHB/n102 }),
    .c({\PWM0/n26 [0],\U_AHB/n99 }),
    .clk(clk100m),
    .d({\PWM0/pnumr [0],pnumcnt6[11]}),
    .e({open_n28293,pnumcnt7[11]}),
    .mi({\U_AHB/h2h_hwdata [0],\U_AHB/h2h_hwdata [28]}),
    .sr(\U_AHB/n45 ),
    .f({_al_u1739_o,_al_u3313_o}),
    .q({pnum0[0],pnum0[28]}));  // src/AHB.v(67)
  // src/AHB.v(67)
  // src/AHB.v(67)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg18_b10|U_AHB/reg18_b32  (
    .a({\PWM0/n24 ,\PWM0/n24 }),
    .b({\PWM0/n25_neg_lutinv ,\PWM0/n25_neg_lutinv }),
    .c(\PWM0/n26 [10:9]),
    .clk(clk100m),
    .d(\PWM0/pnumr [10:9]),
    .mi({\U_AHB/h2h_hwdata [10],1'b1}),
    .sr(\U_AHB/n45 ),
    .f({_al_u1735_o,_al_u1693_o}),
    .q({pnum0[10],pnum0[32]}));  // src/AHB.v(67)
  // src/AHB.v(67)
  // src/AHB.v(67)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg18_b11|U_AHB/reg18_b8  (
    .a({\PWM0/n24 ,\PWM0/n24 }),
    .b({\PWM0/n25_neg_lutinv ,\PWM0/n25_neg_lutinv }),
    .c({\PWM0/n26 [11],\PWM0/n26 [8]}),
    .clk(clk100m),
    .d({\PWM0/pnumr [11],\PWM0/pnumr [8]}),
    .mi({\U_AHB/h2h_hwdata [11],\U_AHB/h2h_hwdata [8]}),
    .sr(\U_AHB/n45 ),
    .f({_al_u1733_o,_al_u1695_o}),
    .q({pnum0[11],pnum0[8]}));  // src/AHB.v(67)
  // src/AHB.v(67)
  // src/AHB.v(67)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg18_b12|U_AHB/reg18_b7  (
    .a({\PWM0/n24 ,\PWM0/n24 }),
    .b({\PWM0/n25_neg_lutinv ,\PWM0/n25_neg_lutinv }),
    .c({\PWM0/n26 [12],\PWM0/n26 [7]}),
    .clk(clk100m),
    .d({\PWM0/pnumr [12],\PWM0/pnumr [7]}),
    .mi({\U_AHB/h2h_hwdata [12],\U_AHB/h2h_hwdata [7]}),
    .sr(\U_AHB/n45 ),
    .f({_al_u1731_o,_al_u1697_o}),
    .q({pnum0[12],pnum0[7]}));  // src/AHB.v(67)
  // src/AHB.v(67)
  // src/AHB.v(67)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg18_b13|U_AHB/reg18_b6  (
    .a({\PWM0/n24 ,\PWM0/n24 }),
    .b({\PWM0/n25_neg_lutinv ,\PWM0/n25_neg_lutinv }),
    .c({\PWM0/n26 [13],\PWM0/n26 [6]}),
    .clk(clk100m),
    .d({\PWM0/pnumr [13],\PWM0/pnumr [6]}),
    .mi({\U_AHB/h2h_hwdata [13],\U_AHB/h2h_hwdata [6]}),
    .sr(\U_AHB/n45 ),
    .f({_al_u1729_o,_al_u1699_o}),
    .q({pnum0[13],pnum0[6]}));  // src/AHB.v(67)
  // src/AHB.v(67)
  // src/AHB.v(67)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg18_b14|U_AHB/reg18_b5  (
    .a({\PWM0/n24 ,\PWM0/n24 }),
    .b({\PWM0/n25_neg_lutinv ,\PWM0/n25_neg_lutinv }),
    .c({\PWM0/n26 [14],\PWM0/n26 [5]}),
    .clk(clk100m),
    .d({\PWM0/pnumr [14],\PWM0/pnumr [5]}),
    .mi({\U_AHB/h2h_hwdata [14],\U_AHB/h2h_hwdata [5]}),
    .sr(\U_AHB/n45 ),
    .f({_al_u1727_o,_al_u1701_o}),
    .q({pnum0[14],pnum0[5]}));  // src/AHB.v(67)
  // src/AHB.v(67)
  // src/AHB.v(67)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg18_b15|U_AHB/reg18_b4  (
    .a({\PWM0/n24 ,\PWM0/n24 }),
    .b({\PWM0/n25_neg_lutinv ,\PWM0/n25_neg_lutinv }),
    .c({\PWM0/n26 [15],\PWM0/n26 [4]}),
    .clk(clk100m),
    .d({\PWM0/pnumr [15],\PWM0/pnumr [4]}),
    .mi({\U_AHB/h2h_hwdata [15],\U_AHB/h2h_hwdata [4]}),
    .sr(\U_AHB/n45 ),
    .f({_al_u1725_o,_al_u1703_o}),
    .q({pnum0[15],pnum0[4]}));  // src/AHB.v(67)
  // src/AHB.v(67)
  // src/AHB.v(67)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg18_b16|U_AHB/reg18_b3  (
    .a({\PWM0/n24 ,\PWM0/n24 }),
    .b({\PWM0/n25_neg_lutinv ,\PWM0/n25_neg_lutinv }),
    .c({\PWM0/n26 [16],\PWM0/n26 [3]}),
    .clk(clk100m),
    .d({\PWM0/pnumr [16],\PWM0/pnumr [3]}),
    .mi({\U_AHB/h2h_hwdata [16],\U_AHB/h2h_hwdata [3]}),
    .sr(\U_AHB/n45 ),
    .f({_al_u1723_o,_al_u1705_o}),
    .q({pnum0[16],pnum0[3]}));  // src/AHB.v(67)
  // src/AHB.v(67)
  // src/AHB.v(67)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg18_b17|U_AHB/reg18_b23  (
    .a({\PWM0/n24 ,\PWM0/n24 }),
    .b({\PWM0/n25_neg_lutinv ,\PWM0/n25_neg_lutinv }),
    .c({\PWM0/n26 [17],\PWM0/n26 [23]}),
    .clk(clk100m),
    .d({\PWM0/pnumr [17],\PWM0/pnumr [23]}),
    .mi({\U_AHB/h2h_hwdata [17],\U_AHB/h2h_hwdata [23]}),
    .sr(\U_AHB/n45 ),
    .f({_al_u1721_o,_al_u1707_o}),
    .q({pnum0[17],pnum0[23]}));  // src/AHB.v(67)
  // src/AHB.v(67)
  // src/AHB.v(67)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg18_b18|U_AHB/reg18_b22  (
    .a({\PWM0/n24 ,\PWM0/n24 }),
    .b({\PWM0/n25_neg_lutinv ,\PWM0/n25_neg_lutinv }),
    .c({\PWM0/n26 [18],\PWM0/n26 [22]}),
    .clk(clk100m),
    .d({\PWM0/pnumr [18],\PWM0/pnumr [22]}),
    .mi({\U_AHB/h2h_hwdata [18],\U_AHB/h2h_hwdata [22]}),
    .sr(\U_AHB/n45 ),
    .f({_al_u1719_o,_al_u1709_o}),
    .q({pnum0[18],pnum0[22]}));  // src/AHB.v(67)
  // src/AHB.v(67)
  // src/AHB.v(67)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg18_b19|U_AHB/reg18_b21  (
    .a({\PWM0/n24 ,\PWM0/n24 }),
    .b({\PWM0/n25_neg_lutinv ,\PWM0/n25_neg_lutinv }),
    .c({\PWM0/n26 [19],\PWM0/n26 [21]}),
    .clk(clk100m),
    .d({\PWM0/pnumr [19],\PWM0/pnumr [21]}),
    .mi({\U_AHB/h2h_hwdata [19],\U_AHB/h2h_hwdata [21]}),
    .sr(\U_AHB/n45 ),
    .f({_al_u1717_o,_al_u1711_o}),
    .q({pnum0[19],pnum0[21]}));  // src/AHB.v(67)
  // src/AHB.v(67)
  // src/AHB.v(67)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg18_b1|U_AHB/reg18_b20  (
    .a({\PWM0/n24 ,\PWM0/n24 }),
    .b({\PWM0/n25_neg_lutinv ,\PWM0/n25_neg_lutinv }),
    .c({\PWM0/n26 [1],\PWM0/n26 [20]}),
    .clk(clk100m),
    .d({\PWM0/pnumr [1],\PWM0/pnumr [20]}),
    .mi({\U_AHB/h2h_hwdata [1],\U_AHB/h2h_hwdata [20]}),
    .sr(\U_AHB/n45 ),
    .f({_al_u1737_o,_al_u1713_o}),
    .q({pnum0[1],pnum0[20]}));  // src/AHB.v(67)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg18_b2  (
    .a({open_n28463,\PWM0/n24 }),
    .b({open_n28464,\PWM0/n25_neg_lutinv }),
    .c({open_n28465,\PWM0/n26 [2]}),
    .clk(clk100m),
    .d({open_n28467,\PWM0/pnumr [2]}),
    .mi({open_n28478,\U_AHB/h2h_hwdata [2]}),
    .sr(\U_AHB/n45 ),
    .f({open_n28479,_al_u1715_o}),
    .q({open_n28483,pnum0[2]}));  // src/AHB.v(67)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg18_b24  (
    .a({open_n28484,_al_u3174_o}),
    .b({open_n28485,\U_AHB/n96 }),
    .c({open_n28486,\U_AHB/n93 }),
    .clk(clk100m),
    .d({open_n28488,pnumcntF[23]}),
    .e({open_n28489,pwm_state_read[7]}),
    .mi({open_n28491,\U_AHB/h2h_hwdata [24]}),
    .sr(\U_AHB/n45 ),
    .f({open_n28503,_al_u3175_o}),
    .q({open_n28507,pnum0[24]}));  // src/AHB.v(67)
  // src/AHB.v(67)
  // src/AHB.v(67)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg18_b26|U_AHB/reg18_b9  (
    .a({_al_u3334_o,_al_u3268_o}),
    .b({\U_AHB/n102 ,\U_AHB/n102 }),
    .c({\U_AHB/n99 ,\U_AHB/n99 }),
    .clk(clk100m),
    .d({pnumcnt6[1],pnumcnt6[15]}),
    .e({pnumcnt7[1],pnumcnt7[15]}),
    .mi({\U_AHB/h2h_hwdata [26],\U_AHB/h2h_hwdata [9]}),
    .sr(\U_AHB/n45 ),
    .f({_al_u3335_o,_al_u3269_o}),
    .q({pnum0[26],pnum0[9]}));  // src/AHB.v(67)
  // src/AHB.v(67)
  // src/AHB.v(67)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg18_b27|U_AHB/reg18_b31  (
    .a({_al_u3323_o,_al_u3279_o}),
    .b({\U_AHB/n102 ,\U_AHB/n102 }),
    .c({\U_AHB/n99 ,\U_AHB/n99 }),
    .clk(clk100m),
    .d({pnumcnt6[10],pnumcnt6[14]}),
    .e({pnumcnt7[10],pnumcnt7[14]}),
    .mi({\U_AHB/h2h_hwdata [27],\U_AHB/h2h_hwdata [31]}),
    .sr(\U_AHB/n45 ),
    .f({_al_u3324_o,_al_u3280_o}),
    .q({pnum0[27],pnum0[31]}));  // src/AHB.v(67)
  // src/AHB.v(68)
  // src/AHB.v(68)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b1010100000100000),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b1010100000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg19_b0|U_AHB/reg19_b28  (
    .a({\PWM1/n24 ,_al_u3213_o}),
    .b({\PWM1/n25_neg_lutinv ,\U_AHB/n102 }),
    .c({\PWM1/n26 [0],\U_AHB/n99 }),
    .clk(clk100m),
    .d({\PWM1/pnumr [0],pnumcnt6[2]}),
    .e({open_n28541,pnumcnt7[2]}),
    .mi({\U_AHB/h2h_hwdata [0],\U_AHB/h2h_hwdata [28]}),
    .sr(\U_AHB/n47 ),
    .f({_al_u1821_o,_al_u3214_o}),
    .q({pnum1[0],pnum1[28]}));  // src/AHB.v(68)
  // src/AHB.v(68)
  // src/AHB.v(68)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg19_b10|U_AHB/reg19_b32  (
    .a({\PWM1/n24 ,\PWM1/n24 }),
    .b({\PWM1/n25_neg_lutinv ,\PWM1/n25_neg_lutinv }),
    .c(\PWM1/n26 [10:9]),
    .clk(clk100m),
    .d(\PWM1/pnumr [10:9]),
    .mi({\U_AHB/h2h_hwdata [10],1'b1}),
    .sr(\U_AHB/n47 ),
    .f({_al_u1817_o,_al_u1775_o}),
    .q({pnum1[10],pnum1[32]}));  // src/AHB.v(68)
  // src/AHB.v(68)
  // src/AHB.v(68)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg19_b11|U_AHB/reg19_b8  (
    .a({\PWM1/n24 ,\PWM1/n24 }),
    .b({\PWM1/n25_neg_lutinv ,\PWM1/n25_neg_lutinv }),
    .c({\PWM1/n26 [11],\PWM1/n26 [8]}),
    .clk(clk100m),
    .d({\PWM1/pnumr [11],\PWM1/pnumr [8]}),
    .mi({\U_AHB/h2h_hwdata [11],\U_AHB/h2h_hwdata [8]}),
    .sr(\U_AHB/n47 ),
    .f({_al_u1815_o,_al_u1777_o}),
    .q({pnum1[11],pnum1[8]}));  // src/AHB.v(68)
  // src/AHB.v(68)
  // src/AHB.v(68)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg19_b12|U_AHB/reg19_b7  (
    .a({\PWM1/n24 ,\PWM1/n24 }),
    .b({\PWM1/n25_neg_lutinv ,\PWM1/n25_neg_lutinv }),
    .c({\PWM1/n26 [12],\PWM1/n26 [7]}),
    .clk(clk100m),
    .d({\PWM1/pnumr [12],\PWM1/pnumr [7]}),
    .mi({\U_AHB/h2h_hwdata [12],\U_AHB/h2h_hwdata [7]}),
    .sr(\U_AHB/n47 ),
    .f({_al_u1813_o,_al_u1779_o}),
    .q({pnum1[12],pnum1[7]}));  // src/AHB.v(68)
  // src/AHB.v(68)
  // src/AHB.v(68)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg19_b13|U_AHB/reg19_b6  (
    .a({\PWM1/n24 ,\PWM1/n24 }),
    .b({\PWM1/n25_neg_lutinv ,\PWM1/n25_neg_lutinv }),
    .c({\PWM1/n26 [13],\PWM1/n26 [6]}),
    .clk(clk100m),
    .d({\PWM1/pnumr [13],\PWM1/pnumr [6]}),
    .mi({\U_AHB/h2h_hwdata [13],\U_AHB/h2h_hwdata [6]}),
    .sr(\U_AHB/n47 ),
    .f({_al_u1811_o,_al_u1781_o}),
    .q({pnum1[13],pnum1[6]}));  // src/AHB.v(68)
  // src/AHB.v(68)
  // src/AHB.v(68)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg19_b14|U_AHB/reg19_b5  (
    .a({\PWM1/n24 ,\PWM1/n24 }),
    .b({\PWM1/n25_neg_lutinv ,\PWM1/n25_neg_lutinv }),
    .c({\PWM1/n26 [14],\PWM1/n26 [5]}),
    .clk(clk100m),
    .d({\PWM1/pnumr [14],\PWM1/pnumr [5]}),
    .mi({\U_AHB/h2h_hwdata [14],\U_AHB/h2h_hwdata [5]}),
    .sr(\U_AHB/n47 ),
    .f({_al_u1809_o,_al_u1783_o}),
    .q({pnum1[14],pnum1[5]}));  // src/AHB.v(68)
  // src/AHB.v(68)
  // src/AHB.v(68)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg19_b15|U_AHB/reg19_b4  (
    .a({\PWM1/n24 ,\PWM1/n24 }),
    .b({\PWM1/n25_neg_lutinv ,\PWM1/n25_neg_lutinv }),
    .c({\PWM1/n26 [15],\PWM1/n26 [4]}),
    .clk(clk100m),
    .d({\PWM1/pnumr [15],\PWM1/pnumr [4]}),
    .mi({\U_AHB/h2h_hwdata [15],\U_AHB/h2h_hwdata [4]}),
    .sr(\U_AHB/n47 ),
    .f({_al_u1807_o,_al_u1785_o}),
    .q({pnum1[15],pnum1[4]}));  // src/AHB.v(68)
  // src/AHB.v(68)
  // src/AHB.v(68)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg19_b16|U_AHB/reg19_b3  (
    .a({\PWM1/n24 ,\PWM1/n24 }),
    .b({\PWM1/n25_neg_lutinv ,\PWM1/n25_neg_lutinv }),
    .c({\PWM1/n26 [16],\PWM1/n26 [3]}),
    .clk(clk100m),
    .d({\PWM1/pnumr [16],\PWM1/pnumr [3]}),
    .mi({\U_AHB/h2h_hwdata [16],\U_AHB/h2h_hwdata [3]}),
    .sr(\U_AHB/n47 ),
    .f({_al_u1805_o,_al_u1787_o}),
    .q({pnum1[16],pnum1[3]}));  // src/AHB.v(68)
  // src/AHB.v(68)
  // src/AHB.v(68)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg19_b17|U_AHB/reg19_b23  (
    .a({\PWM1/n24 ,\PWM1/n24 }),
    .b({\PWM1/n25_neg_lutinv ,\PWM1/n25_neg_lutinv }),
    .c({\PWM1/n26 [17],\PWM1/n26 [23]}),
    .clk(clk100m),
    .d({\PWM1/pnumr [17],\PWM1/pnumr [23]}),
    .mi({\U_AHB/h2h_hwdata [17],\U_AHB/h2h_hwdata [23]}),
    .sr(\U_AHB/n47 ),
    .f({_al_u1803_o,_al_u1789_o}),
    .q({pnum1[17],pnum1[23]}));  // src/AHB.v(68)
  // src/AHB.v(68)
  // src/AHB.v(68)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg19_b18|U_AHB/reg19_b22  (
    .a({\PWM1/n24 ,\PWM1/n24 }),
    .b({\PWM1/n25_neg_lutinv ,\PWM1/n25_neg_lutinv }),
    .c({\PWM1/n26 [18],\PWM1/n26 [22]}),
    .clk(clk100m),
    .d({\PWM1/pnumr [18],\PWM1/pnumr [22]}),
    .mi({\U_AHB/h2h_hwdata [18],\U_AHB/h2h_hwdata [22]}),
    .sr(\U_AHB/n47 ),
    .f({_al_u1801_o,_al_u1791_o}),
    .q({pnum1[18],pnum1[22]}));  // src/AHB.v(68)
  // src/AHB.v(68)
  // src/AHB.v(68)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg19_b19|U_AHB/reg19_b21  (
    .a({\PWM1/n24 ,\PWM1/n24 }),
    .b({\PWM1/n25_neg_lutinv ,\PWM1/n25_neg_lutinv }),
    .c({\PWM1/n26 [19],\PWM1/n26 [21]}),
    .clk(clk100m),
    .d({\PWM1/pnumr [19],\PWM1/pnumr [21]}),
    .mi({\U_AHB/h2h_hwdata [19],\U_AHB/h2h_hwdata [21]}),
    .sr(\U_AHB/n47 ),
    .f({_al_u1799_o,_al_u1793_o}),
    .q({pnum1[19],pnum1[21]}));  // src/AHB.v(68)
  // src/AHB.v(68)
  // src/AHB.v(68)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg19_b1|U_AHB/reg19_b20  (
    .a({\PWM1/n24 ,\PWM1/n24 }),
    .b({\PWM1/n25_neg_lutinv ,\PWM1/n25_neg_lutinv }),
    .c({\PWM1/n26 [1],\PWM1/n26 [20]}),
    .clk(clk100m),
    .d({\PWM1/pnumr [1],\PWM1/pnumr [20]}),
    .mi({\U_AHB/h2h_hwdata [1],\U_AHB/h2h_hwdata [20]}),
    .sr(\U_AHB/n47 ),
    .f({_al_u1819_o,_al_u1795_o}),
    .q({pnum1[1],pnum1[20]}));  // src/AHB.v(68)
  // src/AHB.v(68)
  // src/AHB.v(68)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg19_b27|U_AHB/reg19_b30  (
    .a({_al_u3224_o,_al_u3191_o}),
    .b({\U_AHB/n102 ,\U_AHB/n102 }),
    .c({\U_AHB/n99 ,\U_AHB/n99 }),
    .clk(clk100m),
    .d({pnumcnt6[19],pnumcnt6[21]}),
    .e({pnumcnt7[19],pnumcnt7[21]}),
    .mi({\U_AHB/h2h_hwdata [27],\U_AHB/h2h_hwdata [30]}),
    .sr(\U_AHB/n47 ),
    .f({_al_u3225_o,_al_u3192_o}),
    .q({pnum1[27],pnum1[30]}));  // src/AHB.v(68)
  // src/AHB.v(46)
  // src/AHB.v(46)
  EF2_PHY_MSLICE #(
    //.LUT0("(D*~C*B*A)"),
    //.LUT1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100000000000),
    .INIT_LUT1(16'b1000010000100001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg1_b10|U_AHB/reg1_b0  (
    .a({\PWM0/FreCnt [10],\U_AHB/h2h_hwrite }),
    .b({\PWM0/FreCnt [2],\U_AHB/h2h_haddr [13]}),
    .c({\PWM0/FreCntr [10],\U_AHB/h2h_haddr [14]}),
    .ce(\U_AHB/n2 ),
    .clk(clk100m),
    .d({\PWM0/FreCntr [2],\U_AHB/h2h_haddr [5]}),
    .mi({\U_AHB/h2h_hwdata [10],\U_AHB/h2h_hwdata [0]}),
    .f({_al_u1367_o,\U_AHB/n2 }),
    .q({freq0[10],freq0[0]}));  // src/AHB.v(46)
  // src/AHB.v(46)
  // src/AHB.v(46)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg1_b11|U_AHB/reg1_b22  (
    .a({open_n28741,_al_u739_o}),
    .b({_al_u738_o,\PWM0/FreCnt [2]}),
    .c({_al_u740_o,\PWM0/FreCnt [20]}),
    .ce(\U_AHB/n2 ),
    .clk(clk100m),
    .d({_al_u736_o,\PWM0/FreCnt [21]}),
    .e({open_n28742,\PWM0/FreCnt [22]}),
    .mi({\U_AHB/h2h_hwdata [11],\U_AHB/h2h_hwdata [22]}),
    .f({\PWM0/n0_lutinv ,_al_u740_o}),
    .q({freq0[11],freq0[22]}));  // src/AHB.v(46)
  // src/AHB.v(46)
  // src/AHB.v(46)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~(D*~B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1000110010101111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg1_b15|U_AHB/reg1_b17  (
    .a({\PWM0/FreCnt [12],open_n28759}),
    .b({\PWM0/FreCnt [15],open_n28760}),
    .c({\PWM0/FreCntr [12],pwm_state_read[0]}),
    .ce(\U_AHB/n2 ),
    .clk(clk100m),
    .d({\PWM0/FreCntr [15],\PWM0/n0_lutinv }),
    .mi({\U_AHB/h2h_hwdata [15],\U_AHB/h2h_hwdata [17]}),
    .f({_al_u1366_o,\PWM0/n24 }),
    .q({freq0[15],freq0[17]}));  // src/AHB.v(46)
  // src/AHB.v(46)
  // src/AHB.v(46)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*~C)*~(D*~B))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(A*~(1*~C)*~(D*~B))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000100010101010),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000000010100000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg1_b16|U_AHB/reg1_b14  (
    .a({\PWM0/FreCnt [16],_al_u1745_o}),
    .b({\PWM0/FreCnt [26],\PWM0/FreCnt [13]}),
    .c({\PWM0/FreCntr [16],\PWM0/FreCnt [25]}),
    .ce(\U_AHB/n2 ),
    .clk(clk100m),
    .d({\PWM0/FreCntr [26],\PWM0/FreCntr [14]}),
    .e({open_n28775,\PWM0/FreCntr [26]}),
    .mi({\U_AHB/h2h_hwdata [16],\U_AHB/h2h_hwdata [14]}),
    .f({_al_u1375_o,_al_u1746_o}),
    .q({freq0[16],freq0[14]}));  // src/AHB.v(46)
  // src/AHB.v(46)
  // src/AHB.v(46)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*~C)*~(D*~B))"),
    //.LUTF1("(A*~(0@C)*~(D@B))"),
    //.LUTG0("(A*~(1*~C)*~(D*~B))"),
    //.LUTG1("(A*~(1@C)*~(D@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000100010101010),
    .INIT_LUTF1(16'b0000100000000010),
    .INIT_LUTG0(16'b1000000010100000),
    .INIT_LUTG1(16'b1000000000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg1_b19|U_AHB/reg1_b13  (
    .a({_al_u1375_o,_al_u1741_o}),
    .b(\PWM0/FreCnt [13:12]),
    .c({\PWM0/FreCnt [19],\PWM0/FreCnt [5]}),
    .ce(\U_AHB/n2 ),
    .clk(clk100m),
    .d({\PWM0/FreCntr [13],\PWM0/FreCntr [13]}),
    .e({\PWM0/FreCntr [19],\PWM0/FreCntr [6]}),
    .mi({\U_AHB/h2h_hwdata [19],\U_AHB/h2h_hwdata [13]}),
    .f({_al_u1376_o,_al_u1742_o}),
    .q({freq0[19],freq0[13]}));  // src/AHB.v(46)
  // src/AHB.v(46)
  // src/AHB.v(46)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(~(~D*B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b1111010100110001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg1_b1|U_AHB/reg1_b18  (
    .a({\PWM0/FreCnt [1],open_n28808}),
    .b({\PWM0/FreCnt [15],limit_r_pad[0]}),
    .c({\PWM0/FreCntr [1],limit_l_pad[0]}),
    .ce(\U_AHB/n2 ),
    .clk(clk100m),
    .d({\PWM0/FreCntr [15],\PWM0/n11 }),
    .mi({\U_AHB/h2h_hwdata [1],\U_AHB/h2h_hwdata [18]}),
    .f({_al_u1371_o,_al_u3008_o}),
    .q({freq0[1],freq0[18]}));  // src/AHB.v(46)
  // src/AHB.v(46)
  // src/AHB.v(46)
  EF2_PHY_MSLICE #(
    //.LUT0("(~D*~C*~B*A)"),
    //.LUT1("(B*A*~(D@C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000010),
    .INIT_LUT1(16'b1000000000001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg1_b21|U_AHB/reg1_b7  (
    .a({_al_u1366_o,_al_u735_o}),
    .b({_al_u1367_o,\PWM0/FreCnt [7]}),
    .c({\PWM0/FreCnt [21],\PWM0/FreCnt [8]}),
    .ce(\U_AHB/n2 ),
    .clk(clk100m),
    .d({\PWM0/FreCntr [21],\PWM0/FreCnt [9]}),
    .mi({\U_AHB/h2h_hwdata [21],\U_AHB/h2h_hwdata [7]}),
    .f({_al_u1368_o,_al_u736_o}),
    .q({freq0[21],freq0[7]}));  // src/AHB.v(46)
  // src/AHB.v(46)
  // src/AHB.v(46)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg1_b23|U_AHB/reg1_b3  (
    .a({\PWM0/FreCnt [23],_al_u734_o}),
    .b({\PWM0/FreCnt [24],\PWM0/FreCnt [3]}),
    .c({\PWM0/FreCnt [25],\PWM0/FreCnt [4]}),
    .ce(\U_AHB/n2 ),
    .clk(clk100m),
    .d({\PWM0/FreCnt [26],\PWM0/FreCnt [5]}),
    .e({open_n28837,\PWM0/FreCnt [6]}),
    .mi({\U_AHB/h2h_hwdata [23],\U_AHB/h2h_hwdata [3]}),
    .f({_al_u734_o,_al_u735_o}),
    .q({freq0[23],freq0[3]}));  // src/AHB.v(46)
  // src/AHB.v(46)
  // src/AHB.v(46)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg1_b24|U_AHB/reg1_b9  (
    .a({_al_u3333_o,_al_u3306_o}),
    .b({\U_AHB/n96 ,\U_AHB/n96 }),
    .c({\U_AHB/n93 ,\U_AHB/n93 }),
    .ce(\U_AHB/n2 ),
    .clk(clk100m),
    .d({pnumcnt4[1],pnumcntF[12]}),
    .e({pnumcnt5[1],pwm_state_read[12]}),
    .mi({\U_AHB/h2h_hwdata [24],\U_AHB/h2h_hwdata [9]}),
    .f({_al_u3334_o,_al_u3307_o}),
    .q({freq0[24],freq0[9]}));  // src/AHB.v(46)
  // src/AHB.v(46)
  // src/AHB.v(46)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg1_b25|U_AHB/reg1_b5  (
    .a({_al_u3328_o,_al_u3317_o}),
    .b({\U_AHB/n96 ,\U_AHB/n96 }),
    .c({\U_AHB/n93 ,\U_AHB/n93 }),
    .ce(\U_AHB/n2 ),
    .clk(clk100m),
    .d({pnumcntF[10],pnumcntF[11]}),
    .e({pwm_state_read[10],pwm_state_read[11]}),
    .mi({\U_AHB/h2h_hwdata [25],\U_AHB/h2h_hwdata [5]}),
    .f({_al_u3329_o,_al_u3318_o}),
    .q({freq0[25],freq0[5]}));  // src/AHB.v(46)
  // src/AHB.v(46)
  // src/AHB.v(46)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg1_b6|U_AHB/reg1_b4  (
    .a({\PWM0/FreCnt [6],_al_u1362_o}),
    .b({\PWM0/FreCnt [7],\PWM0/FreCnt [4]}),
    .c({\PWM0/FreCntr [6],\PWM0/FreCnt [9]}),
    .ce(\U_AHB/n2 ),
    .clk(clk100m),
    .d({\PWM0/FreCntr [7],\PWM0/FreCntr [4]}),
    .e({open_n28886,\PWM0/FreCntr [9]}),
    .mi({\U_AHB/h2h_hwdata [6],\U_AHB/h2h_hwdata [4]}),
    .f({_al_u1362_o,_al_u1363_o}),
    .q({freq0[6],freq0[4]}));  // src/AHB.v(46)
  // src/AHB.v(69)
  // src/AHB.v(69)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(D*~C*B*A)"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(D*~C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000100000000000),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000100000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg20_b0|U_AHB/reg20_b28  (
    .a({\U_AHB/h2h_hwrite ,_al_u3113_o}),
    .b({\U_AHB/h2h_haddr [2],\U_AHB/n102 }),
    .c({\U_AHB/h2h_haddr [13],\U_AHB/n99 }),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [14],pnumcnt6[7]}),
    .e({open_n28904,pnumcnt7[7]}),
    .mi({\U_AHB/h2h_hwdata [0],\U_AHB/h2h_hwdata [28]}),
    .sr(\U_AHB/n51 ),
    .f({\U_AHB/n51 ,_al_u3114_o}),
    .q({pnum2[0],pnum2[28]}));  // src/AHB.v(69)
  // src/AHB.v(69)
  // src/AHB.v(69)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b1010100000100000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1010100000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg20_b10|U_AHB/reg20_b9  (
    .a({\PWM2/n24 ,_al_u2500_o}),
    .b({\PWM2/n25_neg_lutinv ,pnumcntA[21]}),
    .c({\PWM2/n26 [10],pnumcntA[22]}),
    .clk(clk100m),
    .d({\PWM2/pnumr [10],pnumcntA[23]}),
    .e({open_n28921,pnumcntA[2]}),
    .mi(\U_AHB/h2h_hwdata [10:9]),
    .sr(\U_AHB/n51 ),
    .f({_al_u1899_o,_al_u2501_o}),
    .q(pnum2[10:9]));  // src/AHB.v(69)
  // src/AHB.v(69)
  // src/AHB.v(69)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg20_b11|U_AHB/reg20_b32  (
    .a({\PWM2/n24 ,\PWM2/n24 }),
    .b({\PWM2/n25_neg_lutinv ,\PWM2/n25_neg_lutinv }),
    .c({\PWM2/n26 [11],\PWM2/n26 [9]}),
    .clk(clk100m),
    .d({\PWM2/pnumr [11],\PWM2/pnumr [9]}),
    .mi({\U_AHB/h2h_hwdata [11],1'b1}),
    .sr(\U_AHB/n51 ),
    .f({_al_u1897_o,_al_u1857_o}),
    .q({pnum2[11],pnum2[32]}));  // src/AHB.v(69)
  // src/AHB.v(69)
  // src/AHB.v(69)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg20_b12|U_AHB/reg20_b8  (
    .a({\PWM2/n24 ,\PWM2/n24 }),
    .b({\PWM2/n25_neg_lutinv ,\PWM2/n25_neg_lutinv }),
    .c({\PWM2/n26 [12],\PWM2/n26 [8]}),
    .clk(clk100m),
    .d({\PWM2/pnumr [12],\PWM2/pnumr [8]}),
    .mi({\U_AHB/h2h_hwdata [12],\U_AHB/h2h_hwdata [8]}),
    .sr(\U_AHB/n51 ),
    .f({_al_u1895_o,_al_u1859_o}),
    .q({pnum2[12],pnum2[8]}));  // src/AHB.v(69)
  // src/AHB.v(69)
  // src/AHB.v(69)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg20_b13|U_AHB/reg20_b7  (
    .a({\PWM2/n24 ,\PWM2/n24 }),
    .b({\PWM2/n25_neg_lutinv ,\PWM2/n25_neg_lutinv }),
    .c({\PWM2/n26 [13],\PWM2/n26 [7]}),
    .clk(clk100m),
    .d({\PWM2/pnumr [13],\PWM2/pnumr [7]}),
    .mi({\U_AHB/h2h_hwdata [13],\U_AHB/h2h_hwdata [7]}),
    .sr(\U_AHB/n51 ),
    .f({_al_u1893_o,_al_u1861_o}),
    .q({pnum2[13],pnum2[7]}));  // src/AHB.v(69)
  // src/AHB.v(69)
  // src/AHB.v(69)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg20_b14|U_AHB/reg20_b6  (
    .a({\PWM2/n24 ,\PWM2/n24 }),
    .b({\PWM2/n25_neg_lutinv ,\PWM2/n25_neg_lutinv }),
    .c({\PWM2/n26 [14],\PWM2/n26 [6]}),
    .clk(clk100m),
    .d({\PWM2/pnumr [14],\PWM2/pnumr [6]}),
    .mi({\U_AHB/h2h_hwdata [14],\U_AHB/h2h_hwdata [6]}),
    .sr(\U_AHB/n51 ),
    .f({_al_u1891_o,_al_u1863_o}),
    .q({pnum2[14],pnum2[6]}));  // src/AHB.v(69)
  // src/AHB.v(69)
  // src/AHB.v(69)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg20_b15|U_AHB/reg20_b5  (
    .a({\PWM2/n24 ,\PWM2/n24 }),
    .b({\PWM2/n25_neg_lutinv ,\PWM2/n25_neg_lutinv }),
    .c({\PWM2/n26 [15],\PWM2/n26 [5]}),
    .clk(clk100m),
    .d({\PWM2/pnumr [15],\PWM2/pnumr [5]}),
    .mi({\U_AHB/h2h_hwdata [15],\U_AHB/h2h_hwdata [5]}),
    .sr(\U_AHB/n51 ),
    .f({_al_u1889_o,_al_u1865_o}),
    .q({pnum2[15],pnum2[5]}));  // src/AHB.v(69)
  // src/AHB.v(69)
  // src/AHB.v(69)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg20_b16|U_AHB/reg20_b4  (
    .a({\PWM2/n24 ,\PWM2/n24 }),
    .b({\PWM2/n25_neg_lutinv ,\PWM2/n25_neg_lutinv }),
    .c({\PWM2/n26 [16],\PWM2/n26 [4]}),
    .clk(clk100m),
    .d({\PWM2/pnumr [16],\PWM2/pnumr [4]}),
    .mi({\U_AHB/h2h_hwdata [16],\U_AHB/h2h_hwdata [4]}),
    .sr(\U_AHB/n51 ),
    .f({_al_u1887_o,_al_u1867_o}),
    .q({pnum2[16],pnum2[4]}));  // src/AHB.v(69)
  // src/AHB.v(69)
  // src/AHB.v(69)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg20_b17|U_AHB/reg20_b3  (
    .a({\PWM2/n24 ,\PWM2/n24 }),
    .b({\PWM2/n25_neg_lutinv ,\PWM2/n25_neg_lutinv }),
    .c({\PWM2/n26 [17],\PWM2/n26 [3]}),
    .clk(clk100m),
    .d({\PWM2/pnumr [17],\PWM2/pnumr [3]}),
    .mi({\U_AHB/h2h_hwdata [17],\U_AHB/h2h_hwdata [3]}),
    .sr(\U_AHB/n51 ),
    .f({_al_u1885_o,_al_u1869_o}),
    .q({pnum2[17],pnum2[3]}));  // src/AHB.v(69)
  // src/AHB.v(69)
  // src/AHB.v(69)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg20_b18|U_AHB/reg20_b23  (
    .a({\PWM2/n24 ,\PWM2/n24 }),
    .b({\PWM2/n25_neg_lutinv ,\PWM2/n25_neg_lutinv }),
    .c({\PWM2/n26 [18],\PWM2/n26 [23]}),
    .clk(clk100m),
    .d({\PWM2/pnumr [18],\PWM2/pnumr [23]}),
    .mi({\U_AHB/h2h_hwdata [18],\U_AHB/h2h_hwdata [23]}),
    .sr(\U_AHB/n51 ),
    .f({_al_u1883_o,_al_u1871_o}),
    .q({pnum2[18],pnum2[23]}));  // src/AHB.v(69)
  // src/AHB.v(69)
  // src/AHB.v(69)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg20_b19|U_AHB/reg20_b22  (
    .a({\PWM2/n24 ,\PWM2/n24 }),
    .b({\PWM2/n25_neg_lutinv ,\PWM2/n25_neg_lutinv }),
    .c({\PWM2/n26 [19],\PWM2/n26 [22]}),
    .clk(clk100m),
    .d({\PWM2/pnumr [19],\PWM2/pnumr [22]}),
    .mi({\U_AHB/h2h_hwdata [19],\U_AHB/h2h_hwdata [22]}),
    .sr(\U_AHB/n51 ),
    .f({_al_u1881_o,_al_u1873_o}),
    .q({pnum2[19],pnum2[22]}));  // src/AHB.v(69)
  // src/AHB.v(69)
  // src/AHB.v(69)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg20_b1|U_AHB/reg20_b21  (
    .a({\PWM2/n24 ,\PWM2/n24 }),
    .b({\PWM2/n25_neg_lutinv ,\PWM2/n25_neg_lutinv }),
    .c({\PWM2/n26 [1],\PWM2/n26 [21]}),
    .clk(clk100m),
    .d({\PWM2/pnumr [1],\PWM2/pnumr [21]}),
    .mi({\U_AHB/h2h_hwdata [1],\U_AHB/h2h_hwdata [21]}),
    .sr(\U_AHB/n51 ),
    .f({_al_u1901_o,_al_u1875_o}),
    .q({pnum2[1],pnum2[21]}));  // src/AHB.v(69)
  // src/AHB.v(69)
  // src/AHB.v(69)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg20_b27|U_AHB/reg20_b24  (
    .a({_al_u3124_o,_al_u3158_o}),
    .b({\U_AHB/n102 ,\U_AHB/n102 }),
    .c({\U_AHB/n99 ,\U_AHB/n99 }),
    .clk(clk100m),
    .d({pnumcnt6[6],pnumcnt6[3]}),
    .e({pnumcnt7[6],pnumcnt7[3]}),
    .mi({\U_AHB/h2h_hwdata [27],\U_AHB/h2h_hwdata [24]}),
    .sr(\U_AHB/n51 ),
    .f({_al_u3125_o,_al_u3159_o}),
    .q({pnum2[27],pnum2[24]}));  // src/AHB.v(69)
  // src/AHB.v(69)
  // src/AHB.v(69)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg20_b2|U_AHB/reg20_b20  (
    .a({\PWM2/n24 ,\PWM2/n24 }),
    .b({\PWM2/n25_neg_lutinv ,\PWM2/n25_neg_lutinv }),
    .c({\PWM2/n26 [2],\PWM2/n26 [20]}),
    .clk(clk100m),
    .d({\PWM2/pnumr [2],\PWM2/pnumr [20]}),
    .mi({\U_AHB/h2h_hwdata [2],\U_AHB/h2h_hwdata [20]}),
    .sr(\U_AHB/n51 ),
    .f({_al_u1879_o,_al_u1877_o}),
    .q({pnum2[2],pnum2[20]}));  // src/AHB.v(69)
  // src/AHB.v(70)
  // src/AHB.v(70)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg21_b10|U_AHB/reg21_b32  (
    .a({\PWM3/n24 ,\PWM3/n24 }),
    .b({\PWM3/n25_neg_lutinv ,\PWM3/n25_neg_lutinv }),
    .c(\PWM3/n26 [10:9]),
    .clk(clk100m),
    .d(\PWM3/pnumr [10:9]),
    .mi({\U_AHB/h2h_hwdata [10],1'b1}),
    .sr(\U_AHB/n53 ),
    .f({_al_u1979_o,_al_u1937_o}),
    .q({pnum3[10],pnum3[32]}));  // src/AHB.v(70)
  // src/AHB.v(70)
  // src/AHB.v(70)
  EF2_PHY_MSLICE #(
    //.LUT0("(D*~C*B*A)"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100000000000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg21_b11|U_AHB/reg21_b0  (
    .a({\PWM3/n24 ,\U_AHB/h2h_hwrite }),
    .b({\PWM3/n25_neg_lutinv ,\U_AHB/h2h_haddr [3]}),
    .c({\PWM3/n26 [11],\U_AHB/h2h_haddr [13]}),
    .clk(clk100m),
    .d({\PWM3/pnumr [11],\U_AHB/h2h_haddr [14]}),
    .mi({\U_AHB/h2h_hwdata [11],\U_AHB/h2h_hwdata [0]}),
    .sr(\U_AHB/n53 ),
    .f({_al_u1977_o,\U_AHB/n53 }),
    .q({pnum3[11],pnum3[0]}));  // src/AHB.v(70)
  // src/AHB.v(70)
  // src/AHB.v(70)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg21_b12|U_AHB/reg21_b8  (
    .a({\PWM3/n24 ,\PWM3/n24 }),
    .b({\PWM3/n25_neg_lutinv ,\PWM3/n25_neg_lutinv }),
    .c({\PWM3/n26 [12],\PWM3/n26 [8]}),
    .clk(clk100m),
    .d({\PWM3/pnumr [12],\PWM3/pnumr [8]}),
    .mi({\U_AHB/h2h_hwdata [12],\U_AHB/h2h_hwdata [8]}),
    .sr(\U_AHB/n53 ),
    .f({_al_u1975_o,_al_u1939_o}),
    .q({pnum3[12],pnum3[8]}));  // src/AHB.v(70)
  // src/AHB.v(70)
  // src/AHB.v(70)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg21_b13|U_AHB/reg21_b7  (
    .a({\PWM3/n24 ,\PWM3/n24 }),
    .b({\PWM3/n25_neg_lutinv ,\PWM3/n25_neg_lutinv }),
    .c({\PWM3/n26 [13],\PWM3/n26 [7]}),
    .clk(clk100m),
    .d({\PWM3/pnumr [13],\PWM3/pnumr [7]}),
    .mi({\U_AHB/h2h_hwdata [13],\U_AHB/h2h_hwdata [7]}),
    .sr(\U_AHB/n53 ),
    .f({_al_u1973_o,_al_u1941_o}),
    .q({pnum3[13],pnum3[7]}));  // src/AHB.v(70)
  // src/AHB.v(70)
  // src/AHB.v(70)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg21_b14|U_AHB/reg21_b6  (
    .a({\PWM3/n24 ,\PWM3/n24 }),
    .b({\PWM3/n25_neg_lutinv ,\PWM3/n25_neg_lutinv }),
    .c({\PWM3/n26 [14],\PWM3/n26 [6]}),
    .clk(clk100m),
    .d({\PWM3/pnumr [14],\PWM3/pnumr [6]}),
    .mi({\U_AHB/h2h_hwdata [14],\U_AHB/h2h_hwdata [6]}),
    .sr(\U_AHB/n53 ),
    .f({_al_u1971_o,_al_u1943_o}),
    .q({pnum3[14],pnum3[6]}));  // src/AHB.v(70)
  // src/AHB.v(70)
  // src/AHB.v(70)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg21_b15|U_AHB/reg21_b5  (
    .a({\PWM3/n24 ,\PWM3/n24 }),
    .b({\PWM3/n25_neg_lutinv ,\PWM3/n25_neg_lutinv }),
    .c({\PWM3/n26 [15],\PWM3/n26 [5]}),
    .clk(clk100m),
    .d({\PWM3/pnumr [15],\PWM3/pnumr [5]}),
    .mi({\U_AHB/h2h_hwdata [15],\U_AHB/h2h_hwdata [5]}),
    .sr(\U_AHB/n53 ),
    .f({_al_u1969_o,_al_u1945_o}),
    .q({pnum3[15],pnum3[5]}));  // src/AHB.v(70)
  // src/AHB.v(70)
  // src/AHB.v(70)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg21_b16|U_AHB/reg21_b4  (
    .a({\PWM3/n24 ,\PWM3/n24 }),
    .b({\PWM3/n25_neg_lutinv ,\PWM3/n25_neg_lutinv }),
    .c({\PWM3/n26 [16],\PWM3/n26 [4]}),
    .clk(clk100m),
    .d({\PWM3/pnumr [16],\PWM3/pnumr [4]}),
    .mi({\U_AHB/h2h_hwdata [16],\U_AHB/h2h_hwdata [4]}),
    .sr(\U_AHB/n53 ),
    .f({_al_u1967_o,_al_u1947_o}),
    .q({pnum3[16],pnum3[4]}));  // src/AHB.v(70)
  // src/AHB.v(70)
  // src/AHB.v(70)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg21_b17|U_AHB/reg21_b3  (
    .a({\PWM3/n24 ,\PWM3/n24 }),
    .b({\PWM3/n25_neg_lutinv ,\PWM3/n25_neg_lutinv }),
    .c({\PWM3/n26 [17],\PWM3/n26 [3]}),
    .clk(clk100m),
    .d({\PWM3/pnumr [17],\PWM3/pnumr [3]}),
    .mi({\U_AHB/h2h_hwdata [17],\U_AHB/h2h_hwdata [3]}),
    .sr(\U_AHB/n53 ),
    .f({_al_u1965_o,_al_u1949_o}),
    .q({pnum3[17],pnum3[3]}));  // src/AHB.v(70)
  // src/AHB.v(70)
  // src/AHB.v(70)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg21_b18|U_AHB/reg21_b23  (
    .a({\PWM3/n24 ,\PWM3/n24 }),
    .b({\PWM3/n25_neg_lutinv ,\PWM3/n25_neg_lutinv }),
    .c({\PWM3/n26 [18],\PWM3/n26 [23]}),
    .clk(clk100m),
    .d({\PWM3/pnumr [18],\PWM3/pnumr [23]}),
    .mi({\U_AHB/h2h_hwdata [18],\U_AHB/h2h_hwdata [23]}),
    .sr(\U_AHB/n53 ),
    .f({_al_u1963_o,_al_u1951_o}),
    .q({pnum3[18],pnum3[23]}));  // src/AHB.v(70)
  // src/AHB.v(70)
  // src/AHB.v(70)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg21_b19|U_AHB/reg21_b22  (
    .a({\PWM3/n24 ,\PWM3/n24 }),
    .b({\PWM3/n25_neg_lutinv ,\PWM3/n25_neg_lutinv }),
    .c({\PWM3/n26 [19],\PWM3/n26 [22]}),
    .clk(clk100m),
    .d({\PWM3/pnumr [19],\PWM3/pnumr [22]}),
    .mi({\U_AHB/h2h_hwdata [19],\U_AHB/h2h_hwdata [22]}),
    .sr(\U_AHB/n53 ),
    .f({_al_u1961_o,_al_u1953_o}),
    .q({pnum3[19],pnum3[22]}));  // src/AHB.v(70)
  // src/AHB.v(70)
  // src/AHB.v(70)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg21_b1|U_AHB/reg21_b21  (
    .a({\PWM3/n24 ,\PWM3/n24 }),
    .b({\PWM3/n25_neg_lutinv ,\PWM3/n25_neg_lutinv }),
    .c({\PWM3/n26 [1],\PWM3/n26 [21]}),
    .clk(clk100m),
    .d({\PWM3/pnumr [1],\PWM3/pnumr [21]}),
    .mi({\U_AHB/h2h_hwdata [1],\U_AHB/h2h_hwdata [21]}),
    .sr(\U_AHB/n53 ),
    .f({_al_u1981_o,_al_u1955_o}),
    .q({pnum3[1],pnum3[21]}));  // src/AHB.v(70)
  // src/AHB.v(70)
  // src/AHB.v(70)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg21_b27|U_AHB/reg21_b29  (
    .a({_al_u3192_o,_al_u3203_o}),
    .b({\U_AHB/n108 ,\U_AHB/n108 }),
    .c({\U_AHB/n105 ,\U_AHB/n105 }),
    .clk(clk100m),
    .d(pnumcnt8[21:20]),
    .e(pnumcnt9[21:20]),
    .mi({\U_AHB/h2h_hwdata [27],\U_AHB/h2h_hwdata [29]}),
    .sr(\U_AHB/n53 ),
    .f({_al_u3193_o,_al_u3204_o}),
    .q({pnum3[27],pnum3[29]}));  // src/AHB.v(70)
  // src/AHB.v(70)
  // src/AHB.v(70)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg21_b28|U_AHB/reg21_b31  (
    .a({_al_u3207_o,_al_u3229_o}),
    .b({\U_AHB/n96 ,\U_AHB/n96 }),
    .c({\U_AHB/n93 ,\U_AHB/n93 }),
    .clk(clk100m),
    .d(pnumcntF[20:19]),
    .e(pwm_state_read[4:3]),
    .mi({\U_AHB/h2h_hwdata [28],\U_AHB/h2h_hwdata [31]}),
    .sr(\U_AHB/n53 ),
    .f({_al_u3208_o,_al_u3230_o}),
    .q({pnum3[28],pnum3[31]}));  // src/AHB.v(70)
  // src/AHB.v(70)
  // src/AHB.v(70)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg21_b2|U_AHB/reg21_b20  (
    .a({\PWM3/n24 ,\PWM3/n24 }),
    .b({\PWM3/n25_neg_lutinv ,\PWM3/n25_neg_lutinv }),
    .c({\PWM3/n26 [2],\PWM3/n26 [20]}),
    .clk(clk100m),
    .d({\PWM3/pnumr [2],\PWM3/pnumr [20]}),
    .mi({\U_AHB/h2h_hwdata [2],\U_AHB/h2h_hwdata [20]}),
    .sr(\U_AHB/n53 ),
    .f({_al_u1959_o,_al_u1957_o}),
    .q({pnum3[2],pnum3[20]}));  // src/AHB.v(70)
  // src/AHB.v(71)
  // src/AHB.v(71)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b1010100000100000),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b1010100000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg22_b0|U_AHB/reg22_b30  (
    .a({\PWM4/n24 ,_al_u3273_o}),
    .b({\PWM4/n25_neg_lutinv ,\U_AHB/n96 }),
    .c({\PWM4/n26 [0],\U_AHB/n93 }),
    .clk(clk100m),
    .d({\PWM4/pnumr [0],pnumcntF[15]}),
    .e({open_n29308,pwm_state_read[15]}),
    .mi({\U_AHB/h2h_hwdata [0],\U_AHB/h2h_hwdata [30]}),
    .sr(\U_AHB/n55 ),
    .f({_al_u2065_o,_al_u3274_o}),
    .q({pnum4[0],pnum4[30]}));  // src/AHB.v(71)
  // src/AHB.v(71)
  // src/AHB.v(71)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b1010100000100000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1010100000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg22_b10|U_AHB/reg22_b27  (
    .a({\PWM4/n24 ,_al_u2503_o}),
    .b({\PWM4/n25_neg_lutinv ,pnumcntA[14]}),
    .c({\PWM4/n26 [10],pnumcntA[15]}),
    .clk(clk100m),
    .d({\PWM4/pnumr [10],pnumcntA[16]}),
    .e({open_n29325,pnumcntA[17]}),
    .mi({\U_AHB/h2h_hwdata [10],\U_AHB/h2h_hwdata [27]}),
    .sr(\U_AHB/n55 ),
    .f({_al_u2061_o,_al_u2504_o}),
    .q({pnum4[10],pnum4[27]}));  // src/AHB.v(71)
  // src/AHB.v(71)
  // src/AHB.v(71)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg22_b11|U_AHB/reg22_b32  (
    .a({\PWM4/n24 ,\PWM4/n24 }),
    .b({\PWM4/n25_neg_lutinv ,\PWM4/n25_neg_lutinv }),
    .c({\PWM4/n26 [11],\PWM4/n26 [9]}),
    .clk(clk100m),
    .d({\PWM4/pnumr [11],\PWM4/pnumr [9]}),
    .mi({\U_AHB/h2h_hwdata [11],1'b1}),
    .sr(\U_AHB/n55 ),
    .f({_al_u2059_o,_al_u2019_o}),
    .q({pnum4[11],pnum4[32]}));  // src/AHB.v(71)
  // src/AHB.v(71)
  // src/AHB.v(71)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg22_b12|U_AHB/reg22_b8  (
    .a({\PWM4/n24 ,\PWM4/n24 }),
    .b({\PWM4/n25_neg_lutinv ,\PWM4/n25_neg_lutinv }),
    .c({\PWM4/n26 [12],\PWM4/n26 [8]}),
    .clk(clk100m),
    .d({\PWM4/pnumr [12],\PWM4/pnumr [8]}),
    .mi({\U_AHB/h2h_hwdata [12],\U_AHB/h2h_hwdata [8]}),
    .sr(\U_AHB/n55 ),
    .f({_al_u2057_o,_al_u2021_o}),
    .q({pnum4[12],pnum4[8]}));  // src/AHB.v(71)
  // src/AHB.v(71)
  // src/AHB.v(71)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg22_b13|U_AHB/reg22_b7  (
    .a({\PWM4/n24 ,\PWM4/n24 }),
    .b({\PWM4/n25_neg_lutinv ,\PWM4/n25_neg_lutinv }),
    .c({\PWM4/n26 [13],\PWM4/n26 [7]}),
    .clk(clk100m),
    .d({\PWM4/pnumr [13],\PWM4/pnumr [7]}),
    .mi({\U_AHB/h2h_hwdata [13],\U_AHB/h2h_hwdata [7]}),
    .sr(\U_AHB/n55 ),
    .f({_al_u2055_o,_al_u2023_o}),
    .q({pnum4[13],pnum4[7]}));  // src/AHB.v(71)
  // src/AHB.v(71)
  // src/AHB.v(71)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg22_b14|U_AHB/reg22_b6  (
    .a({\PWM4/n24 ,\PWM4/n24 }),
    .b({\PWM4/n25_neg_lutinv ,\PWM4/n25_neg_lutinv }),
    .c({\PWM4/n26 [14],\PWM4/n26 [6]}),
    .clk(clk100m),
    .d({\PWM4/pnumr [14],\PWM4/pnumr [6]}),
    .mi({\U_AHB/h2h_hwdata [14],\U_AHB/h2h_hwdata [6]}),
    .sr(\U_AHB/n55 ),
    .f({_al_u2053_o,_al_u2025_o}),
    .q({pnum4[14],pnum4[6]}));  // src/AHB.v(71)
  // src/AHB.v(71)
  // src/AHB.v(71)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg22_b15|U_AHB/reg22_b5  (
    .a({\PWM4/n24 ,\PWM4/n24 }),
    .b({\PWM4/n25_neg_lutinv ,\PWM4/n25_neg_lutinv }),
    .c({\PWM4/n26 [15],\PWM4/n26 [5]}),
    .clk(clk100m),
    .d({\PWM4/pnumr [15],\PWM4/pnumr [5]}),
    .mi({\U_AHB/h2h_hwdata [15],\U_AHB/h2h_hwdata [5]}),
    .sr(\U_AHB/n55 ),
    .f({_al_u2051_o,_al_u2027_o}),
    .q({pnum4[15],pnum4[5]}));  // src/AHB.v(71)
  // src/AHB.v(71)
  // src/AHB.v(71)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg22_b16|U_AHB/reg22_b4  (
    .a({\PWM4/n24 ,\PWM4/n24 }),
    .b({\PWM4/n25_neg_lutinv ,\PWM4/n25_neg_lutinv }),
    .c({\PWM4/n26 [16],\PWM4/n26 [4]}),
    .clk(clk100m),
    .d({\PWM4/pnumr [16],\PWM4/pnumr [4]}),
    .mi({\U_AHB/h2h_hwdata [16],\U_AHB/h2h_hwdata [4]}),
    .sr(\U_AHB/n55 ),
    .f({_al_u2049_o,_al_u2029_o}),
    .q({pnum4[16],pnum4[4]}));  // src/AHB.v(71)
  // src/AHB.v(71)
  // src/AHB.v(71)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg22_b17|U_AHB/reg22_b3  (
    .a({\PWM4/n24 ,\PWM4/n24 }),
    .b({\PWM4/n25_neg_lutinv ,\PWM4/n25_neg_lutinv }),
    .c({\PWM4/n26 [17],\PWM4/n26 [3]}),
    .clk(clk100m),
    .d({\PWM4/pnumr [17],\PWM4/pnumr [3]}),
    .mi({\U_AHB/h2h_hwdata [17],\U_AHB/h2h_hwdata [3]}),
    .sr(\U_AHB/n55 ),
    .f({_al_u2047_o,_al_u2031_o}),
    .q({pnum4[17],pnum4[3]}));  // src/AHB.v(71)
  // src/AHB.v(71)
  // src/AHB.v(71)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg22_b18|U_AHB/reg22_b23  (
    .a({\PWM4/n24 ,\PWM4/n24 }),
    .b({\PWM4/n25_neg_lutinv ,\PWM4/n25_neg_lutinv }),
    .c({\PWM4/n26 [18],\PWM4/n26 [23]}),
    .clk(clk100m),
    .d({\PWM4/pnumr [18],\PWM4/pnumr [23]}),
    .mi({\U_AHB/h2h_hwdata [18],\U_AHB/h2h_hwdata [23]}),
    .sr(\U_AHB/n55 ),
    .f({_al_u2045_o,_al_u2033_o}),
    .q({pnum4[18],pnum4[23]}));  // src/AHB.v(71)
  // src/AHB.v(71)
  // src/AHB.v(71)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg22_b19|U_AHB/reg22_b22  (
    .a({\PWM4/n24 ,\PWM4/n24 }),
    .b({\PWM4/n25_neg_lutinv ,\PWM4/n25_neg_lutinv }),
    .c({\PWM4/n26 [19],\PWM4/n26 [22]}),
    .clk(clk100m),
    .d({\PWM4/pnumr [19],\PWM4/pnumr [22]}),
    .mi({\U_AHB/h2h_hwdata [19],\U_AHB/h2h_hwdata [22]}),
    .sr(\U_AHB/n55 ),
    .f({_al_u2043_o,_al_u2035_o}),
    .q({pnum4[19],pnum4[22]}));  // src/AHB.v(71)
  // src/AHB.v(71)
  // src/AHB.v(71)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg22_b1|U_AHB/reg22_b21  (
    .a({\PWM4/n24 ,\PWM4/n24 }),
    .b({\PWM4/n25_neg_lutinv ,\PWM4/n25_neg_lutinv }),
    .c({\PWM4/n26 [1],\PWM4/n26 [21]}),
    .clk(clk100m),
    .d({\PWM4/pnumr [1],\PWM4/pnumr [21]}),
    .mi({\U_AHB/h2h_hwdata [1],\U_AHB/h2h_hwdata [21]}),
    .sr(\U_AHB/n55 ),
    .f({_al_u2063_o,_al_u2037_o}),
    .q({pnum4[1],pnum4[21]}));  // src/AHB.v(71)
  // src/AHB.v(71)
  // src/AHB.v(71)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg22_b28|U_AHB/reg22_b25  (
    .a({_al_u3262_o,_al_u3251_o}),
    .b({\U_AHB/n96 ,\U_AHB/n96 }),
    .c({\U_AHB/n93 ,\U_AHB/n93 }),
    .clk(clk100m),
    .d({pnumcntF[16],pnumcntF[17]}),
    .e({pwm_state_read[0],pwm_state_read[1]}),
    .mi({\U_AHB/h2h_hwdata [28],\U_AHB/h2h_hwdata [25]}),
    .sr(\U_AHB/n55 ),
    .f({_al_u3263_o,_al_u3252_o}),
    .q({pnum4[28],pnum4[25]}));  // src/AHB.v(71)
  // src/AHB.v(71)
  // src/AHB.v(71)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg22_b29|U_AHB/reg22_b31  (
    .a({_al_u3258_o,_al_u3269_o}),
    .b({\U_AHB/n108 ,\U_AHB/n108 }),
    .c({\U_AHB/n105 ,\U_AHB/n105 }),
    .clk(clk100m),
    .d(pnumcnt8[16:15]),
    .e(pnumcnt9[16:15]),
    .mi({\U_AHB/h2h_hwdata [29],\U_AHB/h2h_hwdata [31]}),
    .sr(\U_AHB/n55 ),
    .f({_al_u3259_o,_al_u3270_o}),
    .q({pnum4[29],pnum4[31]}));  // src/AHB.v(71)
  // src/AHB.v(71)
  // src/AHB.v(71)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg22_b2|U_AHB/reg22_b20  (
    .a({\PWM4/n24 ,\PWM4/n24 }),
    .b({\PWM4/n25_neg_lutinv ,\PWM4/n25_neg_lutinv }),
    .c({\PWM4/n26 [2],\PWM4/n26 [20]}),
    .clk(clk100m),
    .d({\PWM4/pnumr [2],\PWM4/pnumr [20]}),
    .mi({\U_AHB/h2h_hwdata [2],\U_AHB/h2h_hwdata [20]}),
    .sr(\U_AHB/n55 ),
    .f({_al_u2041_o,_al_u2039_o}),
    .q({pnum4[2],pnum4[20]}));  // src/AHB.v(71)
  // src/AHB.v(72)
  // src/AHB.v(72)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b1010100000100000),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b1010100000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg23_b0|U_AHB/reg23_b28  (
    .a({\PWM5/n24 ,_al_u3291_o}),
    .b({\PWM5/n25_neg_lutinv ,\U_AHB/n108 }),
    .c({\PWM5/n26 [0],\U_AHB/n105 }),
    .clk(clk100m),
    .d({\PWM5/pnumr [0],pnumcnt8[13]}),
    .e({open_n29528,pnumcnt9[13]}),
    .mi({\U_AHB/h2h_hwdata [0],\U_AHB/h2h_hwdata [28]}),
    .sr(\U_AHB/n57 ),
    .f({_al_u2147_o,_al_u3292_o}),
    .q({pnum5[0],pnum5[28]}));  // src/AHB.v(72)
  // src/AHB.v(72)
  // src/AHB.v(72)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg23_b10|U_AHB/reg23_b32  (
    .a({\PWM5/n24 ,\PWM5/n24 }),
    .b({\PWM5/n25_neg_lutinv ,\PWM5/n25_neg_lutinv }),
    .c(\PWM5/n26 [10:9]),
    .clk(clk100m),
    .d(\PWM5/pnumr [10:9]),
    .mi({\U_AHB/h2h_hwdata [10],1'b1}),
    .sr(\U_AHB/n57 ),
    .f({_al_u2143_o,_al_u2101_o}),
    .q({pnum5[10],pnum5[32]}));  // src/AHB.v(72)
  // src/AHB.v(72)
  // src/AHB.v(72)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg23_b11|U_AHB/reg23_b8  (
    .a({\PWM5/n24 ,\PWM5/n24 }),
    .b({\PWM5/n25_neg_lutinv ,\PWM5/n25_neg_lutinv }),
    .c({\PWM5/n26 [11],\PWM5/n26 [8]}),
    .clk(clk100m),
    .d({\PWM5/pnumr [11],\PWM5/pnumr [8]}),
    .mi({\U_AHB/h2h_hwdata [11],\U_AHB/h2h_hwdata [8]}),
    .sr(\U_AHB/n57 ),
    .f({_al_u2141_o,_al_u2103_o}),
    .q({pnum5[11],pnum5[8]}));  // src/AHB.v(72)
  // src/AHB.v(72)
  // src/AHB.v(72)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg23_b12|U_AHB/reg23_b7  (
    .a({\PWM5/n24 ,\PWM5/n24 }),
    .b({\PWM5/n25_neg_lutinv ,\PWM5/n25_neg_lutinv }),
    .c({\PWM5/n26 [12],\PWM5/n26 [7]}),
    .clk(clk100m),
    .d({\PWM5/pnumr [12],\PWM5/pnumr [7]}),
    .mi({\U_AHB/h2h_hwdata [12],\U_AHB/h2h_hwdata [7]}),
    .sr(\U_AHB/n57 ),
    .f({_al_u2139_o,_al_u2105_o}),
    .q({pnum5[12],pnum5[7]}));  // src/AHB.v(72)
  // src/AHB.v(72)
  // src/AHB.v(72)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg23_b13|U_AHB/reg23_b6  (
    .a({\PWM5/n24 ,\PWM5/n24 }),
    .b({\PWM5/n25_neg_lutinv ,\PWM5/n25_neg_lutinv }),
    .c({\PWM5/n26 [13],\PWM5/n26 [6]}),
    .clk(clk100m),
    .d({\PWM5/pnumr [13],\PWM5/pnumr [6]}),
    .mi({\U_AHB/h2h_hwdata [13],\U_AHB/h2h_hwdata [6]}),
    .sr(\U_AHB/n57 ),
    .f({_al_u2137_o,_al_u2107_o}),
    .q({pnum5[13],pnum5[6]}));  // src/AHB.v(72)
  // src/AHB.v(72)
  // src/AHB.v(72)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg23_b14|U_AHB/reg23_b5  (
    .a({\PWM5/n24 ,\PWM5/n24 }),
    .b({\PWM5/n25_neg_lutinv ,\PWM5/n25_neg_lutinv }),
    .c({\PWM5/n26 [14],\PWM5/n26 [5]}),
    .clk(clk100m),
    .d({\PWM5/pnumr [14],\PWM5/pnumr [5]}),
    .mi({\U_AHB/h2h_hwdata [14],\U_AHB/h2h_hwdata [5]}),
    .sr(\U_AHB/n57 ),
    .f({_al_u2135_o,_al_u2109_o}),
    .q({pnum5[14],pnum5[5]}));  // src/AHB.v(72)
  // src/AHB.v(72)
  // src/AHB.v(72)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg23_b15|U_AHB/reg23_b4  (
    .a({\PWM5/n24 ,\PWM5/n24 }),
    .b({\PWM5/n25_neg_lutinv ,\PWM5/n25_neg_lutinv }),
    .c({\PWM5/n26 [15],\PWM5/n26 [4]}),
    .clk(clk100m),
    .d({\PWM5/pnumr [15],\PWM5/pnumr [4]}),
    .mi({\U_AHB/h2h_hwdata [15],\U_AHB/h2h_hwdata [4]}),
    .sr(\U_AHB/n57 ),
    .f({_al_u2133_o,_al_u2111_o}),
    .q({pnum5[15],pnum5[4]}));  // src/AHB.v(72)
  // src/AHB.v(72)
  // src/AHB.v(72)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg23_b16|U_AHB/reg23_b3  (
    .a({\PWM5/n24 ,\PWM5/n24 }),
    .b({\PWM5/n25_neg_lutinv ,\PWM5/n25_neg_lutinv }),
    .c({\PWM5/n26 [16],\PWM5/n26 [3]}),
    .clk(clk100m),
    .d({\PWM5/pnumr [16],\PWM5/pnumr [3]}),
    .mi({\U_AHB/h2h_hwdata [16],\U_AHB/h2h_hwdata [3]}),
    .sr(\U_AHB/n57 ),
    .f({_al_u2131_o,_al_u2113_o}),
    .q({pnum5[16],pnum5[3]}));  // src/AHB.v(72)
  // src/AHB.v(72)
  // src/AHB.v(72)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg23_b17|U_AHB/reg23_b23  (
    .a({\PWM5/n24 ,\PWM5/n24 }),
    .b({\PWM5/n25_neg_lutinv ,\PWM5/n25_neg_lutinv }),
    .c({\PWM5/n26 [17],\PWM5/n26 [23]}),
    .clk(clk100m),
    .d({\PWM5/pnumr [17],\PWM5/pnumr [23]}),
    .mi({\U_AHB/h2h_hwdata [17],\U_AHB/h2h_hwdata [23]}),
    .sr(\U_AHB/n57 ),
    .f({_al_u2129_o,_al_u2115_o}),
    .q({pnum5[17],pnum5[23]}));  // src/AHB.v(72)
  // src/AHB.v(72)
  // src/AHB.v(72)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg23_b18|U_AHB/reg23_b22  (
    .a({\PWM5/n24 ,\PWM5/n24 }),
    .b({\PWM5/n25_neg_lutinv ,\PWM5/n25_neg_lutinv }),
    .c({\PWM5/n26 [18],\PWM5/n26 [22]}),
    .clk(clk100m),
    .d({\PWM5/pnumr [18],\PWM5/pnumr [22]}),
    .mi({\U_AHB/h2h_hwdata [18],\U_AHB/h2h_hwdata [22]}),
    .sr(\U_AHB/n57 ),
    .f({_al_u2127_o,_al_u2117_o}),
    .q({pnum5[18],pnum5[22]}));  // src/AHB.v(72)
  // src/AHB.v(72)
  // src/AHB.v(72)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg23_b19|U_AHB/reg23_b21  (
    .a({\PWM5/n24 ,\PWM5/n24 }),
    .b({\PWM5/n25_neg_lutinv ,\PWM5/n25_neg_lutinv }),
    .c({\PWM5/n26 [19],\PWM5/n26 [21]}),
    .clk(clk100m),
    .d({\PWM5/pnumr [19],\PWM5/pnumr [21]}),
    .mi({\U_AHB/h2h_hwdata [19],\U_AHB/h2h_hwdata [21]}),
    .sr(\U_AHB/n57 ),
    .f({_al_u2125_o,_al_u2119_o}),
    .q({pnum5[19],pnum5[21]}));  // src/AHB.v(72)
  // src/AHB.v(72)
  // src/AHB.v(72)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg23_b1|U_AHB/reg23_b20  (
    .a({\PWM5/n24 ,\PWM5/n24 }),
    .b({\PWM5/n25_neg_lutinv ,\PWM5/n25_neg_lutinv }),
    .c({\PWM5/n26 [1],\PWM5/n26 [20]}),
    .clk(clk100m),
    .d({\PWM5/pnumr [1],\PWM5/pnumr [20]}),
    .mi({\U_AHB/h2h_hwdata [1],\U_AHB/h2h_hwdata [20]}),
    .sr(\U_AHB/n57 ),
    .f({_al_u2145_o,_al_u2121_o}),
    .q({pnum5[1],pnum5[20]}));  // src/AHB.v(72)
  // src/AHB.v(72)
  // src/AHB.v(72)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg23_b24|U_AHB/reg23_b2  (
    .a({open_n29698,\PWM5/n24 }),
    .b({limit_l_pad[14],\PWM5/n25_neg_lutinv }),
    .c({limit_r_pad[14],\PWM5/n26 [2]}),
    .clk(clk100m),
    .d({\PWME/n11 ,\PWM5/pnumr [2]}),
    .mi({\U_AHB/h2h_hwdata [24],\U_AHB/h2h_hwdata [2]}),
    .sr(\U_AHB/n57 ),
    .f({_al_u3050_o,_al_u2123_o}),
    .q({pnum5[24],pnum5[2]}));  // src/AHB.v(72)
  // src/AHB.v(72)
  // src/AHB.v(72)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(C*B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg23_b27|U_AHB/reg23_b9  (
    .b({limit_l_pad[13],limit_l_pad[10]}),
    .c({limit_r_pad[13],limit_r_pad[10]}),
    .clk(clk100m),
    .d({\PWMD/n11 ,\PWMA/n11 }),
    .mi({\U_AHB/h2h_hwdata [27],\U_AHB/h2h_hwdata [9]}),
    .sr(\U_AHB/n57 ),
    .f({_al_u3047_o,_al_u3038_o}),
    .q({pnum5[27],pnum5[9]}));  // src/AHB.v(72)
  // src/AHB.v(73)
  // src/AHB.v(73)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(D*C*~B*A)"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(D*C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0010000000000000),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0010000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg24_b0|U_AHB/reg24_b31  (
    .a({\U_AHB/h2h_hwrite ,_al_u3118_o}),
    .b({\U_AHB/h2h_haddr [13],\U_AHB/n96 }),
    .c({\U_AHB/h2h_haddr [14],\U_AHB/n93 }),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [6],pnumcntF[7]}),
    .e({open_n29730,pwm_state_read[7]}),
    .mi({\U_AHB/h2h_hwdata [0],\U_AHB/h2h_hwdata [31]}),
    .sr(\U_AHB/n59 ),
    .f({\U_AHB/n59 ,_al_u3119_o}),
    .q({pnum6[0],pnum6[31]}));  // src/AHB.v(73)
  // src/AHB.v(73)
  // src/AHB.v(73)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b1010100000100000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1010100000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg24_b10|U_AHB/reg24_b28  (
    .a({\PWM6/n24 ,_al_u2501_o}),
    .b({\PWM6/n25_neg_lutinv ,pnumcntA[6]}),
    .c({\PWM6/n26 [10],pnumcntA[7]}),
    .clk(clk100m),
    .d({\PWM6/pnumr [10],pnumcntA[8]}),
    .e({open_n29747,pnumcntA[9]}),
    .mi({\U_AHB/h2h_hwdata [10],\U_AHB/h2h_hwdata [28]}),
    .sr(\U_AHB/n59 ),
    .f({_al_u2225_o,_al_u2502_o}),
    .q({pnum6[10],pnum6[28]}));  // src/AHB.v(73)
  // src/AHB.v(73)
  // src/AHB.v(73)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg24_b11|U_AHB/reg24_b32  (
    .a({\PWM6/n24 ,\PWM6/n24 }),
    .b({\PWM6/n25_neg_lutinv ,\PWM6/n25_neg_lutinv }),
    .c({\PWM6/n26 [11],\PWM6/n26 [9]}),
    .clk(clk100m),
    .d({\PWM6/pnumr [11],\PWM6/pnumr [9]}),
    .mi({\U_AHB/h2h_hwdata [11],1'b1}),
    .sr(\U_AHB/n59 ),
    .f({_al_u2223_o,_al_u2183_o}),
    .q({pnum6[11],pnum6[32]}));  // src/AHB.v(73)
  // src/AHB.v(73)
  // src/AHB.v(73)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg24_b12|U_AHB/reg24_b8  (
    .a({\PWM6/n24 ,\PWM6/n24 }),
    .b({\PWM6/n25_neg_lutinv ,\PWM6/n25_neg_lutinv }),
    .c({\PWM6/n26 [12],\PWM6/n26 [8]}),
    .clk(clk100m),
    .d({\PWM6/pnumr [12],\PWM6/pnumr [8]}),
    .mi({\U_AHB/h2h_hwdata [12],\U_AHB/h2h_hwdata [8]}),
    .sr(\U_AHB/n59 ),
    .f({_al_u2221_o,_al_u2185_o}),
    .q({pnum6[12],pnum6[8]}));  // src/AHB.v(73)
  // src/AHB.v(73)
  // src/AHB.v(73)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg24_b13|U_AHB/reg24_b7  (
    .a({\PWM6/n24 ,\PWM6/n24 }),
    .b({\PWM6/n25_neg_lutinv ,\PWM6/n25_neg_lutinv }),
    .c({\PWM6/n26 [13],\PWM6/n26 [7]}),
    .clk(clk100m),
    .d({\PWM6/pnumr [13],\PWM6/pnumr [7]}),
    .mi({\U_AHB/h2h_hwdata [13],\U_AHB/h2h_hwdata [7]}),
    .sr(\U_AHB/n59 ),
    .f({_al_u2219_o,_al_u2187_o}),
    .q({pnum6[13],pnum6[7]}));  // src/AHB.v(73)
  // src/AHB.v(73)
  // src/AHB.v(73)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg24_b14|U_AHB/reg24_b6  (
    .a({\PWM6/n24 ,\PWM6/n24 }),
    .b({\PWM6/n25_neg_lutinv ,\PWM6/n25_neg_lutinv }),
    .c({\PWM6/n26 [14],\PWM6/n26 [6]}),
    .clk(clk100m),
    .d({\PWM6/pnumr [14],\PWM6/pnumr [6]}),
    .mi({\U_AHB/h2h_hwdata [14],\U_AHB/h2h_hwdata [6]}),
    .sr(\U_AHB/n59 ),
    .f({_al_u2217_o,_al_u2189_o}),
    .q({pnum6[14],pnum6[6]}));  // src/AHB.v(73)
  // src/AHB.v(73)
  // src/AHB.v(73)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg24_b15|U_AHB/reg24_b5  (
    .a({\PWM6/n24 ,\PWM6/n24 }),
    .b({\PWM6/n25_neg_lutinv ,\PWM6/n25_neg_lutinv }),
    .c({\PWM6/n26 [15],\PWM6/n26 [5]}),
    .clk(clk100m),
    .d({\PWM6/pnumr [15],\PWM6/pnumr [5]}),
    .mi({\U_AHB/h2h_hwdata [15],\U_AHB/h2h_hwdata [5]}),
    .sr(\U_AHB/n59 ),
    .f({_al_u2215_o,_al_u2191_o}),
    .q({pnum6[15],pnum6[5]}));  // src/AHB.v(73)
  // src/AHB.v(73)
  // src/AHB.v(73)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg24_b16|U_AHB/reg24_b4  (
    .a({\PWM6/n24 ,\PWM6/n24 }),
    .b({\PWM6/n25_neg_lutinv ,\PWM6/n25_neg_lutinv }),
    .c({\PWM6/n26 [16],\PWM6/n26 [4]}),
    .clk(clk100m),
    .d({\PWM6/pnumr [16],\PWM6/pnumr [4]}),
    .mi({\U_AHB/h2h_hwdata [16],\U_AHB/h2h_hwdata [4]}),
    .sr(\U_AHB/n59 ),
    .f({_al_u2213_o,_al_u2193_o}),
    .q({pnum6[16],pnum6[4]}));  // src/AHB.v(73)
  // src/AHB.v(73)
  // src/AHB.v(73)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg24_b17|U_AHB/reg24_b3  (
    .a({\PWM6/n24 ,\PWM6/n24 }),
    .b({\PWM6/n25_neg_lutinv ,\PWM6/n25_neg_lutinv }),
    .c({\PWM6/n26 [17],\PWM6/n26 [3]}),
    .clk(clk100m),
    .d({\PWM6/pnumr [17],\PWM6/pnumr [3]}),
    .mi({\U_AHB/h2h_hwdata [17],\U_AHB/h2h_hwdata [3]}),
    .sr(\U_AHB/n59 ),
    .f({_al_u2211_o,_al_u2195_o}),
    .q({pnum6[17],pnum6[3]}));  // src/AHB.v(73)
  // src/AHB.v(73)
  // src/AHB.v(73)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg24_b18|U_AHB/reg24_b23  (
    .a({\PWM6/n24 ,\PWM6/n24 }),
    .b({\PWM6/n25_neg_lutinv ,\PWM6/n25_neg_lutinv }),
    .c({\PWM6/n26 [18],\PWM6/n26 [23]}),
    .clk(clk100m),
    .d({\PWM6/pnumr [18],\PWM6/pnumr [23]}),
    .mi({\U_AHB/h2h_hwdata [18],\U_AHB/h2h_hwdata [23]}),
    .sr(\U_AHB/n59 ),
    .f({_al_u2209_o,_al_u2197_o}),
    .q({pnum6[18],pnum6[23]}));  // src/AHB.v(73)
  // src/AHB.v(73)
  // src/AHB.v(73)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg24_b19|U_AHB/reg24_b22  (
    .a({\PWM6/n24 ,\PWM6/n24 }),
    .b({\PWM6/n25_neg_lutinv ,\PWM6/n25_neg_lutinv }),
    .c({\PWM6/n26 [19],\PWM6/n26 [22]}),
    .clk(clk100m),
    .d({\PWM6/pnumr [19],\PWM6/pnumr [22]}),
    .mi({\U_AHB/h2h_hwdata [19],\U_AHB/h2h_hwdata [22]}),
    .sr(\U_AHB/n59 ),
    .f({_al_u2207_o,_al_u2199_o}),
    .q({pnum6[19],pnum6[22]}));  // src/AHB.v(73)
  // src/AHB.v(73)
  // src/AHB.v(73)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg24_b1|U_AHB/reg24_b21  (
    .a({\PWM6/n24 ,\PWM6/n24 }),
    .b({\PWM6/n25_neg_lutinv ,\PWM6/n25_neg_lutinv }),
    .c({\PWM6/n26 [1],\PWM6/n26 [21]}),
    .clk(clk100m),
    .d({\PWM6/pnumr [1],\PWM6/pnumr [21]}),
    .mi({\U_AHB/h2h_hwdata [1],\U_AHB/h2h_hwdata [21]}),
    .sr(\U_AHB/n59 ),
    .f({_al_u2227_o,_al_u2201_o}),
    .q({pnum6[1],pnum6[21]}));  // src/AHB.v(73)
  // src/AHB.v(73)
  // src/AHB.v(73)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg24_b24|U_AHB/reg24_b9  (
    .a({_al_u3324_o,_al_u3114_o}),
    .b({\U_AHB/n108 ,\U_AHB/n108 }),
    .c({\U_AHB/n105 ,\U_AHB/n105 }),
    .clk(clk100m),
    .d({pnumcnt8[10],pnumcnt8[7]}),
    .e({pnumcnt9[10],pnumcnt9[7]}),
    .mi({\U_AHB/h2h_hwdata [24],\U_AHB/h2h_hwdata [9]}),
    .sr(\U_AHB/n59 ),
    .f({_al_u3325_o,_al_u3115_o}),
    .q({pnum6[24],pnum6[9]}));  // src/AHB.v(73)
  // src/AHB.v(73)
  // src/AHB.v(73)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg24_b27|U_AHB/reg24_b30  (
    .a({_al_u3089_o,_al_u3103_o}),
    .b({\U_AHB/n108 ,\U_AHB/n108 }),
    .c({\U_AHB/n105 ,\U_AHB/n105 }),
    .clk(clk100m),
    .d(pnumcnt8[9:8]),
    .e(pnumcnt9[9:8]),
    .mi({\U_AHB/h2h_hwdata [27],\U_AHB/h2h_hwdata [30]}),
    .sr(\U_AHB/n59 ),
    .f({_al_u3092_o,_al_u3104_o}),
    .q({pnum6[27],pnum6[30]}));  // src/AHB.v(73)
  // src/AHB.v(73)
  // src/AHB.v(73)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg24_b29|U_AHB/reg24_b25  (
    .a({_al_u3107_o,_al_u3096_o}),
    .b({\U_AHB/n96 ,\U_AHB/n96 }),
    .c({\U_AHB/n93 ,\U_AHB/n93 }),
    .clk(clk100m),
    .d({pnumcntF[8],pnumcntF[9]}),
    .e({pwm_state_read[8],pwm_state_read[9]}),
    .mi({\U_AHB/h2h_hwdata [29],\U_AHB/h2h_hwdata [25]}),
    .sr(\U_AHB/n59 ),
    .f({_al_u3108_o,_al_u3097_o}),
    .q({pnum6[29],pnum6[25]}));  // src/AHB.v(73)
  // src/AHB.v(73)
  // src/AHB.v(73)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg24_b2|U_AHB/reg24_b20  (
    .a({\PWM6/n24 ,\PWM6/n24 }),
    .b({\PWM6/n25_neg_lutinv ,\PWM6/n25_neg_lutinv }),
    .c({\PWM6/n26 [2],\PWM6/n26 [20]}),
    .clk(clk100m),
    .d({\PWM6/pnumr [2],\PWM6/pnumr [20]}),
    .mi({\U_AHB/h2h_hwdata [2],\U_AHB/h2h_hwdata [20]}),
    .sr(\U_AHB/n59 ),
    .f({_al_u2205_o,_al_u2203_o}),
    .q({pnum6[2],pnum6[20]}));  // src/AHB.v(73)
  // src/AHB.v(74)
  // src/AHB.v(74)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*~B*D)"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*~B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0011000000000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b0011000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg25_b0|U_AHB/reg25_b1  (
    .b({\U_AHB/h2h_haddr [7],open_n29967}),
    .c(\U_AHB/h2h_haddr [8:7]),
    .clk(clk100m),
    .d({\U_AHB/n95_lutinv ,\U_AHB/n95_lutinv }),
    .mi({\U_AHB/h2h_hwdata [0],\U_AHB/h2h_hwdata [1]}),
    .sr(\U_AHB/n61 ),
    .f({\U_AHB/n99 ,\U_AHB/n96 }),
    .q({pnum7[0],pnum7[1]}));  // src/AHB.v(74)
  // src/AHB.v(74)
  // src/AHB.v(74)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg25_b10|U_AHB/reg25_b32  (
    .a({\PWM7/n24 ,\PWM7/n24 }),
    .b({\PWM7/n25_neg_lutinv ,\PWM7/n25_neg_lutinv }),
    .c(\PWM7/n26 [10:9]),
    .clk(clk100m),
    .d(\PWM7/pnumr [10:9]),
    .mi({\U_AHB/h2h_hwdata [10],1'b1}),
    .sr(\U_AHB/n61 ),
    .f({_al_u2305_o,_al_u2263_o}),
    .q({pnum7[10],pnum7[32]}));  // src/AHB.v(74)
  // src/AHB.v(74)
  // src/AHB.v(74)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg25_b11|U_AHB/reg25_b8  (
    .a({\PWM7/n24 ,\PWM7/n24 }),
    .b({\PWM7/n25_neg_lutinv ,\PWM7/n25_neg_lutinv }),
    .c({\PWM7/n26 [11],\PWM7/n26 [8]}),
    .clk(clk100m),
    .d({\PWM7/pnumr [11],\PWM7/pnumr [8]}),
    .mi({\U_AHB/h2h_hwdata [11],\U_AHB/h2h_hwdata [8]}),
    .sr(\U_AHB/n61 ),
    .f({_al_u2303_o,_al_u2265_o}),
    .q({pnum7[11],pnum7[8]}));  // src/AHB.v(74)
  // src/AHB.v(74)
  // src/AHB.v(74)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg25_b12|U_AHB/reg25_b7  (
    .a({\PWM7/n24 ,\PWM7/n24 }),
    .b({\PWM7/n25_neg_lutinv ,\PWM7/n25_neg_lutinv }),
    .c({\PWM7/n26 [12],\PWM7/n26 [7]}),
    .clk(clk100m),
    .d({\PWM7/pnumr [12],\PWM7/pnumr [7]}),
    .mi({\U_AHB/h2h_hwdata [12],\U_AHB/h2h_hwdata [7]}),
    .sr(\U_AHB/n61 ),
    .f({_al_u2301_o,_al_u2267_o}),
    .q({pnum7[12],pnum7[7]}));  // src/AHB.v(74)
  // src/AHB.v(74)
  // src/AHB.v(74)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg25_b13|U_AHB/reg25_b6  (
    .a({\PWM7/n24 ,\PWM7/n24 }),
    .b({\PWM7/n25_neg_lutinv ,\PWM7/n25_neg_lutinv }),
    .c({\PWM7/n26 [13],\PWM7/n26 [6]}),
    .clk(clk100m),
    .d({\PWM7/pnumr [13],\PWM7/pnumr [6]}),
    .mi({\U_AHB/h2h_hwdata [13],\U_AHB/h2h_hwdata [6]}),
    .sr(\U_AHB/n61 ),
    .f({_al_u2299_o,_al_u2269_o}),
    .q({pnum7[13],pnum7[6]}));  // src/AHB.v(74)
  // src/AHB.v(74)
  // src/AHB.v(74)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg25_b14|U_AHB/reg25_b5  (
    .a({\PWM7/n24 ,\PWM7/n24 }),
    .b({\PWM7/n25_neg_lutinv ,\PWM7/n25_neg_lutinv }),
    .c({\PWM7/n26 [14],\PWM7/n26 [5]}),
    .clk(clk100m),
    .d({\PWM7/pnumr [14],\PWM7/pnumr [5]}),
    .mi({\U_AHB/h2h_hwdata [14],\U_AHB/h2h_hwdata [5]}),
    .sr(\U_AHB/n61 ),
    .f({_al_u2297_o,_al_u2271_o}),
    .q({pnum7[14],pnum7[5]}));  // src/AHB.v(74)
  // src/AHB.v(74)
  // src/AHB.v(74)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg25_b15|U_AHB/reg25_b4  (
    .a({\PWM7/n24 ,\PWM7/n24 }),
    .b({\PWM7/n25_neg_lutinv ,\PWM7/n25_neg_lutinv }),
    .c({\PWM7/n26 [15],\PWM7/n26 [4]}),
    .clk(clk100m),
    .d({\PWM7/pnumr [15],\PWM7/pnumr [4]}),
    .mi({\U_AHB/h2h_hwdata [15],\U_AHB/h2h_hwdata [4]}),
    .sr(\U_AHB/n61 ),
    .f({_al_u2295_o,_al_u2273_o}),
    .q({pnum7[15],pnum7[4]}));  // src/AHB.v(74)
  // src/AHB.v(74)
  // src/AHB.v(74)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg25_b16|U_AHB/reg25_b3  (
    .a({\PWM7/n24 ,\PWM7/n24 }),
    .b({\PWM7/n25_neg_lutinv ,\PWM7/n25_neg_lutinv }),
    .c({\PWM7/n26 [16],\PWM7/n26 [3]}),
    .clk(clk100m),
    .d({\PWM7/pnumr [16],\PWM7/pnumr [3]}),
    .mi({\U_AHB/h2h_hwdata [16],\U_AHB/h2h_hwdata [3]}),
    .sr(\U_AHB/n61 ),
    .f({_al_u2293_o,_al_u2275_o}),
    .q({pnum7[16],pnum7[3]}));  // src/AHB.v(74)
  // src/AHB.v(74)
  // src/AHB.v(74)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg25_b17|U_AHB/reg25_b23  (
    .a({\PWM7/n24 ,\PWM7/n24 }),
    .b({\PWM7/n25_neg_lutinv ,\PWM7/n25_neg_lutinv }),
    .c({\PWM7/n26 [17],\PWM7/n26 [23]}),
    .clk(clk100m),
    .d({\PWM7/pnumr [17],\PWM7/pnumr [23]}),
    .mi({\U_AHB/h2h_hwdata [17],\U_AHB/h2h_hwdata [23]}),
    .sr(\U_AHB/n61 ),
    .f({_al_u2291_o,_al_u2277_o}),
    .q({pnum7[17],pnum7[23]}));  // src/AHB.v(74)
  // src/AHB.v(74)
  // src/AHB.v(74)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg25_b18|U_AHB/reg25_b22  (
    .a({\PWM7/n24 ,\PWM7/n24 }),
    .b({\PWM7/n25_neg_lutinv ,\PWM7/n25_neg_lutinv }),
    .c({\PWM7/n26 [18],\PWM7/n26 [22]}),
    .clk(clk100m),
    .d({\PWM7/pnumr [18],\PWM7/pnumr [22]}),
    .mi({\U_AHB/h2h_hwdata [18],\U_AHB/h2h_hwdata [22]}),
    .sr(\U_AHB/n61 ),
    .f({_al_u2289_o,_al_u2279_o}),
    .q({pnum7[18],pnum7[22]}));  // src/AHB.v(74)
  // src/AHB.v(74)
  // src/AHB.v(74)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg25_b19|U_AHB/reg25_b21  (
    .a({\PWM7/n24 ,\PWM7/n24 }),
    .b({\PWM7/n25_neg_lutinv ,\PWM7/n25_neg_lutinv }),
    .c({\PWM7/n26 [19],\PWM7/n26 [21]}),
    .clk(clk100m),
    .d({\PWM7/pnumr [19],\PWM7/pnumr [21]}),
    .mi({\U_AHB/h2h_hwdata [19],\U_AHB/h2h_hwdata [21]}),
    .sr(\U_AHB/n61 ),
    .f({_al_u2287_o,_al_u2281_o}),
    .q({pnum7[19],pnum7[21]}));  // src/AHB.v(74)
  // src/AHB.v(74)
  // src/AHB.v(74)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg25_b27|U_AHB/reg25_b25  (
    .a({_al_u3136_o,_al_u3125_o}),
    .b({\U_AHB/n108 ,\U_AHB/n108 }),
    .c({\U_AHB/n105 ,\U_AHB/n105 }),
    .clk(clk100m),
    .d({pnumcnt8[5],pnumcnt8[6]}),
    .e({pnumcnt9[5],pnumcnt9[6]}),
    .mi({\U_AHB/h2h_hwdata [27],\U_AHB/h2h_hwdata [25]}),
    .sr(\U_AHB/n61 ),
    .f({_al_u3137_o,_al_u3126_o}),
    .q({pnum7[27],pnum7[25]}));  // src/AHB.v(74)
  // src/AHB.v(74)
  // src/AHB.v(74)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg25_b29|U_AHB/reg25_b24  (
    .a({_al_u3152_o,_al_u3129_o}),
    .b({\U_AHB/n96 ,\U_AHB/n96 }),
    .c({\U_AHB/n93 ,\U_AHB/n93 }),
    .clk(clk100m),
    .d({pnumcntF[4],pnumcntF[6]}),
    .e({pwm_state_read[4],pwm_state_read[6]}),
    .mi({\U_AHB/h2h_hwdata [29],\U_AHB/h2h_hwdata [24]}),
    .sr(\U_AHB/n61 ),
    .f({_al_u3153_o,_al_u3130_o}),
    .q({pnum7[29],pnum7[24]}));  // src/AHB.v(74)
  // src/AHB.v(74)
  // src/AHB.v(74)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg25_b2|U_AHB/reg25_b20  (
    .a({\PWM7/n24 ,\PWM7/n24 }),
    .b({\PWM7/n25_neg_lutinv ,\PWM7/n25_neg_lutinv }),
    .c({\PWM7/n26 [2],\PWM7/n26 [20]}),
    .clk(clk100m),
    .d({\PWM7/pnumr [2],\PWM7/pnumr [20]}),
    .mi({\U_AHB/h2h_hwdata [2],\U_AHB/h2h_hwdata [20]}),
    .sr(\U_AHB/n61 ),
    .f({_al_u2285_o,_al_u2283_o}),
    .q({pnum7[2],pnum7[20]}));  // src/AHB.v(74)
  // src/AHB.v(75)
  // src/AHB.v(75)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg26_b0|U_AHB/reg26_b32  (
    .a({\PWM8/n24 ,\PWM8/n24 }),
    .b({\PWM8/n25_neg_lutinv ,\PWM8/n25_neg_lutinv }),
    .c({\PWM8/n26 [0],\PWM8/n26 [9]}),
    .clk(clk100m),
    .d({\PWM8/pnumr [0],\PWM8/pnumr [9]}),
    .mi({\U_AHB/h2h_hwdata [0],1'b1}),
    .sr(\U_AHB/n63 ),
    .f({_al_u2391_o,_al_u2345_o}),
    .q({pnum8[0],pnum8[32]}));  // src/AHB.v(75)
  // src/AHB.v(75)
  // src/AHB.v(75)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg26_b10|U_AHB/reg26_b8  (
    .a({\PWM8/n24 ,\PWM8/n24 }),
    .b({\PWM8/n25_neg_lutinv ,\PWM8/n25_neg_lutinv }),
    .c({\PWM8/n26 [10],\PWM8/n26 [8]}),
    .clk(clk100m),
    .d({\PWM8/pnumr [10],\PWM8/pnumr [8]}),
    .mi({\U_AHB/h2h_hwdata [10],\U_AHB/h2h_hwdata [8]}),
    .sr(\U_AHB/n63 ),
    .f({_al_u2387_o,_al_u2347_o}),
    .q({pnum8[10],pnum8[8]}));  // src/AHB.v(75)
  // src/AHB.v(75)
  // src/AHB.v(75)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg26_b11|U_AHB/reg26_b7  (
    .a({\PWM8/n24 ,\PWM8/n24 }),
    .b({\PWM8/n25_neg_lutinv ,\PWM8/n25_neg_lutinv }),
    .c({\PWM8/n26 [11],\PWM8/n26 [7]}),
    .clk(clk100m),
    .d({\PWM8/pnumr [11],\PWM8/pnumr [7]}),
    .mi({\U_AHB/h2h_hwdata [11],\U_AHB/h2h_hwdata [7]}),
    .sr(\U_AHB/n63 ),
    .f({_al_u2385_o,_al_u2349_o}),
    .q({pnum8[11],pnum8[7]}));  // src/AHB.v(75)
  // src/AHB.v(75)
  // src/AHB.v(75)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg26_b12|U_AHB/reg26_b6  (
    .a({\PWM8/n24 ,\PWM8/n24 }),
    .b({\PWM8/n25_neg_lutinv ,\PWM8/n25_neg_lutinv }),
    .c({\PWM8/n26 [12],\PWM8/n26 [6]}),
    .clk(clk100m),
    .d({\PWM8/pnumr [12],\PWM8/pnumr [6]}),
    .mi({\U_AHB/h2h_hwdata [12],\U_AHB/h2h_hwdata [6]}),
    .sr(\U_AHB/n63 ),
    .f({_al_u2383_o,_al_u2351_o}),
    .q({pnum8[12],pnum8[6]}));  // src/AHB.v(75)
  // src/AHB.v(75)
  // src/AHB.v(75)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg26_b13|U_AHB/reg26_b5  (
    .a({\PWM8/n24 ,\PWM8/n24 }),
    .b({\PWM8/n25_neg_lutinv ,\PWM8/n25_neg_lutinv }),
    .c({\PWM8/n26 [13],\PWM8/n26 [5]}),
    .clk(clk100m),
    .d({\PWM8/pnumr [13],\PWM8/pnumr [5]}),
    .mi({\U_AHB/h2h_hwdata [13],\U_AHB/h2h_hwdata [5]}),
    .sr(\U_AHB/n63 ),
    .f({_al_u2381_o,_al_u2353_o}),
    .q({pnum8[13],pnum8[5]}));  // src/AHB.v(75)
  // src/AHB.v(75)
  // src/AHB.v(75)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg26_b14|U_AHB/reg26_b4  (
    .a({\PWM8/n24 ,\PWM8/n24 }),
    .b({\PWM8/n25_neg_lutinv ,\PWM8/n25_neg_lutinv }),
    .c({\PWM8/n26 [14],\PWM8/n26 [4]}),
    .clk(clk100m),
    .d({\PWM8/pnumr [14],\PWM8/pnumr [4]}),
    .mi({\U_AHB/h2h_hwdata [14],\U_AHB/h2h_hwdata [4]}),
    .sr(\U_AHB/n63 ),
    .f({_al_u2379_o,_al_u2355_o}),
    .q({pnum8[14],pnum8[4]}));  // src/AHB.v(75)
  // src/AHB.v(75)
  // src/AHB.v(75)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg26_b15|U_AHB/reg26_b3  (
    .a({\PWM8/n24 ,\PWM8/n24 }),
    .b({\PWM8/n25_neg_lutinv ,\PWM8/n25_neg_lutinv }),
    .c({\PWM8/n26 [15],\PWM8/n26 [3]}),
    .clk(clk100m),
    .d({\PWM8/pnumr [15],\PWM8/pnumr [3]}),
    .mi({\U_AHB/h2h_hwdata [15],\U_AHB/h2h_hwdata [3]}),
    .sr(\U_AHB/n63 ),
    .f({_al_u2377_o,_al_u2357_o}),
    .q({pnum8[15],pnum8[3]}));  // src/AHB.v(75)
  // src/AHB.v(75)
  // src/AHB.v(75)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg26_b16|U_AHB/reg26_b23  (
    .a({\PWM8/n24 ,\PWM8/n24 }),
    .b({\PWM8/n25_neg_lutinv ,\PWM8/n25_neg_lutinv }),
    .c({\PWM8/n26 [16],\PWM8/n26 [23]}),
    .clk(clk100m),
    .d({\PWM8/pnumr [16],\PWM8/pnumr [23]}),
    .mi({\U_AHB/h2h_hwdata [16],\U_AHB/h2h_hwdata [23]}),
    .sr(\U_AHB/n63 ),
    .f({_al_u2375_o,_al_u2359_o}),
    .q({pnum8[16],pnum8[23]}));  // src/AHB.v(75)
  // src/AHB.v(75)
  // src/AHB.v(75)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg26_b17|U_AHB/reg26_b22  (
    .a({\PWM8/n24 ,\PWM8/n24 }),
    .b({\PWM8/n25_neg_lutinv ,\PWM8/n25_neg_lutinv }),
    .c({\PWM8/n26 [17],\PWM8/n26 [22]}),
    .clk(clk100m),
    .d({\PWM8/pnumr [17],\PWM8/pnumr [22]}),
    .mi({\U_AHB/h2h_hwdata [17],\U_AHB/h2h_hwdata [22]}),
    .sr(\U_AHB/n63 ),
    .f({_al_u2373_o,_al_u2361_o}),
    .q({pnum8[17],pnum8[22]}));  // src/AHB.v(75)
  // src/AHB.v(75)
  // src/AHB.v(75)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg26_b18|U_AHB/reg26_b21  (
    .a({\PWM8/n24 ,\PWM8/n24 }),
    .b({\PWM8/n25_neg_lutinv ,\PWM8/n25_neg_lutinv }),
    .c({\PWM8/n26 [18],\PWM8/n26 [21]}),
    .clk(clk100m),
    .d({\PWM8/pnumr [18],\PWM8/pnumr [21]}),
    .mi({\U_AHB/h2h_hwdata [18],\U_AHB/h2h_hwdata [21]}),
    .sr(\U_AHB/n63 ),
    .f({_al_u2371_o,_al_u2363_o}),
    .q({pnum8[18],pnum8[21]}));  // src/AHB.v(75)
  // src/AHB.v(75)
  // src/AHB.v(75)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg26_b19|U_AHB/reg26_b20  (
    .a({\PWM8/n24 ,\PWM8/n24 }),
    .b({\PWM8/n25_neg_lutinv ,\PWM8/n25_neg_lutinv }),
    .c({\PWM8/n26 [19],\PWM8/n26 [20]}),
    .clk(clk100m),
    .d({\PWM8/pnumr [19],\PWM8/pnumr [20]}),
    .mi({\U_AHB/h2h_hwdata [19],\U_AHB/h2h_hwdata [20]}),
    .sr(\U_AHB/n63 ),
    .f({_al_u2369_o,_al_u2365_o}),
    .q({pnum8[19],pnum8[20]}));  // src/AHB.v(75)
  // src/AHB.v(75)
  // src/AHB.v(75)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg26_b1|U_AHB/reg26_b2  (
    .a({\PWM8/n24 ,\PWM8/n24 }),
    .b({\PWM8/n25_neg_lutinv ,\PWM8/n25_neg_lutinv }),
    .c({\PWM8/n26 [1],\PWM8/n26 [2]}),
    .clk(clk100m),
    .d({\PWM8/pnumr [1],\PWM8/pnumr [2]}),
    .mi({\U_AHB/h2h_hwdata [1],\U_AHB/h2h_hwdata [2]}),
    .sr(\U_AHB/n63 ),
    .f({_al_u2389_o,_al_u2367_o}),
    .q({pnum8[1],pnum8[2]}));  // src/AHB.v(75)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg26_b24  (
    .a({open_n30340,_al_u3218_o}),
    .b({open_n30341,\U_AHB/n96 }),
    .c({open_n30342,\U_AHB/n93 }),
    .clk(clk100m),
    .d({open_n30344,pnumcntF[2]}),
    .e({open_n30345,pwm_state_read[2]}),
    .mi({open_n30347,\U_AHB/h2h_hwdata [24]}),
    .sr(\U_AHB/n63 ),
    .f({open_n30359,_al_u3219_o}),
    .q({open_n30363,pnum8[24]}));  // src/AHB.v(75)
  // src/AHB.v(75)
  // src/AHB.v(75)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg26_b25|U_AHB/reg26_b26  (
    .a({_al_u3214_o,_al_u3335_o}),
    .b({\U_AHB/n108 ,\U_AHB/n108 }),
    .c({\U_AHB/n105 ,\U_AHB/n105 }),
    .clk(clk100m),
    .d(pnumcnt8[2:1]),
    .e(pnumcnt9[2:1]),
    .mi({\U_AHB/h2h_hwdata [25],\U_AHB/h2h_hwdata [26]}),
    .sr(\U_AHB/n63 ),
    .f({_al_u3215_o,_al_u3336_o}),
    .q({pnum8[25],pnum8[26]}));  // src/AHB.v(75)
  // src/AHB.v(75)
  // src/AHB.v(75)
  EF2_PHY_MSLICE #(
    //.LUT0("(~D*C*B*A)"),
    //.LUT1("(C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000010000000),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg26_b31|U_AHB/reg26_b28  (
    .a({open_n30380,_al_u2502_o}),
    .b({open_n30381,_al_u2504_o}),
    .c({pwm_state_read[15],_al_u2505_o}),
    .clk(clk100m),
    .d({_al_u2978_o,pnumcntA[0]}),
    .mi({\U_AHB/h2h_hwdata [31],\U_AHB/h2h_hwdata [28]}),
    .sr(\U_AHB/n63 ),
    .f({\PWMF/u14_sel_is_1_o ,\PWMA/n25_neg_lutinv }),
    .q({pnum8[31],pnum8[28]}));  // src/AHB.v(75)
  // src/AHB.v(76)
  // src/AHB.v(76)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~(D*C*B*A))"),
    //.LUTF1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("(~1*~(D*C*B*A))"),
    //.LUTG1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111111111111111),
    .INIT_LUTF1(16'b1010100000100000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1010100000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg27_b0|U_AHB/reg27_b31  (
    .a({\PWM9/n24 ,_al_u2420_o}),
    .b({\PWM9/n25_neg_lutinv ,_al_u2422_o}),
    .c({\PWM9/n26 [0],_al_u2423_o}),
    .clk(clk100m),
    .d({\PWM9/pnumr [0],pnumcnt9[0]}),
    .e({open_n30397,\PWM9/stopreq }),
    .mi({\U_AHB/h2h_hwdata [0],\U_AHB/h2h_hwdata [31]}),
    .sr(\U_AHB/n65 ),
    .f({_al_u2471_o,_al_u3034_o}),
    .q({pnum9[0],pnum9[31]}));  // src/AHB.v(76)
  // src/AHB.v(76)
  // src/AHB.v(76)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg27_b10|U_AHB/reg27_b32  (
    .a({\PWM9/n24 ,\PWM9/n24 }),
    .b({\PWM9/n25_neg_lutinv ,\PWM9/n25_neg_lutinv }),
    .c(\PWM9/n26 [10:9]),
    .clk(clk100m),
    .d(\PWM9/pnumr [10:9]),
    .mi({\U_AHB/h2h_hwdata [10],1'b1}),
    .sr(\U_AHB/n65 ),
    .f({_al_u2467_o,_al_u2425_o}),
    .q({pnum9[10],pnum9[32]}));  // src/AHB.v(76)
  // src/AHB.v(76)
  // src/AHB.v(76)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg27_b11|U_AHB/reg27_b8  (
    .a({\PWM9/n24 ,\PWM9/n24 }),
    .b({\PWM9/n25_neg_lutinv ,\PWM9/n25_neg_lutinv }),
    .c({\PWM9/n26 [11],\PWM9/n26 [8]}),
    .clk(clk100m),
    .d({\PWM9/pnumr [11],\PWM9/pnumr [8]}),
    .mi({\U_AHB/h2h_hwdata [11],\U_AHB/h2h_hwdata [8]}),
    .sr(\U_AHB/n65 ),
    .f({_al_u2465_o,_al_u2427_o}),
    .q({pnum9[11],pnum9[8]}));  // src/AHB.v(76)
  // src/AHB.v(76)
  // src/AHB.v(76)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg27_b12|U_AHB/reg27_b7  (
    .a({\PWM9/n24 ,\PWM9/n24 }),
    .b({\PWM9/n25_neg_lutinv ,\PWM9/n25_neg_lutinv }),
    .c({\PWM9/n26 [12],\PWM9/n26 [7]}),
    .clk(clk100m),
    .d({\PWM9/pnumr [12],\PWM9/pnumr [7]}),
    .mi({\U_AHB/h2h_hwdata [12],\U_AHB/h2h_hwdata [7]}),
    .sr(\U_AHB/n65 ),
    .f({_al_u2463_o,_al_u2429_o}),
    .q({pnum9[12],pnum9[7]}));  // src/AHB.v(76)
  // src/AHB.v(76)
  // src/AHB.v(76)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg27_b13|U_AHB/reg27_b6  (
    .a({\PWM9/n24 ,\PWM9/n24 }),
    .b({\PWM9/n25_neg_lutinv ,\PWM9/n25_neg_lutinv }),
    .c({\PWM9/n26 [13],\PWM9/n26 [6]}),
    .clk(clk100m),
    .d({\PWM9/pnumr [13],\PWM9/pnumr [6]}),
    .mi({\U_AHB/h2h_hwdata [13],\U_AHB/h2h_hwdata [6]}),
    .sr(\U_AHB/n65 ),
    .f({_al_u2461_o,_al_u2431_o}),
    .q({pnum9[13],pnum9[6]}));  // src/AHB.v(76)
  // src/AHB.v(76)
  // src/AHB.v(76)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg27_b14|U_AHB/reg27_b5  (
    .a({\PWM9/n24 ,\PWM9/n24 }),
    .b({\PWM9/n25_neg_lutinv ,\PWM9/n25_neg_lutinv }),
    .c({\PWM9/n26 [14],\PWM9/n26 [5]}),
    .clk(clk100m),
    .d({\PWM9/pnumr [14],\PWM9/pnumr [5]}),
    .mi({\U_AHB/h2h_hwdata [14],\U_AHB/h2h_hwdata [5]}),
    .sr(\U_AHB/n65 ),
    .f({_al_u2459_o,_al_u2433_o}),
    .q({pnum9[14],pnum9[5]}));  // src/AHB.v(76)
  // src/AHB.v(76)
  // src/AHB.v(76)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg27_b15|U_AHB/reg27_b4  (
    .a({\PWM9/n24 ,\PWM9/n24 }),
    .b({\PWM9/n25_neg_lutinv ,\PWM9/n25_neg_lutinv }),
    .c({\PWM9/n26 [15],\PWM9/n26 [4]}),
    .clk(clk100m),
    .d({\PWM9/pnumr [15],\PWM9/pnumr [4]}),
    .mi({\U_AHB/h2h_hwdata [15],\U_AHB/h2h_hwdata [4]}),
    .sr(\U_AHB/n65 ),
    .f({_al_u2457_o,_al_u2435_o}),
    .q({pnum9[15],pnum9[4]}));  // src/AHB.v(76)
  // src/AHB.v(76)
  // src/AHB.v(76)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg27_b16|U_AHB/reg27_b3  (
    .a({\PWM9/n24 ,\PWM9/n24 }),
    .b({\PWM9/n25_neg_lutinv ,\PWM9/n25_neg_lutinv }),
    .c({\PWM9/n26 [16],\PWM9/n26 [3]}),
    .clk(clk100m),
    .d({\PWM9/pnumr [16],\PWM9/pnumr [3]}),
    .mi({\U_AHB/h2h_hwdata [16],\U_AHB/h2h_hwdata [3]}),
    .sr(\U_AHB/n65 ),
    .f({_al_u2455_o,_al_u2437_o}),
    .q({pnum9[16],pnum9[3]}));  // src/AHB.v(76)
  // src/AHB.v(76)
  // src/AHB.v(76)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg27_b17|U_AHB/reg27_b23  (
    .a({\PWM9/n24 ,\PWM9/n24 }),
    .b({\PWM9/n25_neg_lutinv ,\PWM9/n25_neg_lutinv }),
    .c({\PWM9/n26 [17],\PWM9/n26 [23]}),
    .clk(clk100m),
    .d({\PWM9/pnumr [17],\PWM9/pnumr [23]}),
    .mi({\U_AHB/h2h_hwdata [17],\U_AHB/h2h_hwdata [23]}),
    .sr(\U_AHB/n65 ),
    .f({_al_u2453_o,_al_u2439_o}),
    .q({pnum9[17],pnum9[23]}));  // src/AHB.v(76)
  // src/AHB.v(76)
  // src/AHB.v(76)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg27_b18|U_AHB/reg27_b22  (
    .a({\PWM9/n24 ,\PWM9/n24 }),
    .b({\PWM9/n25_neg_lutinv ,\PWM9/n25_neg_lutinv }),
    .c({\PWM9/n26 [18],\PWM9/n26 [22]}),
    .clk(clk100m),
    .d({\PWM9/pnumr [18],\PWM9/pnumr [22]}),
    .mi({\U_AHB/h2h_hwdata [18],\U_AHB/h2h_hwdata [22]}),
    .sr(\U_AHB/n65 ),
    .f({_al_u2451_o,_al_u2441_o}),
    .q({pnum9[18],pnum9[22]}));  // src/AHB.v(76)
  // src/AHB.v(76)
  // src/AHB.v(76)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg27_b19|U_AHB/reg27_b21  (
    .a({\PWM9/n24 ,\PWM9/n24 }),
    .b({\PWM9/n25_neg_lutinv ,\PWM9/n25_neg_lutinv }),
    .c({\PWM9/n26 [19],\PWM9/n26 [21]}),
    .clk(clk100m),
    .d({\PWM9/pnumr [19],\PWM9/pnumr [21]}),
    .mi({\U_AHB/h2h_hwdata [19],\U_AHB/h2h_hwdata [21]}),
    .sr(\U_AHB/n65 ),
    .f({_al_u2449_o,_al_u2443_o}),
    .q({pnum9[19],pnum9[21]}));  // src/AHB.v(76)
  // src/AHB.v(76)
  // src/AHB.v(76)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg27_b1|U_AHB/reg27_b20  (
    .a({\PWM9/n24 ,\PWM9/n24 }),
    .b({\PWM9/n25_neg_lutinv ,\PWM9/n25_neg_lutinv }),
    .c({\PWM9/n26 [1],\PWM9/n26 [20]}),
    .clk(clk100m),
    .d({\PWM9/pnumr [1],\PWM9/pnumr [20]}),
    .mi({\U_AHB/h2h_hwdata [1],\U_AHB/h2h_hwdata [20]}),
    .sr(\U_AHB/n65 ),
    .f({_al_u2469_o,_al_u2445_o}),
    .q({pnum9[1],pnum9[20]}));  // src/AHB.v(76)
  // src/AHB.v(76)
  // src/AHB.v(76)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(D*~(C*B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b0111111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg27_b24|U_AHB/reg27_b2  (
    .a({_al_u2880_o,\PWM9/n24 }),
    .b({_al_u2888_o,\PWM9/n25_neg_lutinv }),
    .c({_al_u2896_o,\PWM9/n26 [2]}),
    .clk(clk100m),
    .d({pwm_state_read[14],\PWM9/pnumr [2]}),
    .mi({\U_AHB/h2h_hwdata [24],\U_AHB/h2h_hwdata [2]}),
    .sr(\U_AHB/n65 ),
    .f({\PWME/u14_sel_is_1_o ,_al_u2447_o}),
    .q({pnum9[24],pnum9[2]}));  // src/AHB.v(76)
  // src/AHB.v(76)
  // src/AHB.v(76)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg27_b27|U_AHB/reg27_b25  (
    .c({pwm_state_read[13],pwm_state_read[13]}),
    .clk(clk100m),
    .d({_al_u2817_o,\PWMD/n0_lutinv }),
    .mi({\U_AHB/h2h_hwdata [27],\U_AHB/h2h_hwdata [25]}),
    .sr(\U_AHB/n65 ),
    .f({\PWMD/u14_sel_is_1_o ,\PWMD/n24 }),
    .q({pnum9[27],pnum9[25]}));  // src/AHB.v(76)
  // src/AHB.v(76)
  // src/AHB.v(76)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(D*~(C*B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0111111100000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg27_b28|U_AHB/reg27_b9  (
    .a({_al_u2723_o,open_n30599}),
    .b({_al_u2731_o,open_n30600}),
    .c({_al_u2737_o,pwm_state_read[9]}),
    .clk(clk100m),
    .d({pwm_state_read[12],_al_u2497_o}),
    .mi({\U_AHB/h2h_hwdata [28],\U_AHB/h2h_hwdata [9]}),
    .sr(\U_AHB/n65 ),
    .f({\PWMC/u14_sel_is_1_o ,\PWM9/u14_sel_is_1_o }),
    .q({pnum9[28],pnum9[9]}));  // src/AHB.v(76)
  // src/AHB.v(77)
  // src/AHB.v(77)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~(D*C*B*A))"),
    //.LUTF1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("(~1*~(D*C*B*A))"),
    //.LUTG1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111111111111111),
    .INIT_LUTF1(16'b1010100000100000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1010100000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg28_b0|U_AHB/reg28_b24  (
    .a({\PWMA/n24 ,_al_u2340_o}),
    .b({\PWMA/n25_neg_lutinv ,_al_u2342_o}),
    .c({\PWMA/n26 [0],_al_u2343_o}),
    .clk(clk100m),
    .d({\PWMA/pnumr [0],pnumcnt8[0]}),
    .e({open_n30616,\PWM8/stopreq }),
    .mi({\U_AHB/h2h_hwdata [0],\U_AHB/h2h_hwdata [24]}),
    .sr(\U_AHB/n67 ),
    .f({_al_u2553_o,_al_u3031_o}),
    .q({pnumA[0],pnumA[24]}));  // src/AHB.v(77)
  // src/AHB.v(77)
  // src/AHB.v(77)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~(D*C*B*A))"),
    //.LUTF1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("(~1*~(D*C*B*A))"),
    //.LUTG1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111111111111111),
    .INIT_LUTF1(16'b1010100000100000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1010100000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg28_b10|U_AHB/reg28_b28  (
    .a({\PWMA/n24 ,_al_u2178_o}),
    .b({\PWMA/n25_neg_lutinv ,_al_u2180_o}),
    .c({\PWMA/n26 [10],_al_u2181_o}),
    .clk(clk100m),
    .d({\PWMA/pnumr [10],pnumcnt6[0]}),
    .e({open_n30633,\PWM6/stopreq }),
    .mi({\U_AHB/h2h_hwdata [10],\U_AHB/h2h_hwdata [28]}),
    .sr(\U_AHB/n67 ),
    .f({_al_u2549_o,_al_u3025_o}),
    .q({pnumA[10],pnumA[28]}));  // src/AHB.v(77)
  // src/AHB.v(77)
  // src/AHB.v(77)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg28_b11|U_AHB/reg28_b32  (
    .a({\PWMA/n24 ,\PWMA/n24 }),
    .b({\PWMA/n25_neg_lutinv ,\PWMA/n25_neg_lutinv }),
    .c({\PWMA/n26 [11],\PWMA/n26 [9]}),
    .clk(clk100m),
    .d({\PWMA/pnumr [11],\PWMA/pnumr [9]}),
    .mi({\U_AHB/h2h_hwdata [11],1'b1}),
    .sr(\U_AHB/n67 ),
    .f({_al_u2547_o,_al_u2507_o}),
    .q({pnumA[11],pnumA[32]}));  // src/AHB.v(77)
  // src/AHB.v(77)
  // src/AHB.v(77)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg28_b12|U_AHB/reg28_b8  (
    .a({\PWMA/n24 ,\PWMA/n24 }),
    .b({\PWMA/n25_neg_lutinv ,\PWMA/n25_neg_lutinv }),
    .c({\PWMA/n26 [12],\PWMA/n26 [8]}),
    .clk(clk100m),
    .d({\PWMA/pnumr [12],\PWMA/pnumr [8]}),
    .mi({\U_AHB/h2h_hwdata [12],\U_AHB/h2h_hwdata [8]}),
    .sr(\U_AHB/n67 ),
    .f({_al_u2545_o,_al_u2509_o}),
    .q({pnumA[12],pnumA[8]}));  // src/AHB.v(77)
  // src/AHB.v(77)
  // src/AHB.v(77)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg28_b13|U_AHB/reg28_b7  (
    .a({\PWMA/n24 ,\PWMA/n24 }),
    .b({\PWMA/n25_neg_lutinv ,\PWMA/n25_neg_lutinv }),
    .c({\PWMA/n26 [13],\PWMA/n26 [7]}),
    .clk(clk100m),
    .d({\PWMA/pnumr [13],\PWMA/pnumr [7]}),
    .mi({\U_AHB/h2h_hwdata [13],\U_AHB/h2h_hwdata [7]}),
    .sr(\U_AHB/n67 ),
    .f({_al_u2543_o,_al_u2511_o}),
    .q({pnumA[13],pnumA[7]}));  // src/AHB.v(77)
  // src/AHB.v(77)
  // src/AHB.v(77)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg28_b14|U_AHB/reg28_b6  (
    .a({\PWMA/n24 ,\PWMA/n24 }),
    .b({\PWMA/n25_neg_lutinv ,\PWMA/n25_neg_lutinv }),
    .c({\PWMA/n26 [14],\PWMA/n26 [6]}),
    .clk(clk100m),
    .d({\PWMA/pnumr [14],\PWMA/pnumr [6]}),
    .mi({\U_AHB/h2h_hwdata [14],\U_AHB/h2h_hwdata [6]}),
    .sr(\U_AHB/n67 ),
    .f({_al_u2541_o,_al_u2513_o}),
    .q({pnumA[14],pnumA[6]}));  // src/AHB.v(77)
  // src/AHB.v(77)
  // src/AHB.v(77)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg28_b15|U_AHB/reg28_b5  (
    .a({\PWMA/n24 ,\PWMA/n24 }),
    .b({\PWMA/n25_neg_lutinv ,\PWMA/n25_neg_lutinv }),
    .c({\PWMA/n26 [15],\PWMA/n26 [5]}),
    .clk(clk100m),
    .d({\PWMA/pnumr [15],\PWMA/pnumr [5]}),
    .mi({\U_AHB/h2h_hwdata [15],\U_AHB/h2h_hwdata [5]}),
    .sr(\U_AHB/n67 ),
    .f({_al_u2539_o,_al_u2515_o}),
    .q({pnumA[15],pnumA[5]}));  // src/AHB.v(77)
  // src/AHB.v(77)
  // src/AHB.v(77)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg28_b16|U_AHB/reg28_b4  (
    .a({\PWMA/n24 ,\PWMA/n24 }),
    .b({\PWMA/n25_neg_lutinv ,\PWMA/n25_neg_lutinv }),
    .c({\PWMA/n26 [16],\PWMA/n26 [4]}),
    .clk(clk100m),
    .d({\PWMA/pnumr [16],\PWMA/pnumr [4]}),
    .mi({\U_AHB/h2h_hwdata [16],\U_AHB/h2h_hwdata [4]}),
    .sr(\U_AHB/n67 ),
    .f({_al_u2537_o,_al_u2517_o}),
    .q({pnumA[16],pnumA[4]}));  // src/AHB.v(77)
  // src/AHB.v(77)
  // src/AHB.v(77)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg28_b17|U_AHB/reg28_b3  (
    .a({\PWMA/n24 ,\PWMA/n24 }),
    .b({\PWMA/n25_neg_lutinv ,\PWMA/n25_neg_lutinv }),
    .c({\PWMA/n26 [17],\PWMA/n26 [3]}),
    .clk(clk100m),
    .d({\PWMA/pnumr [17],\PWMA/pnumr [3]}),
    .mi({\U_AHB/h2h_hwdata [17],\U_AHB/h2h_hwdata [3]}),
    .sr(\U_AHB/n67 ),
    .f({_al_u2535_o,_al_u2519_o}),
    .q({pnumA[17],pnumA[3]}));  // src/AHB.v(77)
  // src/AHB.v(77)
  // src/AHB.v(77)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg28_b18|U_AHB/reg28_b23  (
    .a({\PWMA/n24 ,\PWMA/n24 }),
    .b({\PWMA/n25_neg_lutinv ,\PWMA/n25_neg_lutinv }),
    .c({\PWMA/n26 [18],\PWMA/n26 [23]}),
    .clk(clk100m),
    .d({\PWMA/pnumr [18],\PWMA/pnumr [23]}),
    .mi({\U_AHB/h2h_hwdata [18],\U_AHB/h2h_hwdata [23]}),
    .sr(\U_AHB/n67 ),
    .f({_al_u2533_o,_al_u2521_o}),
    .q({pnumA[18],pnumA[23]}));  // src/AHB.v(77)
  // src/AHB.v(77)
  // src/AHB.v(77)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg28_b19|U_AHB/reg28_b22  (
    .a({\PWMA/n24 ,\PWMA/n24 }),
    .b({\PWMA/n25_neg_lutinv ,\PWMA/n25_neg_lutinv }),
    .c({\PWMA/n26 [19],\PWMA/n26 [22]}),
    .clk(clk100m),
    .d({\PWMA/pnumr [19],\PWMA/pnumr [22]}),
    .mi({\U_AHB/h2h_hwdata [19],\U_AHB/h2h_hwdata [22]}),
    .sr(\U_AHB/n67 ),
    .f({_al_u2531_o,_al_u2523_o}),
    .q({pnumA[19],pnumA[22]}));  // src/AHB.v(77)
  // src/AHB.v(77)
  // src/AHB.v(77)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg28_b1|U_AHB/reg28_b21  (
    .a({\PWMA/n24 ,\PWMA/n24 }),
    .b({\PWMA/n25_neg_lutinv ,\PWMA/n25_neg_lutinv }),
    .c({\PWMA/n26 [1],\PWMA/n26 [21]}),
    .clk(clk100m),
    .d({\PWMA/pnumr [1],\PWMA/pnumr [21]}),
    .mi({\U_AHB/h2h_hwdata [1],\U_AHB/h2h_hwdata [21]}),
    .sr(\U_AHB/n67 ),
    .f({_al_u2551_o,_al_u2525_o}),
    .q({pnumA[1],pnumA[21]}));  // src/AHB.v(77)
  // src/AHB.v(77)
  // src/AHB.v(77)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg28_b27|U_AHB/reg28_b25  (
    .c({pwm_state_read[7],pwm_state_read[8]}),
    .clk(clk100m),
    .d({_al_u2335_o,_al_u2415_o}),
    .mi({\U_AHB/h2h_hwdata [27],\U_AHB/h2h_hwdata [25]}),
    .sr(\U_AHB/n67 ),
    .f({\PWM7/u14_sel_is_1_o ,\PWM8/u14_sel_is_1_o }),
    .q({pnumA[27],pnumA[25]}));  // src/AHB.v(77)
  // src/AHB.v(77)
  // src/AHB.v(77)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg28_b2|U_AHB/reg28_b20  (
    .a({\PWMA/n24 ,\PWMA/n24 }),
    .b({\PWMA/n25_neg_lutinv ,\PWMA/n25_neg_lutinv }),
    .c({\PWMA/n26 [2],\PWMA/n26 [20]}),
    .clk(clk100m),
    .d({\PWMA/pnumr [2],\PWMA/pnumr [20]}),
    .mi({\U_AHB/h2h_hwdata [2],\U_AHB/h2h_hwdata [20]}),
    .sr(\U_AHB/n67 ),
    .f({_al_u2529_o,_al_u2527_o}),
    .q({pnumA[2],pnumA[20]}));  // src/AHB.v(77)
  // src/AHB.v(77)
  // src/AHB.v(77)
  EF2_PHY_MSLICE #(
    //.LUT0("(D*~(C*B*A))"),
    //.LUT1("(C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111111100000000),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg28_b31|U_AHB/reg28_b29  (
    .a({open_n30821,_al_u2238_o}),
    .b({open_n30822,_al_u2247_o}),
    .c({pwm_state_read[5],_al_u2253_o}),
    .clk(clk100m),
    .d({_al_u2173_o,pwm_state_read[6]}),
    .mi({\U_AHB/h2h_hwdata [31],\U_AHB/h2h_hwdata [29]}),
    .sr(\U_AHB/n67 ),
    .f({\PWM5/u14_sel_is_1_o ,\PWM6/u14_sel_is_1_o }),
    .q({pnumA[31],pnumA[29]}));  // src/AHB.v(77)
  // src/AHB.v(78)
  // src/AHB.v(78)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg29_b0|U_AHB/reg29_b32  (
    .a({\PWMB/n24 ,\PWMB/n24 }),
    .b({\PWMB/n25_neg_lutinv ,\PWMB/n25_neg_lutinv }),
    .c({\PWMB/n26 [0],\PWMB/n26 [9]}),
    .clk(clk100m),
    .d({\PWMB/pnumr [0],\PWMB/pnumr [9]}),
    .mi({\U_AHB/h2h_hwdata [0],1'b1}),
    .sr(\U_AHB/n69 ),
    .f({_al_u2632_o,_al_u2586_o}),
    .q({pnumB[0],pnumB[32]}));  // src/AHB.v(78)
  // src/AHB.v(78)
  // src/AHB.v(78)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg29_b10|U_AHB/reg29_b8  (
    .a({\PWMB/n24 ,\PWMB/n24 }),
    .b({\PWMB/n25_neg_lutinv ,\PWMB/n25_neg_lutinv }),
    .c({\PWMB/n26 [10],\PWMB/n26 [8]}),
    .clk(clk100m),
    .d({\PWMB/pnumr [10],\PWMB/pnumr [8]}),
    .mi({\U_AHB/h2h_hwdata [10],\U_AHB/h2h_hwdata [8]}),
    .sr(\U_AHB/n69 ),
    .f({_al_u2628_o,_al_u2588_o}),
    .q({pnumB[10],pnumB[8]}));  // src/AHB.v(78)
  // src/AHB.v(78)
  // src/AHB.v(78)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg29_b11|U_AHB/reg29_b7  (
    .a({\PWMB/n24 ,\PWMB/n24 }),
    .b({\PWMB/n25_neg_lutinv ,\PWMB/n25_neg_lutinv }),
    .c({\PWMB/n26 [11],\PWMB/n26 [7]}),
    .clk(clk100m),
    .d({\PWMB/pnumr [11],\PWMB/pnumr [7]}),
    .mi({\U_AHB/h2h_hwdata [11],\U_AHB/h2h_hwdata [7]}),
    .sr(\U_AHB/n69 ),
    .f({_al_u2626_o,_al_u2590_o}),
    .q({pnumB[11],pnumB[7]}));  // src/AHB.v(78)
  // src/AHB.v(78)
  // src/AHB.v(78)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg29_b12|U_AHB/reg29_b6  (
    .a({\PWMB/n24 ,\PWMB/n24 }),
    .b({\PWMB/n25_neg_lutinv ,\PWMB/n25_neg_lutinv }),
    .c({\PWMB/n26 [12],\PWMB/n26 [6]}),
    .clk(clk100m),
    .d({\PWMB/pnumr [12],\PWMB/pnumr [6]}),
    .mi({\U_AHB/h2h_hwdata [12],\U_AHB/h2h_hwdata [6]}),
    .sr(\U_AHB/n69 ),
    .f({_al_u2624_o,_al_u2592_o}),
    .q({pnumB[12],pnumB[6]}));  // src/AHB.v(78)
  // src/AHB.v(78)
  // src/AHB.v(78)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg29_b13|U_AHB/reg29_b5  (
    .a({\PWMB/n24 ,\PWMB/n24 }),
    .b({\PWMB/n25_neg_lutinv ,\PWMB/n25_neg_lutinv }),
    .c({\PWMB/n26 [13],\PWMB/n26 [5]}),
    .clk(clk100m),
    .d({\PWMB/pnumr [13],\PWMB/pnumr [5]}),
    .mi({\U_AHB/h2h_hwdata [13],\U_AHB/h2h_hwdata [5]}),
    .sr(\U_AHB/n69 ),
    .f({_al_u2622_o,_al_u2594_o}),
    .q({pnumB[13],pnumB[5]}));  // src/AHB.v(78)
  // src/AHB.v(78)
  // src/AHB.v(78)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg29_b14|U_AHB/reg29_b4  (
    .a({\PWMB/n24 ,\PWMB/n24 }),
    .b({\PWMB/n25_neg_lutinv ,\PWMB/n25_neg_lutinv }),
    .c({\PWMB/n26 [14],\PWMB/n26 [4]}),
    .clk(clk100m),
    .d({\PWMB/pnumr [14],\PWMB/pnumr [4]}),
    .mi({\U_AHB/h2h_hwdata [14],\U_AHB/h2h_hwdata [4]}),
    .sr(\U_AHB/n69 ),
    .f({_al_u2620_o,_al_u2596_o}),
    .q({pnumB[14],pnumB[4]}));  // src/AHB.v(78)
  // src/AHB.v(78)
  // src/AHB.v(78)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg29_b15|U_AHB/reg29_b3  (
    .a({\PWMB/n24 ,\PWMB/n24 }),
    .b({\PWMB/n25_neg_lutinv ,\PWMB/n25_neg_lutinv }),
    .c({\PWMB/n26 [15],\PWMB/n26 [3]}),
    .clk(clk100m),
    .d({\PWMB/pnumr [15],\PWMB/pnumr [3]}),
    .mi({\U_AHB/h2h_hwdata [15],\U_AHB/h2h_hwdata [3]}),
    .sr(\U_AHB/n69 ),
    .f({_al_u2618_o,_al_u2598_o}),
    .q({pnumB[15],pnumB[3]}));  // src/AHB.v(78)
  // src/AHB.v(78)
  // src/AHB.v(78)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg29_b16|U_AHB/reg29_b23  (
    .a({\PWMB/n24 ,\PWMB/n24 }),
    .b({\PWMB/n25_neg_lutinv ,\PWMB/n25_neg_lutinv }),
    .c({\PWMB/n26 [16],\PWMB/n26 [23]}),
    .clk(clk100m),
    .d({\PWMB/pnumr [16],\PWMB/pnumr [23]}),
    .mi({\U_AHB/h2h_hwdata [16],\U_AHB/h2h_hwdata [23]}),
    .sr(\U_AHB/n69 ),
    .f({_al_u2616_o,_al_u2600_o}),
    .q({pnumB[16],pnumB[23]}));  // src/AHB.v(78)
  // src/AHB.v(78)
  // src/AHB.v(78)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg29_b17|U_AHB/reg29_b22  (
    .a({\PWMB/n24 ,\PWMB/n24 }),
    .b({\PWMB/n25_neg_lutinv ,\PWMB/n25_neg_lutinv }),
    .c({\PWMB/n26 [17],\PWMB/n26 [22]}),
    .clk(clk100m),
    .d({\PWMB/pnumr [17],\PWMB/pnumr [22]}),
    .mi({\U_AHB/h2h_hwdata [17],\U_AHB/h2h_hwdata [22]}),
    .sr(\U_AHB/n69 ),
    .f({_al_u2614_o,_al_u2602_o}),
    .q({pnumB[17],pnumB[22]}));  // src/AHB.v(78)
  // src/AHB.v(78)
  // src/AHB.v(78)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg29_b18|U_AHB/reg29_b21  (
    .a({\PWMB/n24 ,\PWMB/n24 }),
    .b({\PWMB/n25_neg_lutinv ,\PWMB/n25_neg_lutinv }),
    .c({\PWMB/n26 [18],\PWMB/n26 [21]}),
    .clk(clk100m),
    .d({\PWMB/pnumr [18],\PWMB/pnumr [21]}),
    .mi({\U_AHB/h2h_hwdata [18],\U_AHB/h2h_hwdata [21]}),
    .sr(\U_AHB/n69 ),
    .f({_al_u2612_o,_al_u2604_o}),
    .q({pnumB[18],pnumB[21]}));  // src/AHB.v(78)
  // src/AHB.v(78)
  // src/AHB.v(78)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg29_b19|U_AHB/reg29_b20  (
    .a({\PWMB/n24 ,\PWMB/n24 }),
    .b({\PWMB/n25_neg_lutinv ,\PWMB/n25_neg_lutinv }),
    .c({\PWMB/n26 [19],\PWMB/n26 [20]}),
    .clk(clk100m),
    .d({\PWMB/pnumr [19],\PWMB/pnumr [20]}),
    .mi({\U_AHB/h2h_hwdata [19],\U_AHB/h2h_hwdata [20]}),
    .sr(\U_AHB/n69 ),
    .f({_al_u2610_o,_al_u2606_o}),
    .q({pnumB[19],pnumB[20]}));  // src/AHB.v(78)
  // src/AHB.v(78)
  // src/AHB.v(78)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg29_b1|U_AHB/reg29_b2  (
    .a({\PWMB/n24 ,\PWMB/n24 }),
    .b({\PWMB/n25_neg_lutinv ,\PWMB/n25_neg_lutinv }),
    .c({\PWMB/n26 [1],\PWMB/n26 [2]}),
    .clk(clk100m),
    .d({\PWMB/pnumr [1],\PWMB/pnumr [2]}),
    .mi({\U_AHB/h2h_hwdata [1],\U_AHB/h2h_hwdata [2]}),
    .sr(\U_AHB/n69 ),
    .f({_al_u2630_o,_al_u2608_o}),
    .q({pnumB[1],pnumB[2]}));  // src/AHB.v(78)
  // src/AHB.v(78)
  // src/AHB.v(78)
  EF2_PHY_LSLICE #(
    //.LUTF0("(D*C*B*A)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(D*C*B*A)"),
    //.LUTG1("(C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000000000000000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg29_b24|U_AHB/reg29_b9  (
    .a({open_n31005,_al_u1647_o}),
    .b({open_n31006,_al_u1642_o}),
    .c({pwm_state_read[4],_al_u2986_o}),
    .clk(clk100m),
    .d({_al_u2091_o,_al_u2987_o}),
    .mi({\U_AHB/h2h_hwdata [24],\U_AHB/h2h_hwdata [9]}),
    .sr(\U_AHB/n69 ),
    .f({\PWM4/u14_sel_is_1_o ,_al_u2988_o}),
    .q({pnumB[24],pnumB[9]}));  // src/AHB.v(78)
  // src/AHB.v(78)
  // src/AHB.v(78)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(D*~(C*B*A))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(D*~(C*B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0111111100000000),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0111111100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg29_b29|U_AHB/reg29_b28  (
    .a({_al_u1912_o,_al_u3239_o}),
    .b({_al_u1919_o,\U_AHB/n96 }),
    .c({_al_u1927_o,\U_AHB/n93 }),
    .clk(clk100m),
    .d({pwm_state_read[2],pnumcntF[18]}),
    .e({open_n31026,pwm_state_read[2]}),
    .mi(\U_AHB/h2h_hwdata [29:28]),
    .sr(\U_AHB/n69 ),
    .f({\PWM2/u14_sel_is_1_o ,_al_u3240_o}),
    .q(pnumB[29:28]));  // src/AHB.v(78)
  // src/AHB.v(78)
  // src/AHB.v(78)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg29_b30|U_AHB/reg29_b31  (
    .c(pwm_state_read[1:0]),
    .clk(clk100m),
    .d({_al_u1847_o,_al_u1765_o}),
    .mi({\U_AHB/h2h_hwdata [30],\U_AHB/h2h_hwdata [31]}),
    .sr(\U_AHB/n69 ),
    .f({\PWM1/u14_sel_is_1_o ,\PWM0/u14_sel_is_1_o }),
    .q({pnumB[30],pnumB[31]}));  // src/AHB.v(78)
  // src/AHB.v(47)
  // src/AHB.v(47)
  EF2_PHY_MSLICE #(
    //.LUT0("(D*~C*B*A)"),
    //.LUT1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000100000000000),
    .INIT_LUT1(16'b1000010000100001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg2_b10|U_AHB/reg2_b0  (
    .a({\PWM1/FreCnt [0],\U_AHB/h2h_hwrite }),
    .b({\PWM1/FreCnt [10],\U_AHB/h2h_haddr [13]}),
    .c({\PWM1/FreCntr [0],\U_AHB/h2h_haddr [14]}),
    .ce(\U_AHB/n4 ),
    .clk(clk100m),
    .d({\PWM1/FreCntr [10],\U_AHB/h2h_haddr [6]}),
    .mi({\U_AHB/h2h_hwdata [10],\U_AHB/h2h_hwdata [0]}),
    .f({_al_u1384_o,\U_AHB/n4 }),
    .q({freq1[10],freq1[0]}));  // src/AHB.v(47)
  // src/AHB.v(47)
  // src/AHB.v(47)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*~C)*~(~D*B))"),
    //.LUTF1("(~(~D*B)*~(~C*A))"),
    //.LUTG0("(A*~(1*~C)*~(~D*B))"),
    //.LUTG1("(~(~D*B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101000100010),
    .INIT_LUTF1(16'b1111010100110001),
    .INIT_LUTG0(16'b1010000000100000),
    .INIT_LUTG1(16'b1111010100110001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg2_b11|U_AHB/reg2_b2  (
    .a({\PWM1/FreCnt [10],_al_u1823_o}),
    .b({\PWM1/FreCnt [17],\PWM1/FreCnt [1]}),
    .c({\PWM1/FreCntr [11],\PWM1/FreCnt [23]}),
    .ce(\U_AHB/n4 ),
    .clk(clk100m),
    .d({\PWM1/FreCntr [18],\PWM1/FreCntr [2]}),
    .e({open_n31078,\PWM1/FreCntr [24]}),
    .mi({\U_AHB/h2h_hwdata [11],\U_AHB/h2h_hwdata [2]}),
    .f({_al_u1823_o,_al_u1824_o}),
    .q({freq1[11],freq1[2]}));  // src/AHB.v(47)
  // src/AHB.v(47)
  // src/AHB.v(47)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~(~D*B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111010100110001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg2_b12|U_AHB/reg2_b15  (
    .a({\PWM1/FreCnt [12],open_n31095}),
    .b({\PWM1/FreCnt [15],open_n31096}),
    .c({\PWM1/FreCntr [12],pwm_state_read[1]}),
    .ce(\U_AHB/n4 ),
    .clk(clk100m),
    .d({\PWM1/FreCntr [15],\PWM1/n0_lutinv }),
    .mi({\U_AHB/h2h_hwdata [12],\U_AHB/h2h_hwdata [15]}),
    .f({_al_u1385_o,\PWM1/n24 }),
    .q({freq1[12],freq1[15]}));  // src/AHB.v(47)
  // src/AHB.v(47)
  // src/AHB.v(47)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg2_b13|U_AHB/reg2_b19  (
    .a({\PWM1/FreCnt [13],_al_u1392_o}),
    .b({\PWM1/FreCnt [16],\PWM1/FreCnt [19]}),
    .c({\PWM1/FreCntr [13],\PWM1/FreCnt [2]}),
    .ce(\U_AHB/n4 ),
    .clk(clk100m),
    .d({\PWM1/FreCntr [16],\PWM1/FreCntr [19]}),
    .e({open_n31111,\PWM1/FreCntr [2]}),
    .mi({\U_AHB/h2h_hwdata [13],\U_AHB/h2h_hwdata [19]}),
    .f({_al_u1392_o,_al_u1393_o}),
    .q({freq1[13],freq1[19]}));  // src/AHB.v(47)
  // src/AHB.v(47)
  // src/AHB.v(47)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg2_b14|U_AHB/reg2_b20  (
    .a({\PWM1/FreCnt [14],_al_u1390_o}),
    .b({\PWM1/FreCnt [25],\PWM1/FreCnt [20]}),
    .c({\PWM1/FreCntr [14],\PWM1/FreCnt [26]}),
    .ce(\U_AHB/n4 ),
    .clk(clk100m),
    .d({\PWM1/FreCntr [25],\PWM1/FreCntr [20]}),
    .e({open_n31128,\PWM1/FreCntr [26]}),
    .mi({\U_AHB/h2h_hwdata [14],\U_AHB/h2h_hwdata [20]}),
    .f({_al_u1390_o,_al_u1391_o}),
    .q({freq1[14],freq1[20]}));  // src/AHB.v(47)
  // src/AHB.v(47)
  // src/AHB.v(47)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg2_b17|U_AHB/reg2_b24  (
    .a({\PWM1/FreCnt [17],_al_u1380_o}),
    .b({\PWM1/FreCnt [8],\PWM1/FreCnt [11]}),
    .c({\PWM1/FreCntr [17],\PWM1/FreCnt [24]}),
    .ce(\U_AHB/n4 ),
    .clk(clk100m),
    .d({\PWM1/FreCntr [8],\PWM1/FreCntr [11]}),
    .e({open_n31145,\PWM1/FreCntr [24]}),
    .mi({\U_AHB/h2h_hwdata [17],\U_AHB/h2h_hwdata [24]}),
    .f({_al_u1380_o,_al_u1381_o}),
    .q({freq1[17],freq1[24]}));  // src/AHB.v(47)
  // src/AHB.v(47)
  // src/AHB.v(47)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg2_b18|U_AHB/reg2_b16  (
    .a({\PWM1/FreCnt [16],open_n31162}),
    .b({\PWM1/FreCnt [17],limit_r_pad[1]}),
    .c({\PWM1/FreCnt [18],limit_l_pad[1]}),
    .ce(\U_AHB/n4 ),
    .clk(clk100m),
    .d({\PWM1/FreCnt [19],\PWM1/n11 }),
    .mi({\U_AHB/h2h_hwdata [18],\U_AHB/h2h_hwdata [16]}),
    .f({_al_u776_o,_al_u3011_o}),
    .q({freq1[18],freq1[16]}));  // src/AHB.v(47)
  // src/AHB.v(47)
  // src/AHB.v(47)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*B*A*~(0@D))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(C*B*A*~(1@D))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg2_b1|U_AHB/reg2_b6  (
    .a({\PWM1/FreCnt [1],_al_u1386_o}),
    .b({\PWM1/FreCnt [3],_al_u1387_o}),
    .c({\PWM1/FreCntr [1],_al_u1388_o}),
    .ce(\U_AHB/n4 ),
    .clk(clk100m),
    .d({\PWM1/FreCntr [3],\PWM1/FreCnt [6]}),
    .e({open_n31181,\PWM1/FreCntr [6]}),
    .mi({\U_AHB/h2h_hwdata [1],\U_AHB/h2h_hwdata [6]}),
    .f({_al_u1388_o,_al_u1389_o}),
    .q({freq1[1],freq1[6]}));  // src/AHB.v(47)
  // src/AHB.v(47)
  // src/AHB.v(47)
  EF2_PHY_MSLICE #(
    //.LUT0("(~D*~C*~B*A)"),
    //.LUT1("(B*A*~(D@C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000010),
    .INIT_LUT1(16'b1000000000001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg2_b21|U_AHB/reg2_b7  (
    .a({_al_u1384_o,_al_u772_o}),
    .b({_al_u1385_o,\PWM1/FreCnt [7]}),
    .c({\PWM1/FreCnt [21],\PWM1/FreCnt [8]}),
    .ce(\U_AHB/n4 ),
    .clk(clk100m),
    .d({\PWM1/FreCntr [21],\PWM1/FreCnt [9]}),
    .mi({\U_AHB/h2h_hwdata [21],\U_AHB/h2h_hwdata [7]}),
    .f({_al_u1386_o,_al_u773_o}),
    .q({freq1[21],freq1[7]}));  // src/AHB.v(47)
  // src/AHB.v(47)
  // src/AHB.v(47)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg2_b23|U_AHB/reg2_b3  (
    .a({\PWM1/FreCnt [23],_al_u771_o}),
    .b({\PWM1/FreCnt [24],\PWM1/FreCnt [3]}),
    .c({\PWM1/FreCnt [25],\PWM1/FreCnt [4]}),
    .ce(\U_AHB/n4 ),
    .clk(clk100m),
    .d({\PWM1/FreCnt [26],\PWM1/FreCnt [5]}),
    .e({open_n31212,\PWM1/FreCnt [6]}),
    .mi({\U_AHB/h2h_hwdata [23],\U_AHB/h2h_hwdata [3]}),
    .f({_al_u771_o,_al_u772_o}),
    .q({freq1[23],freq1[3]}));  // src/AHB.v(47)
  // src/AHB.v(79)
  // src/AHB.v(79)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*~A)"),
    //.LUTF1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("(~1*~D*~C*~B*~A)"),
    //.LUTG1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000001),
    .INIT_LUTF1(16'b1010100000100000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1010100000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg30_b0|U_AHB/reg30_b30  (
    .a({\PWMC/n24 ,timer[28]}),
    .b({\PWMC/n25_neg_lutinv ,timer[29]}),
    .c({\PWMC/n26 [0],timer[30]}),
    .clk(clk100m),
    .d({\PWMC/pnumr [0],timer[31]}),
    .e({open_n31230,timer[9]}),
    .mi({\U_AHB/h2h_hwdata [0],\U_AHB/h2h_hwdata [30]}),
    .sr(\U_AHB/n71 ),
    .f({_al_u2714_o,_al_u1638_o}),
    .q({pnumC[0],pnumC[30]}));  // src/AHB.v(79)
  // src/AHB.v(79)
  // src/AHB.v(79)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg30_b10|U_AHB/reg30_b32  (
    .a({\PWMC/n24 ,\PWMC/n24 }),
    .b({\PWMC/n25_neg_lutinv ,\PWMC/n25_neg_lutinv }),
    .c(\PWMC/n26 [10:9]),
    .clk(clk100m),
    .d(\PWMC/pnumr [10:9]),
    .mi({\U_AHB/h2h_hwdata [10],1'b1}),
    .sr(\U_AHB/n71 ),
    .f({_al_u2710_o,_al_u2668_o}),
    .q({pnumC[10],pnumC[32]}));  // src/AHB.v(79)
  // src/AHB.v(79)
  // src/AHB.v(79)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg30_b11|U_AHB/reg30_b8  (
    .a({\PWMC/n24 ,\PWMC/n24 }),
    .b({\PWMC/n25_neg_lutinv ,\PWMC/n25_neg_lutinv }),
    .c({\PWMC/n26 [11],\PWMC/n26 [8]}),
    .clk(clk100m),
    .d({\PWMC/pnumr [11],\PWMC/pnumr [8]}),
    .mi({\U_AHB/h2h_hwdata [11],\U_AHB/h2h_hwdata [8]}),
    .sr(\U_AHB/n71 ),
    .f({_al_u2708_o,_al_u2670_o}),
    .q({pnumC[11],pnumC[8]}));  // src/AHB.v(79)
  // src/AHB.v(79)
  // src/AHB.v(79)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg30_b12|U_AHB/reg30_b7  (
    .a({\PWMC/n24 ,\PWMC/n24 }),
    .b({\PWMC/n25_neg_lutinv ,\PWMC/n25_neg_lutinv }),
    .c({\PWMC/n26 [12],\PWMC/n26 [7]}),
    .clk(clk100m),
    .d({\PWMC/pnumr [12],\PWMC/pnumr [7]}),
    .mi({\U_AHB/h2h_hwdata [12],\U_AHB/h2h_hwdata [7]}),
    .sr(\U_AHB/n71 ),
    .f({_al_u2706_o,_al_u2672_o}),
    .q({pnumC[12],pnumC[7]}));  // src/AHB.v(79)
  // src/AHB.v(79)
  // src/AHB.v(79)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg30_b13|U_AHB/reg30_b6  (
    .a({\PWMC/n24 ,\PWMC/n24 }),
    .b({\PWMC/n25_neg_lutinv ,\PWMC/n25_neg_lutinv }),
    .c({\PWMC/n26 [13],\PWMC/n26 [6]}),
    .clk(clk100m),
    .d({\PWMC/pnumr [13],\PWMC/pnumr [6]}),
    .mi({\U_AHB/h2h_hwdata [13],\U_AHB/h2h_hwdata [6]}),
    .sr(\U_AHB/n71 ),
    .f({_al_u2704_o,_al_u2674_o}),
    .q({pnumC[13],pnumC[6]}));  // src/AHB.v(79)
  // src/AHB.v(79)
  // src/AHB.v(79)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg30_b14|U_AHB/reg30_b5  (
    .a({\PWMC/n24 ,\PWMC/n24 }),
    .b({\PWMC/n25_neg_lutinv ,\PWMC/n25_neg_lutinv }),
    .c({\PWMC/n26 [14],\PWMC/n26 [5]}),
    .clk(clk100m),
    .d({\PWMC/pnumr [14],\PWMC/pnumr [5]}),
    .mi({\U_AHB/h2h_hwdata [14],\U_AHB/h2h_hwdata [5]}),
    .sr(\U_AHB/n71 ),
    .f({_al_u2702_o,_al_u2676_o}),
    .q({pnumC[14],pnumC[5]}));  // src/AHB.v(79)
  // src/AHB.v(79)
  // src/AHB.v(79)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg30_b15|U_AHB/reg30_b4  (
    .a({\PWMC/n24 ,\PWMC/n24 }),
    .b({\PWMC/n25_neg_lutinv ,\PWMC/n25_neg_lutinv }),
    .c({\PWMC/n26 [15],\PWMC/n26 [4]}),
    .clk(clk100m),
    .d({\PWMC/pnumr [15],\PWMC/pnumr [4]}),
    .mi({\U_AHB/h2h_hwdata [15],\U_AHB/h2h_hwdata [4]}),
    .sr(\U_AHB/n71 ),
    .f({_al_u2700_o,_al_u2678_o}),
    .q({pnumC[15],pnumC[4]}));  // src/AHB.v(79)
  // src/AHB.v(79)
  // src/AHB.v(79)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg30_b16|U_AHB/reg30_b3  (
    .a({\PWMC/n24 ,\PWMC/n24 }),
    .b({\PWMC/n25_neg_lutinv ,\PWMC/n25_neg_lutinv }),
    .c({\PWMC/n26 [16],\PWMC/n26 [3]}),
    .clk(clk100m),
    .d({\PWMC/pnumr [16],\PWMC/pnumr [3]}),
    .mi({\U_AHB/h2h_hwdata [16],\U_AHB/h2h_hwdata [3]}),
    .sr(\U_AHB/n71 ),
    .f({_al_u2698_o,_al_u2680_o}),
    .q({pnumC[16],pnumC[3]}));  // src/AHB.v(79)
  // src/AHB.v(79)
  // src/AHB.v(79)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg30_b17|U_AHB/reg30_b23  (
    .a({\PWMC/n24 ,\PWMC/n24 }),
    .b({\PWMC/n25_neg_lutinv ,\PWMC/n25_neg_lutinv }),
    .c({\PWMC/n26 [17],\PWMC/n26 [23]}),
    .clk(clk100m),
    .d({\PWMC/pnumr [17],\PWMC/pnumr [23]}),
    .mi({\U_AHB/h2h_hwdata [17],\U_AHB/h2h_hwdata [23]}),
    .sr(\U_AHB/n71 ),
    .f({_al_u2696_o,_al_u2682_o}),
    .q({pnumC[17],pnumC[23]}));  // src/AHB.v(79)
  // src/AHB.v(79)
  // src/AHB.v(79)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg30_b18|U_AHB/reg30_b22  (
    .a({\PWMC/n24 ,\PWMC/n24 }),
    .b({\PWMC/n25_neg_lutinv ,\PWMC/n25_neg_lutinv }),
    .c({\PWMC/n26 [18],\PWMC/n26 [22]}),
    .clk(clk100m),
    .d({\PWMC/pnumr [18],\PWMC/pnumr [22]}),
    .mi({\U_AHB/h2h_hwdata [18],\U_AHB/h2h_hwdata [22]}),
    .sr(\U_AHB/n71 ),
    .f({_al_u2694_o,_al_u2684_o}),
    .q({pnumC[18],pnumC[22]}));  // src/AHB.v(79)
  // src/AHB.v(79)
  // src/AHB.v(79)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg30_b19|U_AHB/reg30_b21  (
    .a({\PWMC/n24 ,\PWMC/n24 }),
    .b({\PWMC/n25_neg_lutinv ,\PWMC/n25_neg_lutinv }),
    .c({\PWMC/n26 [19],\PWMC/n26 [21]}),
    .clk(clk100m),
    .d({\PWMC/pnumr [19],\PWMC/pnumr [21]}),
    .mi({\U_AHB/h2h_hwdata [19],\U_AHB/h2h_hwdata [21]}),
    .sr(\U_AHB/n71 ),
    .f({_al_u2692_o,_al_u2686_o}),
    .q({pnumC[19],pnumC[21]}));  // src/AHB.v(79)
  // src/AHB.v(79)
  // src/AHB.v(79)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg30_b1|U_AHB/reg30_b20  (
    .a({\PWMC/n24 ,\PWMC/n24 }),
    .b({\PWMC/n25_neg_lutinv ,\PWMC/n25_neg_lutinv }),
    .c({\PWMC/n26 [1],\PWMC/n26 [20]}),
    .clk(clk100m),
    .d({\PWMC/pnumr [1],\PWMC/pnumr [20]}),
    .mi({\U_AHB/h2h_hwdata [1],\U_AHB/h2h_hwdata [20]}),
    .sr(\U_AHB/n71 ),
    .f({_al_u2712_o,_al_u2688_o}),
    .q({pnumC[1],pnumC[20]}));  // src/AHB.v(79)
  // src/AHB.v(79)
  // src/AHB.v(79)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b0000000000001111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg30_b24|U_AHB/reg30_b2  (
    .a({open_n31400,\PWMC/n24 }),
    .b({open_n31401,\PWMC/n25_neg_lutinv }),
    .c({_al_u2988_o,\PWMC/n26 [2]}),
    .clk(clk100m),
    .d({_al_u1652_o,\PWMC/pnumr [2]}),
    .mi({\U_AHB/h2h_hwdata [24],\U_AHB/h2h_hwdata [2]}),
    .sr(\U_AHB/n71 ),
    .f({_al_u3055_o,_al_u2690_o}),
    .q({pnumC[24],pnumC[2]}));  // src/AHB.v(79)
  // src/AHB.v(79)
  // src/AHB.v(79)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("~(C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000111111111111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg30_b27|U_AHB/reg30_b26  (
    .c({_al_u3055_o,n4_neg}),
    .clk(clk100m),
    .d({_al_u2984_o,_al_u2983_o}),
    .mi(\U_AHB/h2h_hwdata [27:26]),
    .sr(\U_AHB/n71 ),
    .f({_al_n1_en,_al_u2984_o}),
    .q(pnumC[27:26]));  // src/AHB.v(79)
  // src/AHB.v(79)
  // src/AHB.v(79)
  EF2_PHY_LSLICE #(
    //.LUTF0("(D*C*B*A)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(D*C*B*A)"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000000000000000),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg30_b29|U_AHB/reg30_b25  (
    .a({open_n31434,_al_u1647_o}),
    .b({_al_u1640_o,_al_u1648_o}),
    .c({_al_u1648_o,_al_u1650_o}),
    .clk(clk100m),
    .d({_al_u2982_o,_al_u1651_o}),
    .mi({\U_AHB/h2h_hwdata [29],\U_AHB/h2h_hwdata [25]}),
    .sr(\U_AHB/n71 ),
    .f({_al_u2983_o,_al_u1652_o}),
    .q({pnumC[29],pnumC[25]}));  // src/AHB.v(79)
  // src/AHB.v(79)
  // src/AHB.v(79)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*B*A)"),
    //.LUTF1("(D*~C*~B*A)"),
    //.LUTG0("(~1*~D*~C*B*A)"),
    //.LUTG1("(D*~C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001000),
    .INIT_LUTF1(16'b0000001000000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000001000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg30_b31|U_AHB/reg30_b9  (
    .a({_al_u1638_o,_al_u1638_o}),
    .b({timer[10],_al_u1639_o}),
    .c(timer[11:10]),
    .clk(clk100m),
    .d({timer[8],timer[11]}),
    .e({open_n31454,timer[8]}),
    .mi({\U_AHB/h2h_hwdata [31],\U_AHB/h2h_hwdata [9]}),
    .sr(\U_AHB/n71 ),
    .f({_al_u1647_o,_al_u1640_o}),
    .q({pnumC[31],pnumC[9]}));  // src/AHB.v(79)
  // src/AHB.v(80)
  // src/AHB.v(80)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg31_b0|U_AHB/reg31_b32  (
    .a({\PWMD/n24 ,\PWMD/n24 }),
    .b({\PWMD/n25_neg_lutinv ,\PWMD/n25_neg_lutinv }),
    .c({\PWMD/n26 [0],\PWMD/n26 [9]}),
    .clk(clk100m),
    .d({\PWMD/pnumr [0],\PWMD/pnumr [9]}),
    .mi({\U_AHB/h2h_hwdata [0],1'b1}),
    .sr(\U_AHB/n73 ),
    .f({_al_u2793_o,_al_u2747_o}),
    .q({pnumD[0],pnumD[32]}));  // src/AHB.v(80)
  // src/AHB.v(80)
  // src/AHB.v(80)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg31_b10|U_AHB/reg31_b8  (
    .a({\PWMD/n24 ,\PWMD/n24 }),
    .b({\PWMD/n25_neg_lutinv ,\PWMD/n25_neg_lutinv }),
    .c({\PWMD/n26 [10],\PWMD/n26 [8]}),
    .clk(clk100m),
    .d({\PWMD/pnumr [10],\PWMD/pnumr [8]}),
    .mi({\U_AHB/h2h_hwdata [10],\U_AHB/h2h_hwdata [8]}),
    .sr(\U_AHB/n73 ),
    .f({_al_u2789_o,_al_u2749_o}),
    .q({pnumD[10],pnumD[8]}));  // src/AHB.v(80)
  // src/AHB.v(80)
  // src/AHB.v(80)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg31_b11|U_AHB/reg31_b7  (
    .a({\PWMD/n24 ,\PWMD/n24 }),
    .b({\PWMD/n25_neg_lutinv ,\PWMD/n25_neg_lutinv }),
    .c({\PWMD/n26 [11],\PWMD/n26 [7]}),
    .clk(clk100m),
    .d({\PWMD/pnumr [11],\PWMD/pnumr [7]}),
    .mi({\U_AHB/h2h_hwdata [11],\U_AHB/h2h_hwdata [7]}),
    .sr(\U_AHB/n73 ),
    .f({_al_u2787_o,_al_u2751_o}),
    .q({pnumD[11],pnumD[7]}));  // src/AHB.v(80)
  // src/AHB.v(80)
  // src/AHB.v(80)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg31_b12|U_AHB/reg31_b6  (
    .a({\PWMD/n24 ,\PWMD/n24 }),
    .b({\PWMD/n25_neg_lutinv ,\PWMD/n25_neg_lutinv }),
    .c({\PWMD/n26 [12],\PWMD/n26 [6]}),
    .clk(clk100m),
    .d({\PWMD/pnumr [12],\PWMD/pnumr [6]}),
    .mi({\U_AHB/h2h_hwdata [12],\U_AHB/h2h_hwdata [6]}),
    .sr(\U_AHB/n73 ),
    .f({_al_u2785_o,_al_u2753_o}),
    .q({pnumD[12],pnumD[6]}));  // src/AHB.v(80)
  // src/AHB.v(80)
  // src/AHB.v(80)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg31_b13|U_AHB/reg31_b5  (
    .a({\PWMD/n24 ,\PWMD/n24 }),
    .b({\PWMD/n25_neg_lutinv ,\PWMD/n25_neg_lutinv }),
    .c({\PWMD/n26 [13],\PWMD/n26 [5]}),
    .clk(clk100m),
    .d({\PWMD/pnumr [13],\PWMD/pnumr [5]}),
    .mi({\U_AHB/h2h_hwdata [13],\U_AHB/h2h_hwdata [5]}),
    .sr(\U_AHB/n73 ),
    .f({_al_u2783_o,_al_u2755_o}),
    .q({pnumD[13],pnumD[5]}));  // src/AHB.v(80)
  // src/AHB.v(80)
  // src/AHB.v(80)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg31_b14|U_AHB/reg31_b4  (
    .a({\PWMD/n24 ,\PWMD/n24 }),
    .b({\PWMD/n25_neg_lutinv ,\PWMD/n25_neg_lutinv }),
    .c({\PWMD/n26 [14],\PWMD/n26 [4]}),
    .clk(clk100m),
    .d({\PWMD/pnumr [14],\PWMD/pnumr [4]}),
    .mi({\U_AHB/h2h_hwdata [14],\U_AHB/h2h_hwdata [4]}),
    .sr(\U_AHB/n73 ),
    .f({_al_u2781_o,_al_u2757_o}),
    .q({pnumD[14],pnumD[4]}));  // src/AHB.v(80)
  // src/AHB.v(80)
  // src/AHB.v(80)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg31_b15|U_AHB/reg31_b3  (
    .a({\PWMD/n24 ,\PWMD/n24 }),
    .b({\PWMD/n25_neg_lutinv ,\PWMD/n25_neg_lutinv }),
    .c({\PWMD/n26 [15],\PWMD/n26 [3]}),
    .clk(clk100m),
    .d({\PWMD/pnumr [15],\PWMD/pnumr [3]}),
    .mi({\U_AHB/h2h_hwdata [15],\U_AHB/h2h_hwdata [3]}),
    .sr(\U_AHB/n73 ),
    .f({_al_u2779_o,_al_u2759_o}),
    .q({pnumD[15],pnumD[3]}));  // src/AHB.v(80)
  // src/AHB.v(80)
  // src/AHB.v(80)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg31_b16|U_AHB/reg31_b23  (
    .a({\PWMD/n24 ,\PWMD/n24 }),
    .b({\PWMD/n25_neg_lutinv ,\PWMD/n25_neg_lutinv }),
    .c({\PWMD/n26 [16],\PWMD/n26 [23]}),
    .clk(clk100m),
    .d({\PWMD/pnumr [16],\PWMD/pnumr [23]}),
    .mi({\U_AHB/h2h_hwdata [16],\U_AHB/h2h_hwdata [23]}),
    .sr(\U_AHB/n73 ),
    .f({_al_u2777_o,_al_u2761_o}),
    .q({pnumD[16],pnumD[23]}));  // src/AHB.v(80)
  // src/AHB.v(80)
  // src/AHB.v(80)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg31_b17|U_AHB/reg31_b22  (
    .a({\PWMD/n24 ,\PWMD/n24 }),
    .b({\PWMD/n25_neg_lutinv ,\PWMD/n25_neg_lutinv }),
    .c({\PWMD/n26 [17],\PWMD/n26 [22]}),
    .clk(clk100m),
    .d({\PWMD/pnumr [17],\PWMD/pnumr [22]}),
    .mi({\U_AHB/h2h_hwdata [17],\U_AHB/h2h_hwdata [22]}),
    .sr(\U_AHB/n73 ),
    .f({_al_u2775_o,_al_u2763_o}),
    .q({pnumD[17],pnumD[22]}));  // src/AHB.v(80)
  // src/AHB.v(80)
  // src/AHB.v(80)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg31_b18|U_AHB/reg31_b21  (
    .a({\PWMD/n24 ,\PWMD/n24 }),
    .b({\PWMD/n25_neg_lutinv ,\PWMD/n25_neg_lutinv }),
    .c({\PWMD/n26 [18],\PWMD/n26 [21]}),
    .clk(clk100m),
    .d({\PWMD/pnumr [18],\PWMD/pnumr [21]}),
    .mi({\U_AHB/h2h_hwdata [18],\U_AHB/h2h_hwdata [21]}),
    .sr(\U_AHB/n73 ),
    .f({_al_u2773_o,_al_u2765_o}),
    .q({pnumD[18],pnumD[21]}));  // src/AHB.v(80)
  // src/AHB.v(80)
  // src/AHB.v(80)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg31_b19|U_AHB/reg31_b20  (
    .a({\PWMD/n24 ,\PWMD/n24 }),
    .b({\PWMD/n25_neg_lutinv ,\PWMD/n25_neg_lutinv }),
    .c({\PWMD/n26 [19],\PWMD/n26 [20]}),
    .clk(clk100m),
    .d({\PWMD/pnumr [19],\PWMD/pnumr [20]}),
    .mi({\U_AHB/h2h_hwdata [19],\U_AHB/h2h_hwdata [20]}),
    .sr(\U_AHB/n73 ),
    .f({_al_u2771_o,_al_u2767_o}),
    .q({pnumD[19],pnumD[20]}));  // src/AHB.v(80)
  // src/AHB.v(80)
  // src/AHB.v(80)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg31_b1|U_AHB/reg31_b2  (
    .a({\PWMD/n24 ,\PWMD/n24 }),
    .b({\PWMD/n25_neg_lutinv ,\PWMD/n25_neg_lutinv }),
    .c({\PWMD/n26 [1],\PWMD/n26 [2]}),
    .clk(clk100m),
    .d({\PWMD/pnumr [1],\PWMD/pnumr [2]}),
    .mi({\U_AHB/h2h_hwdata [1],\U_AHB/h2h_hwdata [2]}),
    .sr(\U_AHB/n73 ),
    .f({_al_u2791_o,_al_u2769_o}),
    .q({pnumD[1],pnumD[2]}));  // src/AHB.v(80)
  // src/AHB.v(80)
  // src/AHB.v(80)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*D*C*B*A)"),
    //.LUTF1("(0*D*C*B*A)"),
    //.LUTG0("(~1*D*C*B*A)"),
    //.LUTG1("(1*D*C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000000000000000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg31_b24|U_AHB/reg31_b25  (
    .a({_al_u1641_o,_al_u1641_o}),
    .b({timer[4],timer[4]}),
    .c({timer[5],timer[5]}),
    .clk(clk100m),
    .d({timer[6],timer[6]}),
    .e({timer[7],timer[7]}),
    .mi({\U_AHB/h2h_hwdata [24],\U_AHB/h2h_hwdata [25]}),
    .sr(\U_AHB/n73 ),
    .f({_al_u1648_o,_al_u1642_o}),
    .q({pnumD[24],pnumD[25]}));  // src/AHB.v(80)
  // src/AHB.v(80)
  // src/AHB.v(80)
  EF2_PHY_MSLICE #(
    //.LUT0("(D*C*B*A)"),
    //.LUT1("(D*~C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000000000000000),
    .INIT_LUT1(16'b0000100000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg31_b29|U_AHB/reg31_b26  (
    .a({timer[14],timer[0]}),
    .b({timer[15],timer[1]}),
    .c({timer[26],timer[2]}),
    .clk(clk100m),
    .d({timer[27],timer[3]}),
    .mi({\U_AHB/h2h_hwdata [29],\U_AHB/h2h_hwdata [26]}),
    .sr(\U_AHB/n73 ),
    .f({_al_u2985_o,_al_u1641_o}),
    .q({pnumD[29],pnumD[26]}));  // src/AHB.v(80)
  // src/AHB.v(80)
  // src/AHB.v(80)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*C*~B*A)"),
    //.LUTF1("(~0*D*~C*B*A)"),
    //.LUTG0("(~1*~D*C*~B*A)"),
    //.LUTG1("(~1*D*~C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000100000),
    .INIT_LUTF1(16'b0000100000000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg31_b30|U_AHB/reg31_b9  (
    .a({_al_u2981_o,_al_u1643_o}),
    .b({timer[24],timer[24]}),
    .c({timer[25],timer[25]}),
    .clk(clk100m),
    .d({timer[26],timer[26]}),
    .e({timer[27],timer[27]}),
    .mi({\U_AHB/h2h_hwdata [30],\U_AHB/h2h_hwdata [9]}),
    .sr(\U_AHB/n73 ),
    .f({_al_u2982_o,_al_u1644_o}),
    .q({pnumD[30],pnumD[9]}));  // src/AHB.v(80)
  // src/AHB.v(81)
  // src/AHB.v(81)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg32_b0|U_AHB/reg32_b32  (
    .a({\PWME/n24 ,\PWME/n24 }),
    .b({\PWME/n25_neg_lutinv ,\PWME/n25_neg_lutinv }),
    .c({\PWME/n26 [0],\PWME/n26 [9]}),
    .clk(clk100m),
    .d({\PWME/pnumr [0],\PWME/pnumr [9]}),
    .mi({\U_AHB/h2h_hwdata [0],1'b1}),
    .sr(\U_AHB/n75 ),
    .f({_al_u2873_o,_al_u2827_o}),
    .q({pnumE[0],pnumE[32]}));  // src/AHB.v(81)
  // src/AHB.v(81)
  // src/AHB.v(81)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg32_b10|U_AHB/reg32_b8  (
    .a({\PWME/n24 ,\PWME/n24 }),
    .b({\PWME/n25_neg_lutinv ,\PWME/n25_neg_lutinv }),
    .c({\PWME/n26 [10],\PWME/n26 [8]}),
    .clk(clk100m),
    .d({\PWME/pnumr [10],\PWME/pnumr [8]}),
    .mi({\U_AHB/h2h_hwdata [10],\U_AHB/h2h_hwdata [8]}),
    .sr(\U_AHB/n75 ),
    .f({_al_u2869_o,_al_u2829_o}),
    .q({pnumE[10],pnumE[8]}));  // src/AHB.v(81)
  // src/AHB.v(81)
  // src/AHB.v(81)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg32_b11|U_AHB/reg32_b7  (
    .a({\PWME/n24 ,\PWME/n24 }),
    .b({\PWME/n25_neg_lutinv ,\PWME/n25_neg_lutinv }),
    .c({\PWME/n26 [11],\PWME/n26 [7]}),
    .clk(clk100m),
    .d({\PWME/pnumr [11],\PWME/pnumr [7]}),
    .mi({\U_AHB/h2h_hwdata [11],\U_AHB/h2h_hwdata [7]}),
    .sr(\U_AHB/n75 ),
    .f({_al_u2867_o,_al_u2831_o}),
    .q({pnumE[11],pnumE[7]}));  // src/AHB.v(81)
  // src/AHB.v(81)
  // src/AHB.v(81)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg32_b12|U_AHB/reg32_b6  (
    .a({\PWME/n24 ,\PWME/n24 }),
    .b({\PWME/n25_neg_lutinv ,\PWME/n25_neg_lutinv }),
    .c({\PWME/n26 [12],\PWME/n26 [6]}),
    .clk(clk100m),
    .d({\PWME/pnumr [12],\PWME/pnumr [6]}),
    .mi({\U_AHB/h2h_hwdata [12],\U_AHB/h2h_hwdata [6]}),
    .sr(\U_AHB/n75 ),
    .f({_al_u2865_o,_al_u2833_o}),
    .q({pnumE[12],pnumE[6]}));  // src/AHB.v(81)
  // src/AHB.v(81)
  // src/AHB.v(81)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg32_b13|U_AHB/reg32_b5  (
    .a({\PWME/n24 ,\PWME/n24 }),
    .b({\PWME/n25_neg_lutinv ,\PWME/n25_neg_lutinv }),
    .c({\PWME/n26 [13],\PWME/n26 [5]}),
    .clk(clk100m),
    .d({\PWME/pnumr [13],\PWME/pnumr [5]}),
    .mi({\U_AHB/h2h_hwdata [13],\U_AHB/h2h_hwdata [5]}),
    .sr(\U_AHB/n75 ),
    .f({_al_u2863_o,_al_u2835_o}),
    .q({pnumE[13],pnumE[5]}));  // src/AHB.v(81)
  // src/AHB.v(81)
  // src/AHB.v(81)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg32_b14|U_AHB/reg32_b4  (
    .a({\PWME/n24 ,\PWME/n24 }),
    .b({\PWME/n25_neg_lutinv ,\PWME/n25_neg_lutinv }),
    .c({\PWME/n26 [14],\PWME/n26 [4]}),
    .clk(clk100m),
    .d({\PWME/pnumr [14],\PWME/pnumr [4]}),
    .mi({\U_AHB/h2h_hwdata [14],\U_AHB/h2h_hwdata [4]}),
    .sr(\U_AHB/n75 ),
    .f({_al_u2861_o,_al_u2837_o}),
    .q({pnumE[14],pnumE[4]}));  // src/AHB.v(81)
  // src/AHB.v(81)
  // src/AHB.v(81)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg32_b15|U_AHB/reg32_b3  (
    .a({\PWME/n24 ,\PWME/n24 }),
    .b({\PWME/n25_neg_lutinv ,\PWME/n25_neg_lutinv }),
    .c({\PWME/n26 [15],\PWME/n26 [3]}),
    .clk(clk100m),
    .d({\PWME/pnumr [15],\PWME/pnumr [3]}),
    .mi({\U_AHB/h2h_hwdata [15],\U_AHB/h2h_hwdata [3]}),
    .sr(\U_AHB/n75 ),
    .f({_al_u2859_o,_al_u2839_o}),
    .q({pnumE[15],pnumE[3]}));  // src/AHB.v(81)
  // src/AHB.v(81)
  // src/AHB.v(81)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg32_b16|U_AHB/reg32_b23  (
    .a({\PWME/n24 ,\PWME/n24 }),
    .b({\PWME/n25_neg_lutinv ,\PWME/n25_neg_lutinv }),
    .c({\PWME/n26 [16],\PWME/n26 [23]}),
    .clk(clk100m),
    .d({\PWME/pnumr [16],\PWME/pnumr [23]}),
    .mi({\U_AHB/h2h_hwdata [16],\U_AHB/h2h_hwdata [23]}),
    .sr(\U_AHB/n75 ),
    .f({_al_u2857_o,_al_u2841_o}),
    .q({pnumE[16],pnumE[23]}));  // src/AHB.v(81)
  // src/AHB.v(81)
  // src/AHB.v(81)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg32_b17|U_AHB/reg32_b22  (
    .a({\PWME/n24 ,\PWME/n24 }),
    .b({\PWME/n25_neg_lutinv ,\PWME/n25_neg_lutinv }),
    .c({\PWME/n26 [17],\PWME/n26 [22]}),
    .clk(clk100m),
    .d({\PWME/pnumr [17],\PWME/pnumr [22]}),
    .mi({\U_AHB/h2h_hwdata [17],\U_AHB/h2h_hwdata [22]}),
    .sr(\U_AHB/n75 ),
    .f({_al_u2855_o,_al_u2843_o}),
    .q({pnumE[17],pnumE[22]}));  // src/AHB.v(81)
  // src/AHB.v(81)
  // src/AHB.v(81)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg32_b18|U_AHB/reg32_b21  (
    .a({\PWME/n24 ,\PWME/n24 }),
    .b({\PWME/n25_neg_lutinv ,\PWME/n25_neg_lutinv }),
    .c({\PWME/n26 [18],\PWME/n26 [21]}),
    .clk(clk100m),
    .d({\PWME/pnumr [18],\PWME/pnumr [21]}),
    .mi({\U_AHB/h2h_hwdata [18],\U_AHB/h2h_hwdata [21]}),
    .sr(\U_AHB/n75 ),
    .f({_al_u2853_o,_al_u2845_o}),
    .q({pnumE[18],pnumE[21]}));  // src/AHB.v(81)
  // src/AHB.v(81)
  // src/AHB.v(81)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg32_b19|U_AHB/reg32_b20  (
    .a({\PWME/n24 ,\PWME/n24 }),
    .b({\PWME/n25_neg_lutinv ,\PWME/n25_neg_lutinv }),
    .c({\PWME/n26 [19],\PWME/n26 [20]}),
    .clk(clk100m),
    .d({\PWME/pnumr [19],\PWME/pnumr [20]}),
    .mi({\U_AHB/h2h_hwdata [19],\U_AHB/h2h_hwdata [20]}),
    .sr(\U_AHB/n75 ),
    .f({_al_u2851_o,_al_u2847_o}),
    .q({pnumE[19],pnumE[20]}));  // src/AHB.v(81)
  // src/AHB.v(81)
  // src/AHB.v(81)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg32_b1|U_AHB/reg32_b2  (
    .a({\PWME/n24 ,\PWME/n24 }),
    .b({\PWME/n25_neg_lutinv ,\PWME/n25_neg_lutinv }),
    .c({\PWME/n26 [1],\PWME/n26 [2]}),
    .clk(clk100m),
    .d({\PWME/pnumr [1],\PWME/pnumr [2]}),
    .mi({\U_AHB/h2h_hwdata [1],\U_AHB/h2h_hwdata [2]}),
    .sr(\U_AHB/n75 ),
    .f({_al_u2871_o,_al_u2849_o}),
    .q({pnumE[1],pnumE[2]}));  // src/AHB.v(81)
  // src/AHB.v(81)
  // src/AHB.v(81)
  EF2_PHY_LSLICE #(
    //.LUTF0("(0*D*C*~B*A)"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(1*D*C*~B*A)"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0010000000000000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg32_b26|U_AHB/reg32_b25  (
    .a({timer[20],_al_u1645_o}),
    .b(timer[21:20]),
    .c(timer[22:21]),
    .clk(clk100m),
    .d({timer[23],timer[24]}),
    .e({open_n31853,timer[25]}),
    .mi(\U_AHB/h2h_hwdata [26:25]),
    .sr(\U_AHB/n75 ),
    .f({_al_u1639_o,_al_u1651_o}),
    .q(pnumE[26:25]));  // src/AHB.v(81)
  // src/AHB.v(81)
  // src/AHB.v(81)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(~0*D*~C*B*A)"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(~1*D*~C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000100000000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg32_b27|U_AHB/reg32_b24  (
    .a({_al_u2980_o,_al_u1639_o}),
    .b({timer[16],timer[18]}),
    .c({timer[17],timer[19]}),
    .clk(clk100m),
    .d({timer[18],timer[24]}),
    .e({timer[19],timer[25]}),
    .mi({\U_AHB/h2h_hwdata [27],\U_AHB/h2h_hwdata [24]}),
    .sr(\U_AHB/n75 ),
    .f({_al_u2981_o,_al_u2987_o}),
    .q({pnumE[27],pnumE[24]}));  // src/AHB.v(81)
  // src/AHB.v(81)
  // src/AHB.v(81)
  EF2_PHY_LSLICE #(
    //.LUTF0("(D*C*B*~A)"),
    //.LUTF1("(D*~C*B*A)"),
    //.LUTG0("(D*C*B*~A)"),
    //.LUTG1("(D*~C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100000000000000),
    .INIT_LUTF1(16'b0000100000000000),
    .INIT_LUTG0(16'b0100000000000000),
    .INIT_LUTG1(16'b0000100000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg32_b28|U_AHB/reg32_b9  (
    .a({timer[14],timer[12]}),
    .b({timer[15],timer[13]}),
    .c({timer[18],timer[14]}),
    .clk(clk100m),
    .d({timer[19],timer[15]}),
    .mi({\U_AHB/h2h_hwdata [28],\U_AHB/h2h_hwdata [9]}),
    .sr(\U_AHB/n75 ),
    .f({_al_u1645_o,_al_u2980_o}),
    .q({pnumE[28],pnumE[9]}));  // src/AHB.v(81)
  // src/AHB.v(81)
  // src/AHB.v(81)
  EF2_PHY_LSLICE #(
    //.LUTF0("(0*D*~C*~B*A)"),
    //.LUTF1("(~0*~D*~C*B*A)"),
    //.LUTG0("(1*D*~C*~B*A)"),
    //.LUTG1("(~1*~D*~C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000000000001000),
    .INIT_LUTG0(16'b0000001000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg32_b29|U_AHB/reg32_b30  (
    .a({_al_u2985_o,_al_u1649_o}),
    .b({timer[12],timer[12]}),
    .c({timer[13],timer[13]}),
    .clk(clk100m),
    .d({timer[16],timer[16]}),
    .e({timer[17],timer[17]}),
    .mi({\U_AHB/h2h_hwdata [29],\U_AHB/h2h_hwdata [30]}),
    .sr(\U_AHB/n75 ),
    .f({_al_u2986_o,_al_u1650_o}),
    .q({pnumE[29],pnumE[30]}));  // src/AHB.v(81)
  // src/AHB.v(82)
  // src/AHB.v(82)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b1010100000100000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1010100000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg33_b0|U_AHB/reg33_b24  (
    .a({\PWMF/n24 ,_al_u2339_o}),
    .b({\PWMF/n25_neg_lutinv ,pnumcnt8[6]}),
    .c({\PWMF/n26 [0],pnumcnt8[7]}),
    .clk(clk100m),
    .d({\PWMF/pnumr [0],pnumcnt8[8]}),
    .e({open_n31920,pnumcnt8[9]}),
    .mi({\U_AHB/h2h_hwdata [0],\U_AHB/h2h_hwdata [24]}),
    .sr(\U_AHB/n77 ),
    .f({_al_u2952_o,_al_u2340_o}),
    .q({pnumF[0],pnumF[24]}));  // src/AHB.v(82)
  // src/AHB.v(82)
  // src/AHB.v(82)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b1010100000100000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1010100000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg33_b10|U_AHB/reg33_b31  (
    .a({\PWMF/n24 ,_al_u2900_o}),
    .b({\PWMF/n25_neg_lutinv ,pnumcntF[6]}),
    .c({\PWMF/n26 [10],pnumcntF[7]}),
    .clk(clk100m),
    .d({\PWMF/pnumr [10],pnumcntF[8]}),
    .e({open_n31937,pnumcntF[9]}),
    .mi({\U_AHB/h2h_hwdata [10],\U_AHB/h2h_hwdata [31]}),
    .sr(\U_AHB/n77 ),
    .f({_al_u2948_o,_al_u2901_o}),
    .q({pnumF[10],pnumF[31]}));  // src/AHB.v(82)
  // src/AHB.v(82)
  // src/AHB.v(82)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg33_b11|U_AHB/reg33_b32  (
    .a({\PWMF/n24 ,\PWMF/n24 }),
    .b({\PWMF/n25_neg_lutinv ,\PWMF/n25_neg_lutinv }),
    .c({\PWMF/n26 [11],\PWMF/n26 [9]}),
    .clk(clk100m),
    .d({\PWMF/pnumr [11],\PWMF/pnumr [9]}),
    .mi({\U_AHB/h2h_hwdata [11],1'b1}),
    .sr(\U_AHB/n77 ),
    .f({_al_u2946_o,_al_u2906_o}),
    .q({pnumF[11],pnumF[32]}));  // src/AHB.v(82)
  // src/AHB.v(82)
  // src/AHB.v(82)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg33_b12|U_AHB/reg33_b8  (
    .a({\PWMF/n24 ,\PWMF/n24 }),
    .b({\PWMF/n25_neg_lutinv ,\PWMF/n25_neg_lutinv }),
    .c({\PWMF/n26 [12],\PWMF/n26 [8]}),
    .clk(clk100m),
    .d({\PWMF/pnumr [12],\PWMF/pnumr [8]}),
    .mi({\U_AHB/h2h_hwdata [12],\U_AHB/h2h_hwdata [8]}),
    .sr(\U_AHB/n77 ),
    .f({_al_u2944_o,_al_u2908_o}),
    .q({pnumF[12],pnumF[8]}));  // src/AHB.v(82)
  // src/AHB.v(82)
  // src/AHB.v(82)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg33_b13|U_AHB/reg33_b7  (
    .a({\PWMF/n24 ,\PWMF/n24 }),
    .b({\PWMF/n25_neg_lutinv ,\PWMF/n25_neg_lutinv }),
    .c({\PWMF/n26 [13],\PWMF/n26 [7]}),
    .clk(clk100m),
    .d({\PWMF/pnumr [13],\PWMF/pnumr [7]}),
    .mi({\U_AHB/h2h_hwdata [13],\U_AHB/h2h_hwdata [7]}),
    .sr(\U_AHB/n77 ),
    .f({_al_u2942_o,_al_u2910_o}),
    .q({pnumF[13],pnumF[7]}));  // src/AHB.v(82)
  // src/AHB.v(82)
  // src/AHB.v(82)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg33_b14|U_AHB/reg33_b6  (
    .a({\PWMF/n24 ,\PWMF/n24 }),
    .b({\PWMF/n25_neg_lutinv ,\PWMF/n25_neg_lutinv }),
    .c({\PWMF/n26 [14],\PWMF/n26 [6]}),
    .clk(clk100m),
    .d({\PWMF/pnumr [14],\PWMF/pnumr [6]}),
    .mi({\U_AHB/h2h_hwdata [14],\U_AHB/h2h_hwdata [6]}),
    .sr(\U_AHB/n77 ),
    .f({_al_u2940_o,_al_u2912_o}),
    .q({pnumF[14],pnumF[6]}));  // src/AHB.v(82)
  // src/AHB.v(82)
  // src/AHB.v(82)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg33_b15|U_AHB/reg33_b5  (
    .a({\PWMF/n24 ,\PWMF/n24 }),
    .b({\PWMF/n25_neg_lutinv ,\PWMF/n25_neg_lutinv }),
    .c({\PWMF/n26 [15],\PWMF/n26 [5]}),
    .clk(clk100m),
    .d({\PWMF/pnumr [15],\PWMF/pnumr [5]}),
    .mi({\U_AHB/h2h_hwdata [15],\U_AHB/h2h_hwdata [5]}),
    .sr(\U_AHB/n77 ),
    .f({_al_u2938_o,_al_u2914_o}),
    .q({pnumF[15],pnumF[5]}));  // src/AHB.v(82)
  // src/AHB.v(82)
  // src/AHB.v(82)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg33_b16|U_AHB/reg33_b4  (
    .a({\PWMF/n24 ,\PWMF/n24 }),
    .b({\PWMF/n25_neg_lutinv ,\PWMF/n25_neg_lutinv }),
    .c({\PWMF/n26 [16],\PWMF/n26 [4]}),
    .clk(clk100m),
    .d({\PWMF/pnumr [16],\PWMF/pnumr [4]}),
    .mi({\U_AHB/h2h_hwdata [16],\U_AHB/h2h_hwdata [4]}),
    .sr(\U_AHB/n77 ),
    .f({_al_u2936_o,_al_u2916_o}),
    .q({pnumF[16],pnumF[4]}));  // src/AHB.v(82)
  // src/AHB.v(82)
  // src/AHB.v(82)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg33_b17|U_AHB/reg33_b3  (
    .a({\PWMF/n24 ,\PWMF/n24 }),
    .b({\PWMF/n25_neg_lutinv ,\PWMF/n25_neg_lutinv }),
    .c({\PWMF/n26 [17],\PWMF/n26 [3]}),
    .clk(clk100m),
    .d({\PWMF/pnumr [17],\PWMF/pnumr [3]}),
    .mi({\U_AHB/h2h_hwdata [17],\U_AHB/h2h_hwdata [3]}),
    .sr(\U_AHB/n77 ),
    .f({_al_u2934_o,_al_u2918_o}),
    .q({pnumF[17],pnumF[3]}));  // src/AHB.v(82)
  // src/AHB.v(82)
  // src/AHB.v(82)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg33_b18|U_AHB/reg33_b23  (
    .a({\PWMF/n24 ,\PWMF/n24 }),
    .b({\PWMF/n25_neg_lutinv ,\PWMF/n25_neg_lutinv }),
    .c({\PWMF/n26 [18],\PWMF/n26 [23]}),
    .clk(clk100m),
    .d({\PWMF/pnumr [18],\PWMF/pnumr [23]}),
    .mi({\U_AHB/h2h_hwdata [18],\U_AHB/h2h_hwdata [23]}),
    .sr(\U_AHB/n77 ),
    .f({_al_u2932_o,_al_u2920_o}),
    .q({pnumF[18],pnumF[23]}));  // src/AHB.v(82)
  // src/AHB.v(82)
  // src/AHB.v(82)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg33_b19|U_AHB/reg33_b22  (
    .a({\PWMF/n24 ,\PWMF/n24 }),
    .b({\PWMF/n25_neg_lutinv ,\PWMF/n25_neg_lutinv }),
    .c({\PWMF/n26 [19],\PWMF/n26 [22]}),
    .clk(clk100m),
    .d({\PWMF/pnumr [19],\PWMF/pnumr [22]}),
    .mi({\U_AHB/h2h_hwdata [19],\U_AHB/h2h_hwdata [22]}),
    .sr(\U_AHB/n77 ),
    .f({_al_u2930_o,_al_u2922_o}),
    .q({pnumF[19],pnumF[22]}));  // src/AHB.v(82)
  // src/AHB.v(82)
  // src/AHB.v(82)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg33_b1|U_AHB/reg33_b21  (
    .a({\PWMF/n24 ,\PWMF/n24 }),
    .b({\PWMF/n25_neg_lutinv ,\PWMF/n25_neg_lutinv }),
    .c({\PWMF/n26 [1],\PWMF/n26 [21]}),
    .clk(clk100m),
    .d({\PWMF/pnumr [1],\PWMF/pnumr [21]}),
    .mi({\U_AHB/h2h_hwdata [1],\U_AHB/h2h_hwdata [21]}),
    .sr(\U_AHB/n77 ),
    .f({_al_u2950_o,_al_u2924_o}),
    .q({pnumF[1],pnumF[21]}));  // src/AHB.v(82)
  // src/AHB.v(82)
  // src/AHB.v(82)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg33_b2|U_AHB/reg33_b20  (
    .a({\PWMF/n24 ,\PWMF/n24 }),
    .b({\PWMF/n25_neg_lutinv ,\PWMF/n25_neg_lutinv }),
    .c({\PWMF/n26 [2],\PWMF/n26 [20]}),
    .clk(clk100m),
    .d({\PWMF/pnumr [2],\PWMF/pnumr [20]}),
    .mi({\U_AHB/h2h_hwdata [2],\U_AHB/h2h_hwdata [20]}),
    .sr(\U_AHB/n77 ),
    .f({_al_u2928_o,_al_u2926_o}),
    .q({pnumF[2],pnumF[20]}));  // src/AHB.v(82)
  // src/AHB.v(82)
  // src/AHB.v(82)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg33_b30|U_AHB/reg33_b29  (
    .a({_al_u2821_o,_al_u3095_o}),
    .b({pnumcntE[6],\U_AHB/n90 }),
    .c({pnumcntE[7],\U_AHB/n87 }),
    .clk(clk100m),
    .d({pnumcntE[8],pnumcntD[9]}),
    .e({pnumcntE[9],pnumcntE[9]}),
    .mi(\U_AHB/h2h_hwdata [30:29]),
    .sr(\U_AHB/n77 ),
    .f({_al_u2822_o,_al_u3096_o}),
    .q(pnumF[30:29]));  // src/AHB.v(82)
  // src/AHB.v(82)
  // src/AHB.v(82)
  EF2_PHY_MSLICE #(
    //.LUT0("(~D*~C*~B*~A)"),
    //.LUT1("(~D*~C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000001),
    .INIT_LUT1(16'b0000000000000010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg33_b9|U_AHB/reg33_b26  (
    .a({_al_u1253_o,\PWME/FreCnt [23]}),
    .b({\PWME/FreCnt [7],\PWME/FreCnt [24]}),
    .c({\PWME/FreCnt [8],\PWME/FreCnt [25]}),
    .clk(clk100m),
    .d({\PWME/FreCnt [9],\PWME/FreCnt [26]}),
    .mi({\U_AHB/h2h_hwdata [9],\U_AHB/h2h_hwdata [26]}),
    .sr(\U_AHB/n77 ),
    .f({_al_u1254_o,_al_u1252_o}),
    .q({pnumF[9],pnumF[26]}));  // src/AHB.v(82)
  // src/AHB.v(84)
  // src/AHB.v(84)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~(D*C*B*A))"),
    //.LUTF1("(~0*~(D*C*B*A))"),
    //.LUTG0("(~1*~(D*C*B*A))"),
    //.LUTG1("(~1*~(D*C*B*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111111111111111),
    .INIT_LUTF1(16'b0111111111111111),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg34_b0|U_AHB/reg34_b15  (
    .a({_al_u1688_o,_al_u2901_o}),
    .b({_al_u1690_o,_al_u2903_o}),
    .c({_al_u1691_o,_al_u2904_o}),
    .clk(clk100m),
    .d({pnumcnt0[0],pnumcntF[0]}),
    .e({\PWM0/stopreq ,\PWMF/stopreq }),
    .mi({\U_AHB/h2h_hwdata [0],\U_AHB/h2h_hwdata [15]}),
    .sr(\U_AHB/n79 ),
    .f({_al_u3007_o,_al_u3052_o}),
    .q({pwm_start_stop[0],pwm_start_stop[15]}));  // src/AHB.v(84)
  // src/AHB.v(84)
  // src/AHB.v(84)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~(D*C*B*A))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~1*~(D*C*B*A))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111111111111111),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg34_b13|U_AHB/reg34_b10  (
    .a({open_n32153,_al_u2502_o}),
    .b({_al_u1219_o,_al_u2504_o}),
    .c({_al_u1221_o,_al_u2505_o}),
    .clk(clk100m),
    .d({_al_u1217_o,pnumcntA[0]}),
    .e({open_n32155,\PWMA/stopreq }),
    .mi({\U_AHB/h2h_hwdata [13],\U_AHB/h2h_hwdata [10]}),
    .sr(\U_AHB/n79 ),
    .f({\PWMD/n0_lutinv ,_al_u3037_o}),
    .q({pwm_start_stop[13],pwm_start_stop[10]}));  // src/AHB.v(84)
  // src/AHB.v(84)
  // src/AHB.v(84)
  EF2_PHY_MSLICE #(
    //.LUT0("~(~C*~D)"),
    //.LUT1("(C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg34_b14|U_AHB/reg34_b23  (
    .c({pwm_state_read[14],pwm_start_stop[23]}),
    .clk(clk100m),
    .d({\PWME/n0_lutinv ,pwm_state_read[7]}),
    .mi({\U_AHB/h2h_hwdata [14],\U_AHB/h2h_hwdata [23]}),
    .sr(\U_AHB/n79 ),
    .f({\PWME/n24 ,\PWM7/n11 }),
    .q({pwm_start_stop[14],pwm_start_stop[23]}));  // src/AHB.v(84)
  // src/AHB.v(84)
  // src/AHB.v(84)
  EF2_PHY_MSLICE #(
    //.LUT0("~(~C*~D)"),
    //.LUT1("~(~C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg34_b16|U_AHB/reg34_b20  (
    .c({pwm_start_stop[16],pwm_start_stop[20]}),
    .clk(clk100m),
    .d({pwm_state_read[0],pwm_state_read[4]}),
    .mi({\U_AHB/h2h_hwdata [16],\U_AHB/h2h_hwdata [20]}),
    .sr(\U_AHB/n79 ),
    .f({\PWM0/n11 ,\PWM4/n11 }),
    .q({pwm_start_stop[16],pwm_start_stop[20]}));  // src/AHB.v(84)
  // src/AHB.v(84)
  // src/AHB.v(84)
  EF2_PHY_MSLICE #(
    //.LUT0("~(~C*~D)"),
    //.LUT1("~(~C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg34_b17|U_AHB/reg34_b19  (
    .c({pwm_start_stop[17],pwm_start_stop[19]}),
    .clk(clk100m),
    .d({pwm_state_read[1],pwm_state_read[3]}),
    .mi({\U_AHB/h2h_hwdata [17],\U_AHB/h2h_hwdata [19]}),
    .sr(\U_AHB/n79 ),
    .f({\PWM1/n11 ,\PWM3/n11 }),
    .q({pwm_start_stop[17],pwm_start_stop[19]}));  // src/AHB.v(84)
  // src/AHB.v(84)
  // src/AHB.v(84)
  EF2_PHY_MSLICE #(
    //.LUT0("~(~C*~D)"),
    //.LUT1("~(~C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg34_b21|U_AHB/reg34_b18  (
    .c({pwm_start_stop[21],pwm_start_stop[18]}),
    .clk(clk100m),
    .d({pwm_state_read[5],pwm_state_read[2]}),
    .mi({\U_AHB/h2h_hwdata [21],\U_AHB/h2h_hwdata [18]}),
    .sr(\U_AHB/n79 ),
    .f({\PWM5/n11 ,\PWM2/n11 }),
    .q({pwm_start_stop[21],pwm_start_stop[18]}));  // src/AHB.v(84)
  EF2_PHY_MSLICE #(
    //.LUT0("~(~C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg34_b26  (
    .c({open_n32247,pwm_start_stop[26]}),
    .clk(clk100m),
    .d({open_n32249,pwm_state_read[10]}),
    .mi({open_n32260,\U_AHB/h2h_hwdata [26]}),
    .sr(\U_AHB/n79 ),
    .f({open_n32261,\PWMA/n11 }),
    .q({open_n32265,pwm_start_stop[26]}));  // src/AHB.v(84)
  // src/AHB.v(84)
  // src/AHB.v(84)
  EF2_PHY_MSLICE #(
    //.LUT0("~(~C*~D)"),
    //.LUT1("~(~C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg34_b27|U_AHB/reg34_b31  (
    .c({pwm_start_stop[27],pwm_start_stop[31]}),
    .clk(clk100m),
    .d({pwm_state_read[11],pwm_state_read[15]}),
    .mi({\U_AHB/h2h_hwdata [27],\U_AHB/h2h_hwdata [31]}),
    .sr(\U_AHB/n79 ),
    .f({\PWMB/n11 ,\PWMF/n11 }),
    .q({pwm_start_stop[27],pwm_start_stop[31]}));  // src/AHB.v(84)
  // src/AHB.v(84)
  // src/AHB.v(84)
  EF2_PHY_MSLICE #(
    //.LUT0("~(~C*~D)"),
    //.LUT1("~(~C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1111111111110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg34_b28|U_AHB/reg34_b30  (
    .c({pwm_start_stop[28],pwm_start_stop[30]}),
    .clk(clk100m),
    .d({pwm_state_read[12],pwm_state_read[14]}),
    .mi({\U_AHB/h2h_hwdata [28],\U_AHB/h2h_hwdata [30]}),
    .sr(\U_AHB/n79 ),
    .f({\PWMC/n11 ,\PWME/n11 }),
    .q({pwm_start_stop[28],pwm_start_stop[30]}));  // src/AHB.v(84)
  // src/AHB.v(84)
  // src/AHB.v(84)
  EF2_PHY_MSLICE #(
    //.LUT0("~(~C*~D)"),
    //.LUT1("(C*B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg34_b2|U_AHB/reg34_b29  (
    .b({_al_u812_o,open_n32304}),
    .c({_al_u814_o,pwm_start_stop[29]}),
    .clk(clk100m),
    .d({_al_u810_o,pwm_state_read[13]}),
    .mi({\U_AHB/h2h_hwdata [2],\U_AHB/h2h_hwdata [29]}),
    .sr(\U_AHB/n79 ),
    .f({\PWM2/n0_lutinv ,\PWMD/n11 }),
    .q({pwm_start_stop[2],pwm_start_stop[29]}));  // src/AHB.v(84)
  // src/AHB.v(84)
  // src/AHB.v(84)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(C*B*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg34_b3|U_AHB/reg34_b7  (
    .b({_al_u849_o,_al_u997_o}),
    .c({_al_u851_o,_al_u999_o}),
    .clk(clk100m),
    .d({_al_u847_o,_al_u995_o}),
    .mi({\U_AHB/h2h_hwdata [3],\U_AHB/h2h_hwdata [7]}),
    .sr(\U_AHB/n79 ),
    .f({\PWM3/n0_lutinv ,\PWM7/n0_lutinv }),
    .q({pwm_start_stop[3],pwm_start_stop[7]}));  // src/AHB.v(84)
  // src/AHB.v(84)
  // src/AHB.v(84)
  EF2_PHY_MSLICE #(
    //.LUT0("~(~C*~D)"),
    //.LUT1("(C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg34_b6|U_AHB/reg34_b22  (
    .c({pwm_state_read[6],pwm_start_stop[22]}),
    .clk(clk100m),
    .d({\PWM6/n0_lutinv ,pwm_state_read[6]}),
    .mi({\U_AHB/h2h_hwdata [6],\U_AHB/h2h_hwdata [22]}),
    .sr(\U_AHB/n79 ),
    .f({\PWM6/n24 ,\PWM6/n11 }),
    .q({pwm_start_stop[6],pwm_start_stop[22]}));  // src/AHB.v(84)
  // src/AHB.v(84)
  // src/AHB.v(84)
  EF2_PHY_MSLICE #(
    //.LUT0("~(~C*~D)"),
    //.LUT1("(C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg34_b8|U_AHB/reg34_b24  (
    .c({pwm_state_read[8],pwm_start_stop[24]}),
    .clk(clk100m),
    .d({\PWM8/n0_lutinv ,pwm_state_read[8]}),
    .mi({\U_AHB/h2h_hwdata [8],\U_AHB/h2h_hwdata [24]}),
    .sr(\U_AHB/n79 ),
    .f({\PWM8/n24 ,\PWM8/n11 }),
    .q({pwm_start_stop[8],pwm_start_stop[24]}));  // src/AHB.v(84)
  // src/AHB.v(84)
  // src/AHB.v(84)
  EF2_PHY_MSLICE #(
    //.LUT0("~(~C*~D)"),
    //.LUT1("(C*D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111111111110000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \U_AHB/reg34_b9|U_AHB/reg34_b25  (
    .c({pwm_state_read[9],pwm_start_stop[25]}),
    .clk(clk100m),
    .d({\PWM9/n0_lutinv ,pwm_state_read[9]}),
    .mi({\U_AHB/h2h_hwdata [9],\U_AHB/h2h_hwdata [25]}),
    .sr(\U_AHB/n79 ),
    .f({\PWM9/n24 ,\PWM9/n11 }),
    .q({pwm_start_stop[9],pwm_start_stop[25]}));  // src/AHB.v(84)
  // src/AHB.v(115)
  // src/AHB.v(115)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*C*~(D)*~(0)+~(A)*B*C*~(D)*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0)"),
    //.LUTF1("(~(A)*~(B)*C*~(D)*~(0)+~(A)*B*C*~(D)*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0)"),
    //.LUTG0("(~(A)*~(B)*C*~(D)*~(1)+~(A)*B*C*~(D)*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1)"),
    //.LUTG1("(~(A)*~(B)*C*~(D)*~(1)+~(A)*B*C*~(D)*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011000001010000),
    .INIT_LUTF1(16'b0011000001010000),
    .INIT_LUTG0(16'b0011001101010011),
    .INIT_LUTG1(16'b0011001101010011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg35_b0|U_AHB/reg35_b21  (
    .a({_al_u3348_o,_al_u3194_o}),
    .b({_al_u3352_o,_al_u3198_o}),
    .c({_al_u3061_o,_al_u3061_o}),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [13],\U_AHB/h2h_haddr [13]}),
    .e({\U_AHB/h2h_hrdata [0],\U_AHB/h2h_hrdata [21]}),
    .q({\U_AHB/h2h_hrdata [0],\U_AHB/h2h_hrdata [21]}));  // src/AHB.v(115)
  // src/AHB.v(115)
  // src/AHB.v(115)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*C*~(D)*~(0)+~(A)*B*C*~(D)*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0)"),
    //.LUTF1("(~(A)*~(B)*C*~(D)*~(0)+~(A)*B*C*~(D)*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0)"),
    //.LUTG0("(~(A)*~(B)*C*~(D)*~(1)+~(A)*B*C*~(D)*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1)"),
    //.LUTG1("(~(A)*~(B)*C*~(D)*~(1)+~(A)*B*C*~(D)*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011000001010000),
    .INIT_LUTF1(16'b0011000001010000),
    .INIT_LUTG0(16'b0011001101010011),
    .INIT_LUTG1(16'b0011001101010011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg35_b10|U_AHB/reg35_b20  (
    .a({_al_u3326_o,_al_u3205_o}),
    .b({_al_u3330_o,_al_u3209_o}),
    .c({_al_u3061_o,_al_u3061_o}),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [13],\U_AHB/h2h_haddr [13]}),
    .e({\U_AHB/h2h_hrdata [10],\U_AHB/h2h_hrdata [20]}),
    .q({\U_AHB/h2h_hrdata [10],\U_AHB/h2h_hrdata [20]}));  // src/AHB.v(115)
  // src/AHB.v(115)
  // src/AHB.v(115)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*C*~(D)*~(0)+~(A)*B*C*~(D)*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0)"),
    //.LUTF1("(~(A)*~(B)*C*~(D)*~(0)+~(A)*B*C*~(D)*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0)"),
    //.LUTG0("(~(A)*~(B)*C*~(D)*~(1)+~(A)*B*C*~(D)*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1)"),
    //.LUTG1("(~(A)*~(B)*C*~(D)*~(1)+~(A)*B*C*~(D)*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011000001010000),
    .INIT_LUTF1(16'b0011000001010000),
    .INIT_LUTG0(16'b0011001101010011),
    .INIT_LUTG1(16'b0011001101010011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg35_b11|U_AHB/reg35_b17  (
    .a({_al_u3315_o,_al_u3249_o}),
    .b({_al_u3319_o,_al_u3253_o}),
    .c({_al_u3061_o,_al_u3061_o}),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [13],\U_AHB/h2h_haddr [13]}),
    .e({\U_AHB/h2h_hrdata [11],\U_AHB/h2h_hrdata [17]}),
    .q({\U_AHB/h2h_hrdata [11],\U_AHB/h2h_hrdata [17]}));  // src/AHB.v(115)
  // src/AHB.v(115)
  // src/AHB.v(115)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*C*~(D)*~(0)+~(A)*B*C*~(D)*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0)"),
    //.LUTF1("(~(A)*~(B)*C*~(D)*~(0)+~(A)*B*C*~(D)*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0)"),
    //.LUTG0("(~(A)*~(B)*C*~(D)*~(1)+~(A)*B*C*~(D)*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1)"),
    //.LUTG1("(~(A)*~(B)*C*~(D)*~(1)+~(A)*B*C*~(D)*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011000001010000),
    .INIT_LUTF1(16'b0011000001010000),
    .INIT_LUTG0(16'b0011001101010011),
    .INIT_LUTG1(16'b0011001101010011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg35_b12|U_AHB/reg35_b16  (
    .a({_al_u3304_o,_al_u3260_o}),
    .b({_al_u3308_o,_al_u3264_o}),
    .c({_al_u3061_o,_al_u3061_o}),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [13],\U_AHB/h2h_haddr [13]}),
    .e({\U_AHB/h2h_hrdata [12],\U_AHB/h2h_hrdata [16]}),
    .q({\U_AHB/h2h_hrdata [12],\U_AHB/h2h_hrdata [16]}));  // src/AHB.v(115)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*C*~(D)*~(0)+~(A)*B*C*~(D)*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0)"),
    //.LUT1("(~(A)*~(B)*C*~(D)*~(1)+~(A)*B*C*~(D)*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011000001010000),
    .INIT_LUT1(16'b0011001101010011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg35_b14  (
    .a({_al_u3282_o,_al_u3282_o}),
    .b({_al_u3286_o,_al_u3286_o}),
    .c({_al_u3061_o,_al_u3061_o}),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [13],\U_AHB/h2h_haddr [13]}),
    .mi({open_n32484,\U_AHB/h2h_hrdata [14]}),
    .q({open_n32491,\U_AHB/h2h_hrdata [14]}));  // src/AHB.v(115)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*C*~(D)*~(0)+~(A)*B*C*~(D)*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0)"),
    //.LUT1("(~(A)*~(B)*C*~(D)*~(1)+~(A)*B*C*~(D)*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011000001010000),
    .INIT_LUT1(16'b0011001101010011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg35_b15  (
    .a({_al_u3271_o,_al_u3271_o}),
    .b({_al_u3275_o,_al_u3275_o}),
    .c({_al_u3061_o,_al_u3061_o}),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [13],\U_AHB/h2h_haddr [13]}),
    .mi({open_n32503,\U_AHB/h2h_hrdata [15]}),
    .q({open_n32510,\U_AHB/h2h_hrdata [15]}));  // src/AHB.v(115)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(~(0*~D)*~B)*~(C*A))"),
    //.LUT1("(~(~(1*~D)*~B)*~(C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0100110001001100),
    .INIT_LUT1(16'b0100110001011111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg35_b18  (
    .a({_al_u3237_o,_al_u3237_o}),
    .b({_al_u3241_o,_al_u3241_o}),
    .c({_al_u3242_o,_al_u3242_o}),
    .clk(clk100m),
    .d({_al_u3065_o,_al_u3065_o}),
    .mi({open_n32522,\U_AHB/h2h_hrdata [18]}),
    .q({open_n32529,\U_AHB/h2h_hrdata [18]}));  // src/AHB.v(115)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*C*~(D)*~(0)+~(A)*B*C*~(D)*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0)"),
    //.LUT1("(~(A)*~(B)*C*~(D)*~(1)+~(A)*B*C*~(D)*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011000001010000),
    .INIT_LUT1(16'b0011001101010011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg35_b19  (
    .a({_al_u3227_o,_al_u3227_o}),
    .b({_al_u3231_o,_al_u3231_o}),
    .c({_al_u3061_o,_al_u3061_o}),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [13],\U_AHB/h2h_haddr [13]}),
    .mi({open_n32541,\U_AHB/h2h_hrdata [19]}),
    .q({open_n32548,\U_AHB/h2h_hrdata [19]}));  // src/AHB.v(115)
  // src/AHB.v(115)
  // src/AHB.v(115)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(A)*~(B)*C*~(D)*~(0)+~(A)*B*C*~(D)*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0)"),
    //.LUTF1("(~(A)*~(B)*C*~(D)*~(0)+~(A)*B*C*~(D)*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0)"),
    //.LUTG0("(~(A)*~(B)*C*~(D)*~(1)+~(A)*B*C*~(D)*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1)"),
    //.LUTG1("(~(A)*~(B)*C*~(D)*~(1)+~(A)*B*C*~(D)*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0011000001010000),
    .INIT_LUTF1(16'b0011000001010000),
    .INIT_LUTG0(16'b0011001101010011),
    .INIT_LUTG1(16'b0011001101010011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg35_b1|U_AHB/reg35_b13  (
    .a({_al_u3337_o,_al_u3293_o}),
    .b({_al_u3341_o,_al_u3297_o}),
    .c({_al_u3061_o,_al_u3061_o}),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [13],\U_AHB/h2h_haddr [13]}),
    .e({\U_AHB/h2h_hrdata [1],\U_AHB/h2h_hrdata [13]}),
    .q({\U_AHB/h2h_hrdata [1],\U_AHB/h2h_hrdata [13]}));  // src/AHB.v(115)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*C*~(D)*~(0)+~(A)*B*C*~(D)*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0)"),
    //.LUT1("(~(A)*~(B)*C*~(D)*~(1)+~(A)*B*C*~(D)*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011000001010000),
    .INIT_LUT1(16'b0011001101010011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg35_b2  (
    .a({_al_u3216_o,_al_u3216_o}),
    .b({_al_u3220_o,_al_u3220_o}),
    .c({_al_u3061_o,_al_u3061_o}),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [13],\U_AHB/h2h_haddr [13]}),
    .mi({open_n32581,\U_AHB/h2h_hrdata [2]}),
    .q({open_n32588,\U_AHB/h2h_hrdata [2]}));  // src/AHB.v(115)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*C*~(D)*~(0)+~(A)*B*C*~(D)*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0)"),
    //.LUT1("(~(A)*~(B)*C*~(D)*~(1)+~(A)*B*C*~(D)*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011000001010000),
    .INIT_LUT1(16'b0011001101010011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg35_b22  (
    .a({_al_u3183_o,_al_u3183_o}),
    .b({_al_u3187_o,_al_u3187_o}),
    .c({_al_u3061_o,_al_u3061_o}),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [13],\U_AHB/h2h_haddr [13]}),
    .mi({open_n32600,\U_AHB/h2h_hrdata [22]}),
    .q({open_n32607,\U_AHB/h2h_hrdata [22]}));  // src/AHB.v(115)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*C*~(D)*~(0)+~(A)*B*C*~(D)*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0)"),
    //.LUT1("(~(A)*~(B)*C*~(D)*~(1)+~(A)*B*C*~(D)*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011000001010000),
    .INIT_LUT1(16'b0011001101010011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg35_b23  (
    .a({_al_u3172_o,_al_u3172_o}),
    .b({_al_u3176_o,_al_u3176_o}),
    .c({_al_u3061_o,_al_u3061_o}),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [13],\U_AHB/h2h_haddr [13]}),
    .mi({open_n32619,\U_AHB/h2h_hrdata [23]}),
    .q({open_n32626,\U_AHB/h2h_hrdata [23]}));  // src/AHB.v(115)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+A*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*B*~(C)*~(D)*0+A*B*~(C)*~(D)*0+A*~(B)*C*~(D)*0+A*B*C*~(D)*0+~(A)*B*~(C)*D*0+A*B*~(C)*D*0+A*B*C*D*0)"),
    //.LUT1("(A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+A*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*B*~(C)*~(D)*1+A*B*~(C)*~(D)*1+A*~(B)*C*~(D)*1+A*B*C*~(D)*1+~(A)*B*~(C)*D*1+A*B*~(C)*D*1+A*B*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000010101010),
    .INIT_LUT1(16'b1000110010101111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg35_b24  (
    .a({_al_u3080_o,_al_u3080_o}),
    .b({\U_AHB/n113_lutinv ,\U_AHB/n113_lutinv }),
    .c({_al_u3065_o,_al_u3065_o}),
    .clk(clk100m),
    .d({\U_AHB/n82 ,\U_AHB/n82 }),
    .mi({open_n32638,\U_AHB/h2h_hrdata [24]}),
    .q({open_n32645,\U_AHB/h2h_hrdata [24]}));  // src/AHB.v(115)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+A*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*B*~(C)*~(D)*0+A*B*~(C)*~(D)*0+A*~(B)*C*~(D)*0+A*B*C*~(D)*0+~(A)*B*~(C)*D*0+A*B*~(C)*D*0+A*B*C*D*0)"),
    //.LUT1("(A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+A*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*B*~(C)*~(D)*1+A*B*~(C)*~(D)*1+A*~(B)*C*~(D)*1+A*B*C*~(D)*1+~(A)*B*~(C)*D*1+A*B*~(C)*D*1+A*B*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000010101010),
    .INIT_LUT1(16'b1000110010101111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg35_b25  (
    .a({_al_u3078_o,_al_u3078_o}),
    .b({\U_AHB/n113_lutinv ,\U_AHB/n113_lutinv }),
    .c({_al_u3065_o,_al_u3065_o}),
    .clk(clk100m),
    .d({\U_AHB/n82 ,\U_AHB/n82 }),
    .mi({open_n32657,\U_AHB/h2h_hrdata [25]}),
    .q({open_n32664,\U_AHB/h2h_hrdata [25]}));  // src/AHB.v(115)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+A*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*B*~(C)*~(D)*0+A*B*~(C)*~(D)*0+A*~(B)*C*~(D)*0+A*B*C*~(D)*0+~(A)*B*~(C)*D*0+A*B*~(C)*D*0+A*B*C*D*0)"),
    //.LUT1("(A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+A*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*B*~(C)*~(D)*1+A*B*~(C)*~(D)*1+A*~(B)*C*~(D)*1+A*B*C*~(D)*1+~(A)*B*~(C)*D*1+A*B*~(C)*D*1+A*B*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000010101010),
    .INIT_LUT1(16'b1000110010101111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg35_b26  (
    .a({_al_u3076_o,_al_u3076_o}),
    .b({\U_AHB/n113_lutinv ,\U_AHB/n113_lutinv }),
    .c({_al_u3065_o,_al_u3065_o}),
    .clk(clk100m),
    .d({\U_AHB/n82 ,\U_AHB/n82 }),
    .mi({open_n32676,\U_AHB/h2h_hrdata [26]}),
    .q({open_n32683,\U_AHB/h2h_hrdata [26]}));  // src/AHB.v(115)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+A*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*B*~(C)*~(D)*0+A*B*~(C)*~(D)*0+A*~(B)*C*~(D)*0+A*B*C*~(D)*0+~(A)*B*~(C)*D*0+A*B*~(C)*D*0+A*B*C*D*0)"),
    //.LUT1("(A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+A*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*B*~(C)*~(D)*1+A*B*~(C)*~(D)*1+A*~(B)*C*~(D)*1+A*B*C*~(D)*1+~(A)*B*~(C)*D*1+A*B*~(C)*D*1+A*B*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000010101010),
    .INIT_LUT1(16'b1000110010101111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg35_b27  (
    .a({_al_u3074_o,_al_u3074_o}),
    .b({\U_AHB/n113_lutinv ,\U_AHB/n113_lutinv }),
    .c({_al_u3065_o,_al_u3065_o}),
    .clk(clk100m),
    .d({\U_AHB/n82 ,\U_AHB/n82 }),
    .mi({open_n32695,\U_AHB/h2h_hrdata [27]}),
    .q({open_n32702,\U_AHB/h2h_hrdata [27]}));  // src/AHB.v(115)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+A*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*B*~(C)*~(D)*0+A*B*~(C)*~(D)*0+A*~(B)*C*~(D)*0+A*B*C*~(D)*0+~(A)*B*~(C)*D*0+A*B*~(C)*D*0+A*B*C*D*0)"),
    //.LUT1("(A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+A*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*B*~(C)*~(D)*1+A*B*~(C)*~(D)*1+A*~(B)*C*~(D)*1+A*B*C*~(D)*1+~(A)*B*~(C)*D*1+A*B*~(C)*D*1+A*B*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000010101010),
    .INIT_LUT1(16'b1000110010101111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg35_b28  (
    .a({_al_u3072_o,_al_u3072_o}),
    .b({\U_AHB/n113_lutinv ,\U_AHB/n113_lutinv }),
    .c({_al_u3065_o,_al_u3065_o}),
    .clk(clk100m),
    .d({\U_AHB/n82 ,\U_AHB/n82 }),
    .mi({open_n32714,\U_AHB/h2h_hrdata [28]}),
    .q({open_n32721,\U_AHB/h2h_hrdata [28]}));  // src/AHB.v(115)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+A*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*B*~(C)*~(D)*0+A*B*~(C)*~(D)*0+A*~(B)*C*~(D)*0+A*B*C*~(D)*0+~(A)*B*~(C)*D*0+A*B*~(C)*D*0+A*B*C*D*0)"),
    //.LUT1("(A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+A*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*B*~(C)*~(D)*1+A*B*~(C)*~(D)*1+A*~(B)*C*~(D)*1+A*B*C*~(D)*1+~(A)*B*~(C)*D*1+A*B*~(C)*D*1+A*B*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000010101010),
    .INIT_LUT1(16'b1000110010101111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg35_b29  (
    .a({_al_u3070_o,_al_u3070_o}),
    .b({\U_AHB/n113_lutinv ,\U_AHB/n113_lutinv }),
    .c({_al_u3065_o,_al_u3065_o}),
    .clk(clk100m),
    .d({\U_AHB/n82 ,\U_AHB/n82 }),
    .mi({open_n32733,\U_AHB/h2h_hrdata [29]}),
    .q({open_n32740,\U_AHB/h2h_hrdata [29]}));  // src/AHB.v(115)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*C*~(D)*~(0)+~(A)*B*C*~(D)*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0)"),
    //.LUT1("(~(A)*~(B)*C*~(D)*~(1)+~(A)*B*C*~(D)*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011000001010000),
    .INIT_LUT1(16'b0011001101010011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg35_b3  (
    .a({_al_u3161_o,_al_u3161_o}),
    .b({_al_u3165_o,_al_u3165_o}),
    .c({_al_u3061_o,_al_u3061_o}),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [13],\U_AHB/h2h_haddr [13]}),
    .mi({open_n32752,\U_AHB/h2h_hrdata [3]}),
    .q({open_n32759,\U_AHB/h2h_hrdata [3]}));  // src/AHB.v(115)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+A*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*B*~(C)*~(D)*0+A*B*~(C)*~(D)*0+A*~(B)*C*~(D)*0+A*B*C*~(D)*0+~(A)*B*~(C)*D*0+A*B*~(C)*D*0+A*B*C*D*0)"),
    //.LUT1("(A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+A*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*B*~(C)*~(D)*1+A*B*~(C)*~(D)*1+A*~(B)*C*~(D)*1+A*B*C*~(D)*1+~(A)*B*~(C)*D*1+A*B*~(C)*D*1+A*B*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000010101010),
    .INIT_LUT1(16'b1000110010101111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg35_b30  (
    .a({_al_u3068_o,_al_u3068_o}),
    .b({\U_AHB/n113_lutinv ,\U_AHB/n113_lutinv }),
    .c({_al_u3065_o,_al_u3065_o}),
    .clk(clk100m),
    .d({\U_AHB/n82 ,\U_AHB/n82 }),
    .mi({open_n32771,\U_AHB/h2h_hrdata [30]}),
    .q({open_n32778,\U_AHB/h2h_hrdata [30]}));  // src/AHB.v(115)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*~(B)*~(C)*~(D)*~(0)+A*B*~(C)*~(D)*~(0)+A*~(B)*C*~(D)*~(0)+A*B*C*~(D)*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*B*~(C)*~(D)*0+A*B*~(C)*~(D)*0+A*~(B)*C*~(D)*0+A*B*C*~(D)*0+~(A)*B*~(C)*D*0+A*B*~(C)*D*0+A*B*C*D*0)"),
    //.LUT1("(A*~(B)*~(C)*~(D)*~(1)+A*B*~(C)*~(D)*~(1)+A*~(B)*C*~(D)*~(1)+A*B*C*~(D)*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*B*~(C)*~(D)*1+A*B*~(C)*~(D)*1+A*~(B)*C*~(D)*1+A*B*C*~(D)*1+~(A)*B*~(C)*D*1+A*B*~(C)*D*1+A*B*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000010101010),
    .INIT_LUT1(16'b1000110010101111),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg35_b31  (
    .a({_al_u3062_o,_al_u3062_o}),
    .b({\U_AHB/n113_lutinv ,\U_AHB/n113_lutinv }),
    .c({_al_u3065_o,_al_u3065_o}),
    .clk(clk100m),
    .d({\U_AHB/n82 ,\U_AHB/n82 }),
    .mi({open_n32790,\U_AHB/h2h_hrdata [31]}),
    .q({open_n32797,\U_AHB/h2h_hrdata [31]}));  // src/AHB.v(115)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*C*~(D)*~(0)+~(A)*B*C*~(D)*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0)"),
    //.LUT1("(~(A)*~(B)*C*~(D)*~(1)+~(A)*B*C*~(D)*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011000001010000),
    .INIT_LUT1(16'b0011001101010011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg35_b4  (
    .a({_al_u3150_o,_al_u3150_o}),
    .b({_al_u3154_o,_al_u3154_o}),
    .c({_al_u3061_o,_al_u3061_o}),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [13],\U_AHB/h2h_haddr [13]}),
    .mi({open_n32809,\U_AHB/h2h_hrdata [4]}),
    .q({open_n32816,\U_AHB/h2h_hrdata [4]}));  // src/AHB.v(115)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*C*~(D)*~(0)+~(A)*B*C*~(D)*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0)"),
    //.LUT1("(~(A)*~(B)*C*~(D)*~(1)+~(A)*B*C*~(D)*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011000001010000),
    .INIT_LUT1(16'b0011001101010011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg35_b5  (
    .a({_al_u3138_o,_al_u3138_o}),
    .b({_al_u3143_o,_al_u3143_o}),
    .c({_al_u3061_o,_al_u3061_o}),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [13],\U_AHB/h2h_haddr [13]}),
    .mi({open_n32828,\U_AHB/h2h_hrdata [5]}),
    .q({open_n32835,\U_AHB/h2h_hrdata [5]}));  // src/AHB.v(115)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*C*~(D)*~(0)+~(A)*B*C*~(D)*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0)"),
    //.LUT1("(~(A)*~(B)*C*~(D)*~(1)+~(A)*B*C*~(D)*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011000001010000),
    .INIT_LUT1(16'b0011001101010011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg35_b6  (
    .a({_al_u3127_o,_al_u3127_o}),
    .b({_al_u3131_o,_al_u3131_o}),
    .c({_al_u3061_o,_al_u3061_o}),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [13],\U_AHB/h2h_haddr [13]}),
    .mi({open_n32847,\U_AHB/h2h_hrdata [6]}),
    .q({open_n32854,\U_AHB/h2h_hrdata [6]}));  // src/AHB.v(115)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*C*~(D)*~(0)+~(A)*B*C*~(D)*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0)"),
    //.LUT1("(~(A)*~(B)*C*~(D)*~(1)+~(A)*B*C*~(D)*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011000001010000),
    .INIT_LUT1(16'b0011001101010011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg35_b7  (
    .a({_al_u3116_o,_al_u3116_o}),
    .b({_al_u3120_o,_al_u3120_o}),
    .c({_al_u3061_o,_al_u3061_o}),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [13],\U_AHB/h2h_haddr [13]}),
    .mi({open_n32866,\U_AHB/h2h_hrdata [7]}),
    .q({open_n32873,\U_AHB/h2h_hrdata [7]}));  // src/AHB.v(115)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*C*~(D)*~(0)+~(A)*B*C*~(D)*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0)"),
    //.LUT1("(~(A)*~(B)*C*~(D)*~(1)+~(A)*B*C*~(D)*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011000001010000),
    .INIT_LUT1(16'b0011001101010011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg35_b8  (
    .a({_al_u3105_o,_al_u3105_o}),
    .b({_al_u3109_o,_al_u3109_o}),
    .c({_al_u3061_o,_al_u3061_o}),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [13],\U_AHB/h2h_haddr [13]}),
    .mi({open_n32885,\U_AHB/h2h_hrdata [8]}),
    .q({open_n32892,\U_AHB/h2h_hrdata [8]}));  // src/AHB.v(115)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*C*~(D)*~(0)+~(A)*B*C*~(D)*~(0)+~(A)*~(B)*C*D*~(0)+A*~(B)*C*D*~(0)+~(A)*~(B)*~(C)*~(D)*0+A*~(B)*~(C)*~(D)*0+~(A)*~(B)*C*~(D)*0+~(A)*B*C*~(D)*0+~(A)*~(B)*~(C)*D*0+A*~(B)*~(C)*D*0+~(A)*~(B)*C*D*0+A*~(B)*C*D*0)"),
    //.LUT1("(~(A)*~(B)*C*~(D)*~(1)+~(A)*B*C*~(D)*~(1)+~(A)*~(B)*C*D*~(1)+A*~(B)*C*D*~(1)+~(A)*~(B)*~(C)*~(D)*1+A*~(B)*~(C)*~(D)*1+~(A)*~(B)*C*~(D)*1+~(A)*B*C*~(D)*1+~(A)*~(B)*~(C)*D*1+A*~(B)*~(C)*D*1+~(A)*~(B)*C*D*1+A*~(B)*C*D*1)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011000001010000),
    .INIT_LUT1(16'b0011001101010011),
    .MODE("LOGIC"),
    .MSFXMUX("ON"),
    .REG0_REGSET("RESET"),
    .REG0_SD("FX"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg35_b9  (
    .a({_al_u3094_o,_al_u3094_o}),
    .b({_al_u3098_o,_al_u3098_o}),
    .c({_al_u3061_o,_al_u3061_o}),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [13],\U_AHB/h2h_haddr [13]}),
    .mi({open_n32904,\U_AHB/h2h_hrdata [9]}),
    .q({open_n32911,\U_AHB/h2h_hrdata [9]}));  // src/AHB.v(115)
  // src/AHB.v(48)
  // src/AHB.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(~D*~C*B*A)"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(~D*~C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b0000000000001000),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b0000000000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg3_b0|U_AHB/reg3_b20  (
    .a({\U_AHB/h2h_hwrite ,_al_u1408_o}),
    .b({\U_AHB/h2h_haddr [2],\PWM2/FreCnt [20]}),
    .c({\U_AHB/h2h_haddr [13],\PWM2/FreCnt [26]}),
    .ce(\U_AHB/n8 ),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [14],\PWM2/FreCntr [20]}),
    .e({open_n32912,\PWM2/FreCntr [26]}),
    .mi({\U_AHB/h2h_hwdata [0],\U_AHB/h2h_hwdata [20]}),
    .f({\U_AHB/n8 ,_al_u1409_o}),
    .q({freq2[0],freq2[20]}));  // src/AHB.v(48)
  // src/AHB.v(48)
  // src/AHB.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(B*A*~(~D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1000100000001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg3_b11|U_AHB/reg3_b10  (
    .a({_al_u1906_o,open_n32929}),
    .b({_al_u1907_o,open_n32930}),
    .c({\PWM2/FreCnt [10],pwm_state_read[2]}),
    .ce(\U_AHB/n8 ),
    .clk(clk100m),
    .d({\PWM2/FreCntr [11],\PWM2/n0_lutinv }),
    .mi(\U_AHB/h2h_hwdata [11:10]),
    .f({_al_u1908_o,\PWM2/n24 }),
    .q(freq2[11:10]));  // src/AHB.v(48)
  // src/AHB.v(48)
  // src/AHB.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~D*C*B*A)"),
    //.LUTF1("(~(D*~B)*~(C*~A))"),
    //.LUTG0("(~D*C*B*A)"),
    //.LUTG1("(~(D*~B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b1000110010101111),
    .INIT_LUTG0(16'b0000000010000000),
    .INIT_LUTG1(16'b1000110010101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg3_b12|U_AHB/reg3_b24  (
    .a({\PWM2/FreCnt [12],_al_u2581_o}),
    .b({\PWM2/FreCnt [15],_al_u2583_o}),
    .c({\PWM2/FreCntr [12],_al_u2584_o}),
    .ce(\U_AHB/n8 ),
    .clk(clk100m),
    .d({\PWM2/FreCntr [15],pnumcntB[0]}),
    .mi({\U_AHB/h2h_hwdata [12],\U_AHB/h2h_hwdata [24]}),
    .f({_al_u1401_o,\PWMB/n25_neg_lutinv }),
    .q({freq2[12],freq2[24]}));  // src/AHB.v(48)
  // src/AHB.v(48)
  // src/AHB.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b1000010000100001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg3_b13|U_AHB/reg3_b14  (
    .a({\PWM2/FreCnt [13],open_n32963}),
    .b({\PWM2/FreCnt [16],limit_r_pad[2]}),
    .c({\PWM2/FreCntr [13],limit_l_pad[2]}),
    .ce(\U_AHB/n8 ),
    .clk(clk100m),
    .d({\PWM2/FreCntr [16],\PWM2/n11 }),
    .mi({\U_AHB/h2h_hwdata [13],\U_AHB/h2h_hwdata [14]}),
    .f({_al_u1410_o,_al_u3014_o}),
    .q({freq2[13],freq2[14]}));  // src/AHB.v(48)
  // src/AHB.v(48)
  // src/AHB.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(D@B)*~(C@A))"),
    //.LUT1("(C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000010000100001),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg3_b16|U_AHB/reg3_b18  (
    .a({open_n32978,\PWM2/FreCnt [18]}),
    .b({open_n32979,\PWM2/FreCnt [5]}),
    .c({\PWM2/FreCntr [16],\PWM2/FreCntr [18]}),
    .ce(\U_AHB/n8 ),
    .clk(clk100m),
    .d({\PWM2/FreCnt [15],\PWM2/FreCntr [5]}),
    .mi({\U_AHB/h2h_hwdata [16],\U_AHB/h2h_hwdata [18]}),
    .f({_al_u1913_o,_al_u1399_o}),
    .q({freq2[16],freq2[18]}));  // src/AHB.v(48)
  // src/AHB.v(48)
  // src/AHB.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg3_b19|U_AHB/reg3_b22  (
    .a({\PWM2/FreCnt [16],_al_u813_o}),
    .b({\PWM2/FreCnt [17],\PWM2/FreCnt [2]}),
    .c({\PWM2/FreCnt [18],\PWM2/FreCnt [20]}),
    .ce(\U_AHB/n8 ),
    .clk(clk100m),
    .d({\PWM2/FreCnt [19],\PWM2/FreCnt [21]}),
    .e({open_n32994,\PWM2/FreCnt [22]}),
    .mi({\U_AHB/h2h_hwdata [19],\U_AHB/h2h_hwdata [22]}),
    .f({_al_u813_o,_al_u814_o}),
    .q({freq2[19],freq2[22]}));  // src/AHB.v(48)
  // src/AHB.v(48)
  // src/AHB.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg3_b23|U_AHB/reg3_b3  (
    .a({\PWM2/FreCnt [23],_al_u808_o}),
    .b({\PWM2/FreCnt [24],\PWM2/FreCnt [3]}),
    .c({\PWM2/FreCnt [25],\PWM2/FreCnt [4]}),
    .ce(\U_AHB/n8 ),
    .clk(clk100m),
    .d({\PWM2/FreCnt [26],\PWM2/FreCnt [5]}),
    .e({open_n33011,\PWM2/FreCnt [6]}),
    .mi({\U_AHB/h2h_hwdata [23],\U_AHB/h2h_hwdata [3]}),
    .f({_al_u808_o,_al_u809_o}),
    .q({freq2[23],freq2[3]}));  // src/AHB.v(48)
  // src/AHB.v(48)
  // src/AHB.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(C*B*A*~(0@D))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(C*B*A*~(1@D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg3_b4|U_AHB/reg3_b9  (
    .a({_al_u1396_o,_al_u1397_o}),
    .b({_al_u1398_o,\PWM2/FreCnt [11]}),
    .c({_al_u1399_o,\PWM2/FreCnt [9]}),
    .ce(\U_AHB/n8 ),
    .clk(clk100m),
    .d({\PWM2/FreCnt [4],\PWM2/FreCntr [11]}),
    .e({\PWM2/FreCntr [4],\PWM2/FreCntr [9]}),
    .mi({\U_AHB/h2h_hwdata [4],\U_AHB/h2h_hwdata [9]}),
    .f({_al_u1400_o,_al_u1398_o}),
    .q({freq2[4],freq2[9]}));  // src/AHB.v(48)
  // src/AHB.v(48)
  // src/AHB.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(~D*~C*~B*A)"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(~D*~C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b0000000000000010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg3_b7|U_AHB/reg3_b17  (
    .a({_al_u809_o,_al_u1395_o}),
    .b({\PWM2/FreCnt [7],\PWM2/FreCnt [17]}),
    .c({\PWM2/FreCnt [8],\PWM2/FreCnt [8]}),
    .ce(\U_AHB/n8 ),
    .clk(clk100m),
    .d({\PWM2/FreCnt [9],\PWM2/FreCntr [17]}),
    .e({open_n33044,\PWM2/FreCntr [8]}),
    .mi({\U_AHB/h2h_hwdata [7],\U_AHB/h2h_hwdata [17]}),
    .f({_al_u810_o,_al_u1396_o}),
    .q({freq2[7],freq2[17]}));  // src/AHB.v(48)
  // src/AHB.v(49)
  // src/AHB.v(49)
  EF2_PHY_MSLICE #(
    //.LUT0("(~D*~C*B*A)"),
    //.LUT1("(C*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000001000),
    .INIT_LUT1(16'b1111000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg4_b10|U_AHB/reg4_b0  (
    .a({open_n33061,\U_AHB/h2h_hwrite }),
    .b({open_n33062,\U_AHB/h2h_haddr [3]}),
    .c({pwm_state_read[3],\U_AHB/h2h_haddr [13]}),
    .ce(\U_AHB/n10 ),
    .clk(clk100m),
    .d({\PWM3/n0_lutinv ,\U_AHB/h2h_haddr [14]}),
    .mi({\U_AHB/h2h_hwdata [10],\U_AHB/h2h_hwdata [0]}),
    .f({\PWM3/n24 ,\U_AHB/n10 }),
    .q({freq3[10],freq3[0]}));  // src/AHB.v(49)
  // src/AHB.v(49)
  // src/AHB.v(49)
  EF2_PHY_MSLICE #(
    //.LUT0("(~D*C*B*A)"),
    //.LUT1("(~(~D*B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000010000000),
    .INIT_LUT1(16'b1111010100110001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg4_b12|U_AHB/reg4_b5  (
    .a({\PWM3/FreCnt [12],_al_u1770_o}),
    .b({\PWM3/FreCnt [15],_al_u1772_o}),
    .c({\PWM3/FreCntr [12],_al_u1773_o}),
    .ce(\U_AHB/n10 ),
    .clk(clk100m),
    .d({\PWM3/FreCntr [15],pnumcnt1[0]}),
    .mi({\U_AHB/h2h_hwdata [12],\U_AHB/h2h_hwdata [5]}),
    .f({_al_u1423_o,\PWM1/n25_neg_lutinv }),
    .q({freq3[12],freq3[5]}));  // src/AHB.v(49)
  // src/AHB.v(49)
  // src/AHB.v(49)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(C*B*A*~(0@D))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(C*B*A*~(1@D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg4_b14|U_AHB/reg4_b17  (
    .a({_al_u1414_o,_al_u1415_o}),
    .b({_al_u1416_o,\PWM3/FreCnt [17]}),
    .c({_al_u1417_o,\PWM3/FreCnt [8]}),
    .ce(\U_AHB/n10 ),
    .clk(clk100m),
    .d({\PWM3/FreCnt [14],\PWM3/FreCntr [17]}),
    .e({\PWM3/FreCntr [14],\PWM3/FreCntr [8]}),
    .mi({\U_AHB/h2h_hwdata [14],\U_AHB/h2h_hwdata [17]}),
    .f({_al_u1418_o,_al_u1416_o}),
    .q({freq3[14],freq3[17]}));  // src/AHB.v(49)
  // src/AHB.v(49)
  // src/AHB.v(49)
  EF2_PHY_MSLICE #(
    //.LUT0("(~D*C*B*A)"),
    //.LUT1("(~(D*~B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000010000000),
    .INIT_LUT1(16'b1000110010101111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg4_b15|U_AHB/reg4_b25  (
    .a({\PWM3/FreCnt [12],_al_u1688_o}),
    .b({\PWM3/FreCnt [15],_al_u1690_o}),
    .c({\PWM3/FreCntr [12],_al_u1691_o}),
    .ce(\U_AHB/n10 ),
    .clk(clk100m),
    .d({\PWM3/FreCntr [15],pnumcnt0[0]}),
    .mi({\U_AHB/h2h_hwdata [15],\U_AHB/h2h_hwdata [25]}),
    .f({_al_u1419_o,\PWM0/n25_neg_lutinv }),
    .q({freq3[15],freq3[25]}));  // src/AHB.v(49)
  // src/AHB.v(49)
  // src/AHB.v(49)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg4_b16|U_AHB/reg4_b18  (
    .a({\PWM3/FreCnt [16],_al_u1413_o}),
    .b({\PWM3/FreCnt [3],\PWM3/FreCnt [18]}),
    .c({\PWM3/FreCntr [16],\PWM3/FreCnt [5]}),
    .ce(\U_AHB/n10 ),
    .clk(clk100m),
    .d({\PWM3/FreCntr [3],\PWM3/FreCntr [18]}),
    .e({open_n33121,\PWM3/FreCntr [5]}),
    .mi({\U_AHB/h2h_hwdata [16],\U_AHB/h2h_hwdata [18]}),
    .f({_al_u1413_o,_al_u1414_o}),
    .q({freq3[16],freq3[18]}));  // src/AHB.v(49)
  // src/AHB.v(49)
  // src/AHB.v(49)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(C*B*A*~(0@D))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(C*B*A*~(1@D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg4_b21|U_AHB/reg4_b19  (
    .a({_al_u1420_o,_al_u1421_o}),
    .b({_al_u1422_o,\PWM3/FreCnt [13]}),
    .c({_al_u1423_o,\PWM3/FreCnt [19]}),
    .ce(\U_AHB/n10 ),
    .clk(clk100m),
    .d({\PWM3/FreCnt [21],\PWM3/FreCntr [13]}),
    .e({\PWM3/FreCntr [21],\PWM3/FreCntr [19]}),
    .mi({\U_AHB/h2h_hwdata [21],\U_AHB/h2h_hwdata [19]}),
    .f({_al_u1424_o,_al_u1422_o}),
    .q({freq3[21],freq3[19]}));  // src/AHB.v(49)
  // src/AHB.v(49)
  // src/AHB.v(49)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg4_b23|U_AHB/reg4_b3  (
    .a({\PWM3/FreCnt [23],_al_u845_o}),
    .b({\PWM3/FreCnt [24],\PWM3/FreCnt [3]}),
    .c({\PWM3/FreCnt [25],\PWM3/FreCnt [4]}),
    .ce(\U_AHB/n10 ),
    .clk(clk100m),
    .d({\PWM3/FreCnt [26],\PWM3/FreCnt [5]}),
    .e({open_n33154,\PWM3/FreCnt [6]}),
    .mi({\U_AHB/h2h_hwdata [23],\U_AHB/h2h_hwdata [3]}),
    .f({_al_u845_o,_al_u846_o}),
    .q({freq3[23],freq3[3]}));  // src/AHB.v(49)
  // src/AHB.v(49)
  // src/AHB.v(49)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg4_b7|U_AHB/reg4_b11  (
    .a({\PWM3/FreCnt [7],_al_u1425_o}),
    .b({\PWM3/FreCnt [9],\PWM3/FreCnt [11]}),
    .c({\PWM3/FreCntr [7],\PWM3/FreCnt [4]}),
    .ce(\U_AHB/n10 ),
    .clk(clk100m),
    .d({\PWM3/FreCntr [9],\PWM3/FreCntr [11]}),
    .e({open_n33171,\PWM3/FreCntr [4]}),
    .mi({\U_AHB/h2h_hwdata [7],\U_AHB/h2h_hwdata [11]}),
    .f({_al_u1425_o,_al_u1426_o}),
    .q({freq3[7],freq3[11]}));  // src/AHB.v(49)
  // src/AHB.v(49)
  // src/AHB.v(49)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(~D*~C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b0000000000000010),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg4_b8|U_AHB/reg4_b20  (
    .a({_al_u846_o,open_n33188}),
    .b({\PWM3/FreCnt [7],limit_r_pad[3]}),
    .c({\PWM3/FreCnt [8],limit_l_pad[3]}),
    .ce(\U_AHB/n10 ),
    .clk(clk100m),
    .d({\PWM3/FreCnt [9],\PWM3/n11 }),
    .mi({\U_AHB/h2h_hwdata [8],\U_AHB/h2h_hwdata [20]}),
    .f({_al_u847_o,_al_u3017_o}),
    .q({freq3[8],freq3[20]}));  // src/AHB.v(49)
  // src/AHB.v(50)
  // src/AHB.v(50)
  EF2_PHY_MSLICE #(
    //.LUT0("(D*~C*~B*A)"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg5_b10|U_AHB/reg5_b0  (
    .a({open_n33203,\U_AHB/h2h_hwrite }),
    .b({limit_r_pad[4],\U_AHB/h2h_haddr [13]}),
    .c({limit_l_pad[4],\U_AHB/h2h_haddr [14]}),
    .ce(\U_AHB/n12 ),
    .clk(clk100m),
    .d({\PWM4/n11 ,\U_AHB/h2h_haddr [4]}),
    .mi({\U_AHB/h2h_hwdata [10],\U_AHB/h2h_hwdata [0]}),
    .f({_al_u3020_o,\U_AHB/n12 }),
    .q({freq4[10],freq4[0]}));  // src/AHB.v(50)
  // src/AHB.v(50)
  // src/AHB.v(50)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~(~D*B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111010100110001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg5_b12|U_AHB/reg5_b1  (
    .a({\PWM4/FreCnt [12],open_n33218}),
    .b({\PWM4/FreCnt [15],open_n33219}),
    .c({\PWM4/FreCntr [12],pwm_state_read[4]}),
    .ce(\U_AHB/n12 ),
    .clk(clk100m),
    .d({\PWM4/FreCntr [15],\PWM4/n0_lutinv }),
    .mi({\U_AHB/h2h_hwdata [12],\U_AHB/h2h_hwdata [1]}),
    .f({_al_u1440_o,\PWM4/n24 }),
    .q({freq4[12],freq4[1]}));  // src/AHB.v(50)
  // src/AHB.v(50)
  // src/AHB.v(50)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(D*~B)*~(C*~A))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(~(D*~B)*~(C*~A))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000110010101111),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000110010101111),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg5_b16|U_AHB/reg5_b18  (
    .a({\PWM4/FreCnt [16],\PWM4/FreCnt [17]}),
    .b({\PWM4/FreCnt [4],\PWM4/FreCnt [19]}),
    .c({\PWM4/FreCntr [16],\PWM4/FreCntr [18]}),
    .ce(\U_AHB/n12 ),
    .clk(clk100m),
    .d({\PWM4/FreCntr [4],\PWM4/FreCntr [20]}),
    .mi({\U_AHB/h2h_hwdata [16],\U_AHB/h2h_hwdata [18]}),
    .f({_al_u1430_o,_al_u2069_o}),
    .q({freq4[16],freq4[18]}));  // src/AHB.v(50)
  // src/AHB.v(50)
  // src/AHB.v(50)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg5_b17|U_AHB/reg5_b22  (
    .a({\PWM4/FreCnt [16],_al_u887_o}),
    .b({\PWM4/FreCnt [17],\PWM4/FreCnt [2]}),
    .c({\PWM4/FreCnt [18],\PWM4/FreCnt [20]}),
    .ce(\U_AHB/n12 ),
    .clk(clk100m),
    .d({\PWM4/FreCnt [19],\PWM4/FreCnt [21]}),
    .e({open_n33252,\PWM4/FreCnt [22]}),
    .mi({\U_AHB/h2h_hwdata [17],\U_AHB/h2h_hwdata [22]}),
    .f({_al_u887_o,_al_u888_o}),
    .q({freq4[17],freq4[22]}));  // src/AHB.v(50)
  // src/AHB.v(50)
  // src/AHB.v(50)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*B*A*~(0@D))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(C*B*A*~(1@D))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg5_b20|U_AHB/reg5_b14  (
    .a({\PWM4/FreCnt [20],_al_u1431_o}),
    .b({\PWM4/FreCnt [26],_al_u1433_o}),
    .c({\PWM4/FreCntr [20],_al_u1434_o}),
    .ce(\U_AHB/n12 ),
    .clk(clk100m),
    .d({\PWM4/FreCntr [26],\PWM4/FreCnt [14]}),
    .e({open_n33269,\PWM4/FreCntr [14]}),
    .mi({\U_AHB/h2h_hwdata [20],\U_AHB/h2h_hwdata [14]}),
    .f({_al_u1434_o,_al_u1435_o}),
    .q({freq4[20],freq4[14]}));  // src/AHB.v(50)
  // src/AHB.v(50)
  // src/AHB.v(50)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(C*B*A*~(0@D))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(C*B*A*~(1@D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg5_b21|U_AHB/reg5_b19  (
    .a({_al_u1437_o,_al_u1438_o}),
    .b({_al_u1439_o,\PWM4/FreCnt [13]}),
    .c({_al_u1440_o,\PWM4/FreCnt [19]}),
    .ce(\U_AHB/n12 ),
    .clk(clk100m),
    .d({\PWM4/FreCnt [21],\PWM4/FreCntr [13]}),
    .e({\PWM4/FreCntr [21],\PWM4/FreCntr [19]}),
    .mi({\U_AHB/h2h_hwdata [21],\U_AHB/h2h_hwdata [19]}),
    .f({_al_u1441_o,_al_u1439_o}),
    .q({freq4[21],freq4[19]}));  // src/AHB.v(50)
  // src/AHB.v(50)
  // src/AHB.v(50)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg5_b23|U_AHB/reg5_b3  (
    .a({\PWM4/FreCnt [23],_al_u882_o}),
    .b({\PWM4/FreCnt [24],\PWM4/FreCnt [3]}),
    .c({\PWM4/FreCnt [25],\PWM4/FreCnt [4]}),
    .ce(\U_AHB/n12 ),
    .clk(clk100m),
    .d({\PWM4/FreCnt [26],\PWM4/FreCnt [5]}),
    .e({open_n33302,\PWM4/FreCnt [6]}),
    .mi({\U_AHB/h2h_hwdata [23],\U_AHB/h2h_hwdata [3]}),
    .f({_al_u882_o,_al_u883_o}),
    .q({freq4[23],freq4[3]}));  // src/AHB.v(50)
  // src/AHB.v(50)
  // src/AHB.v(50)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(D*~B)*~(C*~A))"),
    //.LUTF1("(D*~(C@B))"),
    //.LUTG0("(~(D*~B)*~(C*~A))"),
    //.LUTG1("(D*~(C@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000110010101111),
    .INIT_LUTF1(16'b1100001100000000),
    .INIT_LUTG0(16'b1000110010101111),
    .INIT_LUTG1(16'b1100001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg5_b6|U_AHB/reg5_b15  (
    .a({open_n33319,\PWM4/FreCnt [12]}),
    .b({\PWM4/FreCnt [6],\PWM4/FreCnt [15]}),
    .c({\PWM4/FreCntr [6],\PWM4/FreCntr [12]}),
    .ce(\U_AHB/n12 ),
    .clk(clk100m),
    .d({_al_u1436_o,\PWM4/FreCntr [15]}),
    .mi({\U_AHB/h2h_hwdata [6],\U_AHB/h2h_hwdata [15]}),
    .f({_al_u1437_o,_al_u1436_o}),
    .q({freq4[6],freq4[15]}));  // src/AHB.v(50)
  // src/AHB.v(50)
  // src/AHB.v(50)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg5_b7|U_AHB/reg5_b11  (
    .a({\PWM4/FreCnt [7],_al_u1442_o}),
    .b({\PWM4/FreCnt [9],\PWM4/FreCnt [11]}),
    .c({\PWM4/FreCntr [7],\PWM4/FreCnt [25]}),
    .ce(\U_AHB/n12 ),
    .clk(clk100m),
    .d({\PWM4/FreCntr [9],\PWM4/FreCntr [11]}),
    .e({open_n33338,\PWM4/FreCntr [25]}),
    .mi({\U_AHB/h2h_hwdata [7],\U_AHB/h2h_hwdata [11]}),
    .f({_al_u1442_o,_al_u1443_o}),
    .q({freq4[7],freq4[11]}));  // src/AHB.v(50)
  // src/AHB.v(51)
  // src/AHB.v(51)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(D*~C*~B*A)"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(D*~C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b0000001000000000),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b0000001000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg6_b0|U_AHB/reg6_b1  (
    .a({\U_AHB/h2h_hwrite ,_al_u1461_o}),
    .b({\U_AHB/h2h_haddr [13],\PWM5/FreCnt [1]}),
    .c({\U_AHB/h2h_haddr [14],\PWM5/FreCnt [10]}),
    .ce(\U_AHB/n14 ),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [5],\PWM5/FreCntr [1]}),
    .e({open_n33355,\PWM5/FreCntr [10]}),
    .mi({\U_AHB/h2h_hwdata [0],\U_AHB/h2h_hwdata [1]}),
    .f({\U_AHB/n14 ,_al_u1462_o}),
    .q({freq5[0],freq5[1]}));  // src/AHB.v(51)
  // src/AHB.v(51)
  // src/AHB.v(51)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~(~D*B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1111010100110001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg6_b12|U_AHB/reg6_b10  (
    .a({\PWM5/FreCnt [12],open_n33372}),
    .b({\PWM5/FreCnt [15],open_n33373}),
    .c({\PWM5/FreCntr [12],pwm_state_read[5]}),
    .ce(\U_AHB/n14 ),
    .clk(clk100m),
    .d({\PWM5/FreCntr [15],\PWM5/n0_lutinv }),
    .mi({\U_AHB/h2h_hwdata [12],\U_AHB/h2h_hwdata [10]}),
    .f({_al_u1457_o,\PWM5/n24 }),
    .q({freq5[12],freq5[10]}));  // src/AHB.v(51)
  // src/AHB.v(51)
  // src/AHB.v(51)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(C*B*A*~(0@D))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(C*B*A*~(1@D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg6_b14|U_AHB/reg6_b17  (
    .a({_al_u1448_o,_al_u1449_o}),
    .b({_al_u1450_o,\PWM5/FreCnt [17]}),
    .c({_al_u1451_o,\PWM5/FreCnt [8]}),
    .ce(\U_AHB/n14 ),
    .clk(clk100m),
    .d({\PWM5/FreCnt [14],\PWM5/FreCntr [17]}),
    .e({\PWM5/FreCntr [14],\PWM5/FreCntr [8]}),
    .mi({\U_AHB/h2h_hwdata [14],\U_AHB/h2h_hwdata [17]}),
    .f({_al_u1452_o,_al_u1450_o}),
    .q({freq5[14],freq5[17]}));  // src/AHB.v(51)
  // src/AHB.v(51)
  // src/AHB.v(51)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(~(D*~B)*~(C*~A))"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(~(D*~B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b1000110010101111),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b1000110010101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg6_b15|U_AHB/reg6_b13  (
    .a({\PWM5/FreCnt [12],open_n33404}),
    .b({\PWM5/FreCnt [15],limit_r_pad[5]}),
    .c({\PWM5/FreCntr [12],limit_l_pad[5]}),
    .ce(\U_AHB/n14 ),
    .clk(clk100m),
    .d({\PWM5/FreCntr [15],\PWM5/n11 }),
    .mi({\U_AHB/h2h_hwdata [15],\U_AHB/h2h_hwdata [13]}),
    .f({_al_u1453_o,_al_u3023_o}),
    .q({freq5[15],freq5[13]}));  // src/AHB.v(51)
  // src/AHB.v(51)
  // src/AHB.v(51)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg6_b18|U_AHB/reg6_b21  (
    .a({\PWM5/FreCnt [16],_al_u924_o}),
    .b({\PWM5/FreCnt [17],\PWM5/FreCnt [2]}),
    .c({\PWM5/FreCnt [18],\PWM5/FreCnt [20]}),
    .ce(\U_AHB/n14 ),
    .clk(clk100m),
    .d({\PWM5/FreCnt [19],\PWM5/FreCnt [21]}),
    .e({open_n33423,\PWM5/FreCnt [22]}),
    .mi({\U_AHB/h2h_hwdata [18],\U_AHB/h2h_hwdata [21]}),
    .f({_al_u924_o,_al_u925_o}),
    .q({freq5[18],freq5[21]}));  // src/AHB.v(51)
  // src/AHB.v(51)
  // src/AHB.v(51)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(D@B)*~(C@A))"),
    //.LUT1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000010000100001),
    .INIT_LUT1(16'b1000010000100001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg6_b20|U_AHB/reg6_b22  (
    .a({\PWM5/FreCnt [20],\PWM5/FreCnt [22]}),
    .b({\PWM5/FreCnt [26],\PWM5/FreCnt [23]}),
    .c({\PWM5/FreCntr [20],\PWM5/FreCntr [22]}),
    .ce(\U_AHB/n14 ),
    .clk(clk100m),
    .d({\PWM5/FreCntr [26],\PWM5/FreCntr [23]}),
    .mi({\U_AHB/h2h_hwdata [20],\U_AHB/h2h_hwdata [22]}),
    .f({_al_u1451_o,_al_u1449_o}),
    .q({freq5[20],freq5[22]}));  // src/AHB.v(51)
  // src/AHB.v(51)
  // src/AHB.v(51)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg6_b23|U_AHB/reg6_b3  (
    .a({\PWM5/FreCnt [23],_al_u919_o}),
    .b({\PWM5/FreCnt [24],\PWM5/FreCnt [3]}),
    .c({\PWM5/FreCnt [25],\PWM5/FreCnt [4]}),
    .ce(\U_AHB/n14 ),
    .clk(clk100m),
    .d({\PWM5/FreCnt [26],\PWM5/FreCnt [5]}),
    .e({open_n33454,\PWM5/FreCnt [6]}),
    .mi({\U_AHB/h2h_hwdata [23],\U_AHB/h2h_hwdata [3]}),
    .f({_al_u919_o,_al_u920_o}),
    .q({freq5[23],freq5[3]}));  // src/AHB.v(51)
  // src/AHB.v(51)
  // src/AHB.v(51)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~D*~C*~B*A)"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(~D*~C*~B*A)"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b0000000000000010),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg6_b24|U_AHB/reg6_b7  (
    .a({\PWM5/FreCnt [0],_al_u920_o}),
    .b({\PWM5/FreCnt [24],\PWM5/FreCnt [7]}),
    .c({\PWM5/FreCntr [0],\PWM5/FreCnt [8]}),
    .ce(\U_AHB/n14 ),
    .clk(clk100m),
    .d({\PWM5/FreCntr [24],\PWM5/FreCnt [9]}),
    .mi({\U_AHB/h2h_hwdata [24],\U_AHB/h2h_hwdata [7]}),
    .f({_al_u1455_o,_al_u921_o}),
    .q({freq5[24],freq5[7]}));  // src/AHB.v(51)
  // src/AHB.v(51)
  // src/AHB.v(51)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(D@B)*~(C@A))"),
    //.LUTF1("(D*~(C@B))"),
    //.LUTG0("(~(D@B)*~(C@A))"),
    //.LUTG1("(D*~(C@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000010000100001),
    .INIT_LUTF1(16'b1100001100000000),
    .INIT_LUTG0(16'b1000010000100001),
    .INIT_LUTG1(16'b1100001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg6_b6|U_AHB/reg6_b4  (
    .a({open_n33489,\PWM5/FreCnt [16]}),
    .b({\PWM5/FreCnt [6],\PWM5/FreCnt [4]}),
    .c({\PWM5/FreCntr [6],\PWM5/FreCntr [16]}),
    .ce(\U_AHB/n14 ),
    .clk(clk100m),
    .d({_al_u1453_o,\PWM5/FreCntr [4]}),
    .mi({\U_AHB/h2h_hwdata [6],\U_AHB/h2h_hwdata [4]}),
    .f({_al_u1454_o,_al_u1447_o}),
    .q({freq5[6],freq5[4]}));  // src/AHB.v(51)
  // src/AHB.v(52)
  // src/AHB.v(52)
  EF2_PHY_MSLICE #(
    //.LUT0("(D*~C*~B*A)"),
    //.LUT1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000000000),
    .INIT_LUT1(16'b1000010000100001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg7_b10|U_AHB/reg7_b0  (
    .a({\PWM6/FreCnt [0],\U_AHB/h2h_hwrite }),
    .b({\PWM6/FreCnt [10],\U_AHB/h2h_haddr [13]}),
    .c({\PWM6/FreCntr [0],\U_AHB/h2h_haddr [14]}),
    .ce(\U_AHB/n16 ),
    .clk(clk100m),
    .d({\PWM6/FreCntr [10],\U_AHB/h2h_haddr [6]}),
    .mi({\U_AHB/h2h_hwdata [10],\U_AHB/h2h_hwdata [0]}),
    .f({_al_u1472_o,\U_AHB/n16 }),
    .q({freq6[10],freq6[0]}));  // src/AHB.v(52)
  // src/AHB.v(52)
  // src/AHB.v(52)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(~(D*~B)*~(~C*A))"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(~(D*~B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b1100010011110101),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b1100010011110101),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg7_b11|U_AHB/reg7_b12  (
    .a({\PWM6/FreCnt [10],open_n33522}),
    .b({\PWM6/FreCnt [19],limit_l_pad[6]}),
    .c({\PWM6/FreCntr [11],limit_r_pad[6]}),
    .ce(\U_AHB/n16 ),
    .clk(clk100m),
    .d({\PWM6/FreCntr [20],\PWM6/n11 }),
    .mi({\U_AHB/h2h_hwdata [11],\U_AHB/h2h_hwdata [12]}),
    .f({_al_u2231_o,_al_u3026_o}),
    .q({freq6[11],freq6[12]}));  // src/AHB.v(52)
  // src/AHB.v(52)
  // src/AHB.v(52)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(C*B*A*~(0@D))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(C*B*A*~(1@D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg7_b14|U_AHB/reg7_b18  (
    .a({_al_u1465_o,_al_u1464_o}),
    .b({_al_u1467_o,\PWM6/FreCnt [18]}),
    .c({_al_u1468_o,\PWM6/FreCnt [5]}),
    .ce(\U_AHB/n16 ),
    .clk(clk100m),
    .d({\PWM6/FreCnt [14],\PWM6/FreCntr [18]}),
    .e({\PWM6/FreCntr [14],\PWM6/FreCntr [5]}),
    .mi({\U_AHB/h2h_hwdata [14],\U_AHB/h2h_hwdata [18]}),
    .f({_al_u1469_o,_al_u1465_o}),
    .q({freq6[14],freq6[18]}));  // src/AHB.v(52)
  // src/AHB.v(52)
  // src/AHB.v(52)
  EF2_PHY_MSLICE #(
    //.LUT0("(~D*~C*~B*A)"),
    //.LUT1("(C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000010),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg7_b15|U_AHB/reg7_b9  (
    .a({open_n33557,_al_u1216_o}),
    .b({open_n33558,\PWMD/FreCnt [7]}),
    .c({\PWM6/FreCntr [16],\PWMD/FreCnt [8]}),
    .ce(\U_AHB/n16 ),
    .clk(clk100m),
    .d({\PWM6/FreCnt [15],\PWMD/FreCnt [9]}),
    .mi({\U_AHB/h2h_hwdata [15],\U_AHB/h2h_hwdata [9]}),
    .f({_al_u2250_o,_al_u1217_o}),
    .q({freq6[15],freq6[9]}));  // src/AHB.v(52)
  // src/AHB.v(52)
  // src/AHB.v(52)
  EF2_PHY_MSLICE #(
    //.LUT0("(~D*~C*~B*A)"),
    //.LUT1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000010),
    .INIT_LUT1(16'b1000010000100001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg7_b16|U_AHB/reg7_b7  (
    .a({\PWM6/FreCnt [16],_al_u957_o}),
    .b({\PWM6/FreCnt [4],\PWM6/FreCnt [7]}),
    .c({\PWM6/FreCntr [16],\PWM6/FreCnt [8]}),
    .ce(\U_AHB/n16 ),
    .clk(clk100m),
    .d({\PWM6/FreCntr [4],\PWM6/FreCnt [9]}),
    .mi({\U_AHB/h2h_hwdata [16],\U_AHB/h2h_hwdata [7]}),
    .f({_al_u1464_o,_al_u958_o}),
    .q({freq6[16],freq6[7]}));  // src/AHB.v(52)
  // src/AHB.v(52)
  // src/AHB.v(52)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg7_b17|U_AHB/reg7_b6  (
    .a({\PWM6/FreCnt [17],_al_u1474_o}),
    .b({\PWM6/FreCnt [9],\PWM6/FreCnt [6]}),
    .c({\PWM6/FreCntr [17],\PWM6/FreCnt [8]}),
    .ce(\U_AHB/n16 ),
    .clk(clk100m),
    .d({\PWM6/FreCntr [9],\PWM6/FreCntr [6]}),
    .e({open_n33587,\PWM6/FreCntr [8]}),
    .mi({\U_AHB/h2h_hwdata [17],\U_AHB/h2h_hwdata [6]}),
    .f({_al_u1474_o,_al_u1475_o}),
    .q({freq6[17],freq6[6]}));  // src/AHB.v(52)
  // src/AHB.v(52)
  // src/AHB.v(52)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg7_b19|U_AHB/reg7_b21  (
    .a({\PWM6/FreCnt [16],_al_u961_o}),
    .b({\PWM6/FreCnt [17],\PWM6/FreCnt [2]}),
    .c({\PWM6/FreCnt [18],\PWM6/FreCnt [20]}),
    .ce(\U_AHB/n16 ),
    .clk(clk100m),
    .d({\PWM6/FreCnt [19],\PWM6/FreCnt [21]}),
    .e({open_n33604,\PWM6/FreCnt [22]}),
    .mi({\U_AHB/h2h_hwdata [19],\U_AHB/h2h_hwdata [21]}),
    .f({_al_u961_o,_al_u962_o}),
    .q({freq6[19],freq6[21]}));  // src/AHB.v(52)
  // src/AHB.v(52)
  // src/AHB.v(52)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(D@B)*~(C@A))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(~(D@B)*~(C@A))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000010000100001),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000010000100001),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg7_b20|U_AHB/reg7_b22  (
    .a({\PWM6/FreCnt [20],\PWM6/FreCnt [22]}),
    .b({\PWM6/FreCnt [26],\PWM6/FreCnt [23]}),
    .c({\PWM6/FreCntr [20],\PWM6/FreCntr [22]}),
    .ce(\U_AHB/n16 ),
    .clk(clk100m),
    .d({\PWM6/FreCntr [26],\PWM6/FreCntr [23]}),
    .mi({\U_AHB/h2h_hwdata [20],\U_AHB/h2h_hwdata [22]}),
    .f({_al_u1468_o,_al_u1466_o}),
    .q({freq6[20],freq6[22]}));  // src/AHB.v(52)
  // src/AHB.v(52)
  // src/AHB.v(52)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg7_b23|U_AHB/reg7_b3  (
    .a({\PWM6/FreCnt [23],_al_u956_o}),
    .b({\PWM6/FreCnt [24],\PWM6/FreCnt [3]}),
    .c({\PWM6/FreCnt [25],\PWM6/FreCnt [4]}),
    .ce(\U_AHB/n16 ),
    .clk(clk100m),
    .d({\PWM6/FreCnt [26],\PWM6/FreCnt [5]}),
    .e({open_n33639,\PWM6/FreCnt [6]}),
    .mi({\U_AHB/h2h_hwdata [23],\U_AHB/h2h_hwdata [3]}),
    .f({_al_u956_o,_al_u957_o}),
    .q({freq6[23],freq6[3]}));  // src/AHB.v(52)
  // src/AHB.v(52)
  // src/AHB.v(52)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg7_b4|U_AHB/reg7_b13  (
    .a({\PWM6/FreCnt [0],_al_u959_o}),
    .b({\PWM6/FreCnt [1],\PWM6/FreCnt [12]}),
    .c({\PWM6/FreCnt [10],\PWM6/FreCnt [13]}),
    .ce(\U_AHB/n16 ),
    .clk(clk100m),
    .d({\PWM6/FreCnt [11],\PWM6/FreCnt [14]}),
    .e({open_n33656,\PWM6/FreCnt [15]}),
    .mi({\U_AHB/h2h_hwdata [4],\U_AHB/h2h_hwdata [13]}),
    .f({_al_u959_o,_al_u960_o}),
    .q({freq6[4],freq6[13]}));  // src/AHB.v(52)
  // src/AHB.v(52)
  // src/AHB.v(52)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(D@B)*~(C@A))"),
    //.LUT1("(C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000010000100001),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg7_b5|U_AHB/reg7_b25  (
    .a({open_n33673,\PWM6/FreCnt [11]}),
    .b({open_n33674,\PWM6/FreCnt [25]}),
    .c({\PWME/FreCntr [6],\PWM6/FreCntr [11]}),
    .ce(\U_AHB/n16 ),
    .clk(clk100m),
    .d({\PWME/FreCnt [5],\PWM6/FreCntr [25]}),
    .mi({\U_AHB/h2h_hwdata [5],\U_AHB/h2h_hwdata [25]}),
    .f({_al_u2875_o,_al_u1476_o}),
    .q({freq6[5],freq6[25]}));  // src/AHB.v(52)
  // src/AHB.v(53)
  // src/AHB.v(53)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(D*~C*~B*A)"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(D*~C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b0000001000000000),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b0000001000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg8_b0|U_AHB/reg8_b13  (
    .a({\U_AHB/h2h_hwrite ,_al_u1495_o}),
    .b({\U_AHB/h2h_haddr [13],\PWM7/FreCnt [13]}),
    .c({\U_AHB/h2h_haddr [14],\PWM7/FreCnt [19]}),
    .ce(\U_AHB/n18 ),
    .clk(clk100m),
    .d({\U_AHB/h2h_haddr [7],\PWM7/FreCntr [13]}),
    .e({open_n33689,\PWM7/FreCntr [19]}),
    .mi({\U_AHB/h2h_hwdata [0],\U_AHB/h2h_hwdata [13]}),
    .f({\U_AHB/n18 ,_al_u1496_o}),
    .q({freq7[0],freq7[13]}));  // src/AHB.v(53)
  // src/AHB.v(53)
  // src/AHB.v(53)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg8_b10|U_AHB/reg8_b14  (
    .a({\PWM7/FreCnt [10],_al_u1493_o}),
    .b({\PWM7/FreCnt [2],\PWM7/FreCnt [14]}),
    .c({\PWM7/FreCntr [10],\PWM7/FreCnt [20]}),
    .ce(\U_AHB/n18 ),
    .clk(clk100m),
    .d({\PWM7/FreCntr [2],\PWM7/FreCntr [14]}),
    .e({open_n33706,\PWM7/FreCntr [20]}),
    .mi({\U_AHB/h2h_hwdata [10],\U_AHB/h2h_hwdata [14]}),
    .f({_al_u1487_o,_al_u1494_o}),
    .q({freq7[10],freq7[14]}));  // src/AHB.v(53)
  // src/AHB.v(53)
  // src/AHB.v(53)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(~(D*~B)*~(C*~A))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(~(D*~B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b1000110010101111),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1000110010101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg8_b12|U_AHB/reg8_b11  (
    .a({\PWM7/FreCnt [12],open_n33723}),
    .b({\PWM7/FreCnt [15],open_n33724}),
    .c({\PWM7/FreCntr [12],pwm_state_read[7]}),
    .ce(\U_AHB/n18 ),
    .clk(clk100m),
    .d({\PWM7/FreCntr [15],\PWM7/n0_lutinv }),
    .mi(\U_AHB/h2h_hwdata [12:11]),
    .f({_al_u1486_o,\PWM7/n24 }),
    .q(freq7[12:11]));  // src/AHB.v(53)
  // src/AHB.v(53)
  // src/AHB.v(53)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(~(C*~B)*~(D*~A))"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(~(C*~B)*~(D*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b1000101011001111),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b1000101011001111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg8_b16|U_AHB/reg8_b15  (
    .a({\PWM7/FreCnt [1],open_n33743}),
    .b({\PWM7/FreCnt [15],limit_l_pad[7]}),
    .c({\PWM7/FreCntr [16],limit_r_pad[7]}),
    .ce(\U_AHB/n18 ),
    .clk(clk100m),
    .d({\PWM7/FreCntr [2],\PWM7/n11 }),
    .mi(\U_AHB/h2h_hwdata [16:15]),
    .f({_al_u2311_o,_al_u3029_o}),
    .q(freq7[16:15]));  // src/AHB.v(53)
  // src/AHB.v(53)
  // src/AHB.v(53)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*B*A*~(0@D))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(C*B*A*~(1@D))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg8_b18|U_AHB/reg8_b3  (
    .a({\PWM7/FreCnt [18],_al_u1481_o}),
    .b({\PWM7/FreCnt [5],_al_u1483_o}),
    .c({\PWM7/FreCntr [18],_al_u1484_o}),
    .ce(\U_AHB/n18 ),
    .clk(clk100m),
    .d({\PWM7/FreCntr [5],\PWM7/FreCnt [3]}),
    .e({open_n33762,\PWM7/FreCntr [3]}),
    .mi({\U_AHB/h2h_hwdata [18],\U_AHB/h2h_hwdata [3]}),
    .f({_al_u1484_o,_al_u1485_o}),
    .q({freq7[18],freq7[3]}));  // src/AHB.v(53)
  // src/AHB.v(53)
  // src/AHB.v(53)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg8_b19|U_AHB/reg8_b20  (
    .a({\PWM7/FreCnt [16],_al_u998_o}),
    .b({\PWM7/FreCnt [17],\PWM7/FreCnt [2]}),
    .c({\PWM7/FreCnt [18],\PWM7/FreCnt [20]}),
    .ce(\U_AHB/n18 ),
    .clk(clk100m),
    .d({\PWM7/FreCnt [19],\PWM7/FreCnt [21]}),
    .e({open_n33779,\PWM7/FreCnt [22]}),
    .mi({\U_AHB/h2h_hwdata [19],\U_AHB/h2h_hwdata [20]}),
    .f({_al_u998_o,_al_u999_o}),
    .q({freq7[19],freq7[20]}));  // src/AHB.v(53)
  // src/AHB.v(53)
  // src/AHB.v(53)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*B*A*~(0@D))"),
    //.LUTF1("(~(~D*B)*~(~C*A))"),
    //.LUTG0("(C*B*A*~(1@D))"),
    //.LUTG1("(~(~D*B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b1111010100110001),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b1111010100110001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg8_b1|U_AHB/reg8_b6  (
    .a({\PWM7/FreCnt [1],_al_u1488_o}),
    .b({\PWM7/FreCnt [15],_al_u1490_o}),
    .c({\PWM7/FreCntr [1],_al_u1491_o}),
    .ce(\U_AHB/n18 ),
    .clk(clk100m),
    .d({\PWM7/FreCntr [15],\PWM7/FreCnt [0]}),
    .e({open_n33796,\PWM7/FreCntr [0]}),
    .mi({\U_AHB/h2h_hwdata [1],\U_AHB/h2h_hwdata [6]}),
    .f({_al_u1491_o,_al_u1492_o}),
    .q({freq7[1],freq7[6]}));  // src/AHB.v(53)
  // src/AHB.v(53)
  // src/AHB.v(53)
  EF2_PHY_MSLICE #(
    //.LUT0("(~D*~C*~B*A)"),
    //.LUT1("(B*A*~(D@C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000010),
    .INIT_LUT1(16'b1000000000001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg8_b21|U_AHB/reg8_b9  (
    .a({_al_u1486_o,_al_u1105_o}),
    .b({_al_u1487_o,\PWMA/FreCnt [7]}),
    .c({\PWM7/FreCnt [21],\PWMA/FreCnt [8]}),
    .ce(\U_AHB/n18 ),
    .clk(clk100m),
    .d({\PWM7/FreCntr [21],\PWMA/FreCnt [9]}),
    .mi({\U_AHB/h2h_hwdata [21],\U_AHB/h2h_hwdata [9]}),
    .f({_al_u1488_o,_al_u1106_o}),
    .q({freq7[21],freq7[9]}));  // src/AHB.v(53)
  // src/AHB.v(53)
  // src/AHB.v(53)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg8_b22|U_AHB/reg8_b17  (
    .a({\PWM7/FreCnt [22],_al_u1480_o}),
    .b({\PWM7/FreCnt [23],\PWM7/FreCnt [17]}),
    .c({\PWM7/FreCntr [22],\PWM7/FreCnt [8]}),
    .ce(\U_AHB/n18 ),
    .clk(clk100m),
    .d({\PWM7/FreCntr [23],\PWM7/FreCntr [17]}),
    .e({open_n33827,\PWM7/FreCntr [8]}),
    .mi({\U_AHB/h2h_hwdata [22],\U_AHB/h2h_hwdata [17]}),
    .f({_al_u1480_o,_al_u1481_o}),
    .q({freq7[22],freq7[17]}));  // src/AHB.v(53)
  // src/AHB.v(53)
  // src/AHB.v(53)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg8_b23|U_AHB/reg8_b4  (
    .a({\PWM7/FreCnt [23],_al_u993_o}),
    .b({\PWM7/FreCnt [24],\PWM7/FreCnt [3]}),
    .c({\PWM7/FreCnt [25],\PWM7/FreCnt [4]}),
    .ce(\U_AHB/n18 ),
    .clk(clk100m),
    .d({\PWM7/FreCnt [26],\PWM7/FreCnt [5]}),
    .e({open_n33844,\PWM7/FreCnt [6]}),
    .mi({\U_AHB/h2h_hwdata [23],\U_AHB/h2h_hwdata [4]}),
    .f({_al_u993_o,_al_u994_o}),
    .q({freq7[23],freq7[4]}));  // src/AHB.v(53)
  // src/AHB.v(53)
  // src/AHB.v(53)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~D*~C*~B*A)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(~D*~C*~B*A)"),
    //.LUTG1("(C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000000000000010),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg8_b25|U_AHB/reg8_b7  (
    .a({open_n33861,_al_u994_o}),
    .b({open_n33862,\PWM7/FreCnt [7]}),
    .c({\PWM7/FreCntr [1],\PWM7/FreCnt [8]}),
    .ce(\U_AHB/n18 ),
    .clk(clk100m),
    .d({\PWM7/FreCnt [1],\PWM7/FreCnt [9]}),
    .mi({\U_AHB/h2h_hwdata [25],\U_AHB/h2h_hwdata [7]}),
    .f({_al_u1489_o,_al_u995_o}),
    .q({freq7[25],freq7[7]}));  // src/AHB.v(53)
  // src/AHB.v(53)
  // src/AHB.v(53)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg8_b26|U_AHB/reg8_b5  (
    .a({\PWM7/FreCnt [0],_al_u996_o}),
    .b({\PWM7/FreCnt [1],\PWM7/FreCnt [12]}),
    .c({\PWM7/FreCnt [10],\PWM7/FreCnt [13]}),
    .ce(\U_AHB/n18 ),
    .clk(clk100m),
    .d({\PWM7/FreCnt [11],\PWM7/FreCnt [14]}),
    .e({open_n33881,\PWM7/FreCnt [15]}),
    .mi({\U_AHB/h2h_hwdata [26],\U_AHB/h2h_hwdata [5]}),
    .f({_al_u996_o,_al_u997_o}),
    .q({freq7[26],freq7[5]}));  // src/AHB.v(53)
  // src/AHB.v(54)
  // src/AHB.v(54)
  EF2_PHY_MSLICE #(
    //.LUT0("(D*~C*~B*A)"),
    //.LUT1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000001000000000),
    .INIT_LUT1(16'b1000010000100001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg9_b10|U_AHB/reg9_b0  (
    .a({\PWM8/FreCnt [10],\U_AHB/h2h_hwrite }),
    .b({\PWM8/FreCnt [2],\U_AHB/h2h_haddr [13]}),
    .c({\PWM8/FreCntr [10],\U_AHB/h2h_haddr [14]}),
    .ce(\U_AHB/n20 ),
    .clk(clk100m),
    .d({\PWM8/FreCntr [2],\U_AHB/h2h_haddr [8]}),
    .mi({\U_AHB/h2h_hwdata [10],\U_AHB/h2h_hwdata [0]}),
    .f({_al_u1505_o,\U_AHB/n20 }),
    .q({freq8[10],freq8[0]}));  // src/AHB.v(54)
  // src/AHB.v(54)
  // src/AHB.v(54)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    //.LUT1("(~(D*~B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000000000000),
    .INIT_LUT1(16'b1000110010101111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg9_b15|U_AHB/reg9_b14  (
    .a({\PWM8/FreCnt [12],open_n33912}),
    .b({\PWM8/FreCnt [15],limit_l_pad[8]}),
    .c({\PWM8/FreCntr [12],limit_r_pad[8]}),
    .ce(\U_AHB/n20 ),
    .clk(clk100m),
    .d({\PWM8/FreCntr [15],\PWM8/n11 }),
    .mi(\U_AHB/h2h_hwdata [15:14]),
    .f({_al_u1504_o,_al_u3032_o}),
    .q(freq8[15:14]));  // src/AHB.v(54)
  // src/AHB.v(54)
  // src/AHB.v(54)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg9_b16|U_AHB/reg9_b13  (
    .a({\PWM8/FreCnt [16],_al_u1513_o}),
    .b({\PWM8/FreCnt [26],\PWM8/FreCnt [13]}),
    .c({\PWM8/FreCntr [16],\PWM8/FreCnt [19]}),
    .ce(\U_AHB/n20 ),
    .clk(clk100m),
    .d({\PWM8/FreCntr [26],\PWM8/FreCntr [13]}),
    .e({open_n33927,\PWM8/FreCntr [19]}),
    .mi({\U_AHB/h2h_hwdata [16],\U_AHB/h2h_hwdata [13]}),
    .f({_al_u1513_o,_al_u1514_o}),
    .q({freq8[16],freq8[13]}));  // src/AHB.v(54)
  // src/AHB.v(54)
  // src/AHB.v(54)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg9_b17|U_AHB/reg9_b20  (
    .a({\PWM8/FreCnt [16],_al_u1035_o}),
    .b({\PWM8/FreCnt [17],\PWM8/FreCnt [2]}),
    .c({\PWM8/FreCnt [18],\PWM8/FreCnt [20]}),
    .ce(\U_AHB/n20 ),
    .clk(clk100m),
    .d({\PWM8/FreCnt [19],\PWM8/FreCnt [21]}),
    .e({open_n33944,\PWM8/FreCnt [22]}),
    .mi({\U_AHB/h2h_hwdata [17],\U_AHB/h2h_hwdata [20]}),
    .f({_al_u1035_o,_al_u1036_o}),
    .q({freq8[17],freq8[20]}));  // src/AHB.v(54)
  // src/AHB.v(54)
  // src/AHB.v(54)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(~0*C)*~(D*~B))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(A*~(~1*C)*~(D*~B))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000001010),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000100010101010),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg9_b18|U_AHB/reg9_b11  (
    .a({\PWM8/FreCnt [18],_al_u2393_o}),
    .b({\PWM8/FreCnt [5],\PWM8/FreCnt [10]}),
    .c({\PWM8/FreCntr [18],\PWM8/FreCnt [17]}),
    .ce(\U_AHB/n20 ),
    .clk(clk100m),
    .d({\PWM8/FreCntr [5],\PWM8/FreCntr [11]}),
    .e({open_n33961,\PWM8/FreCntr [18]}),
    .mi({\U_AHB/h2h_hwdata [18],\U_AHB/h2h_hwdata [11]}),
    .f({_al_u1502_o,_al_u2394_o}),
    .q({freq8[18],freq8[11]}));  // src/AHB.v(54)
  // src/AHB.v(54)
  // src/AHB.v(54)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*B*A*~(0@D))"),
    //.LUTF1("(~(~D*B)*~(~C*A))"),
    //.LUTG0("(C*B*A*~(1@D))"),
    //.LUTG1("(~(~D*B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b1111010100110001),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b1111010100110001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg9_b1|U_AHB/reg9_b5  (
    .a({\PWM8/FreCnt [1],_al_u1506_o}),
    .b({\PWM8/FreCnt [15],_al_u1508_o}),
    .c({\PWM8/FreCntr [1],_al_u1509_o}),
    .ce(\U_AHB/n20 ),
    .clk(clk100m),
    .d({\PWM8/FreCntr [15],\PWM8/FreCnt [0]}),
    .e({open_n33978,\PWM8/FreCntr [0]}),
    .mi({\U_AHB/h2h_hwdata [1],\U_AHB/h2h_hwdata [5]}),
    .f({_al_u1509_o,_al_u1510_o}),
    .q({freq8[1],freq8[5]}));  // src/AHB.v(54)
  // src/AHB.v(54)
  // src/AHB.v(54)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(D@B)*~(C@A))"),
    //.LUT1("(~(~D*B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000010000100001),
    .INIT_LUT1(16'b1010111100100011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg9_b21|U_AHB/reg9_b22  (
    .a({\PWM8/FreCnt [21],\PWM8/FreCnt [22]}),
    .b({\PWM8/FreCnt [7],\PWM8/FreCnt [23]}),
    .c({\PWM8/FreCntr [22],\PWM8/FreCntr [22]}),
    .ce(\U_AHB/n20 ),
    .clk(clk100m),
    .d({\PWM8/FreCntr [8],\PWM8/FreCntr [23]}),
    .mi({\U_AHB/h2h_hwdata [21],\U_AHB/h2h_hwdata [22]}),
    .f({_al_u2403_o,_al_u1498_o}),
    .q({freq8[21],freq8[22]}));  // src/AHB.v(54)
  // src/AHB.v(54)
  // src/AHB.v(54)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg9_b23|U_AHB/reg9_b3  (
    .a({\PWM8/FreCnt [23],_al_u1030_o}),
    .b({\PWM8/FreCnt [24],\PWM8/FreCnt [3]}),
    .c({\PWM8/FreCnt [25],\PWM8/FreCnt [4]}),
    .ce(\U_AHB/n20 ),
    .clk(clk100m),
    .d({\PWM8/FreCnt [26],\PWM8/FreCnt [5]}),
    .e({open_n34009,\PWM8/FreCnt [6]}),
    .mi({\U_AHB/h2h_hwdata [23],\U_AHB/h2h_hwdata [3]}),
    .f({_al_u1030_o,_al_u1031_o}),
    .q({freq8[23],freq8[3]}));  // src/AHB.v(54)
  // src/AHB.v(54)
  // src/AHB.v(54)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~A*~(0@C)*~(~D*B))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(~A*~(1@C)*~(~D*B))"),
    //.LUTG1("(C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010100000001),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0101000000010000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg9_b24|U_AHB/reg9_b12  (
    .a({open_n34026,_al_u1507_o}),
    .b({open_n34027,\PWM8/FreCnt [12]}),
    .c({\PWM8/FreCntr [1],\PWM8/FreCnt [24]}),
    .ce(\U_AHB/n20 ),
    .clk(clk100m),
    .d({\PWM8/FreCnt [1],\PWM8/FreCntr [12]}),
    .e({open_n34028,\PWM8/FreCntr [24]}),
    .mi({\U_AHB/h2h_hwdata [24],\U_AHB/h2h_hwdata [12]}),
    .f({_al_u1507_o,_al_u1508_o}),
    .q({freq8[24],freq8[12]}));  // src/AHB.v(54)
  // src/AHB.v(54)
  // src/AHB.v(54)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~D*~C*~B*A)"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(~D*~C*~B*A)"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b0000000000000010),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg9_b25|U_AHB/reg9_b7  (
    .a({\PWM8/FreCnt [11],_al_u1031_o}),
    .b({\PWM8/FreCnt [25],\PWM8/FreCnt [7]}),
    .c({\PWM8/FreCntr [11],\PWM8/FreCnt [8]}),
    .ce(\U_AHB/n20 ),
    .clk(clk100m),
    .d({\PWM8/FreCntr [25],\PWM8/FreCnt [9]}),
    .mi({\U_AHB/h2h_hwdata [25],\U_AHB/h2h_hwdata [7]}),
    .f({_al_u1511_o,_al_u1032_o}),
    .q({freq8[25],freq8[7]}));  // src/AHB.v(54)
  // src/AHB.v(54)
  // src/AHB.v(54)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \U_AHB/reg9_b26|U_AHB/reg9_b4  (
    .a({\PWM8/FreCnt [0],_al_u1033_o}),
    .b({\PWM8/FreCnt [1],\PWM8/FreCnt [12]}),
    .c({\PWM8/FreCnt [10],\PWM8/FreCnt [13]}),
    .ce(\U_AHB/n20 ),
    .clk(clk100m),
    .d({\PWM8/FreCnt [11],\PWM8/FreCnt [14]}),
    .e({open_n34063,\PWM8/FreCnt [15]}),
    .mi({\U_AHB/h2h_hwdata [26],\U_AHB/h2h_hwdata [4]}),
    .f({_al_u1033_o,_al_u1034_o}),
    .q({freq8[26],freq8[4]}));  // src/AHB.v(54)
  EF2_PHY_PLL #(
    .CLKC0_CPHASE(4),
    .CLKC0_DIV(5),
    .CLKC0_DIV2_ENABLE("DISABLE"),
    .CLKC0_DUTY(0.500000),
    .CLKC0_DUTY50("ENABLE"),
    .CLKC0_DUTY_INT(3),
    .CLKC0_ENABLE("ENABLE"),
    .CLKC0_FPHASE(0),
    .CLKC1_CPHASE(9),
    .CLKC1_DIV(10),
    .CLKC1_DIV2_ENABLE("DISABLE"),
    .CLKC1_DUTY(0.500000),
    .CLKC1_DUTY50("ENABLE"),
    .CLKC1_DUTY_INT(5),
    .CLKC1_ENABLE("ENABLE"),
    .CLKC1_FPHASE(0),
    .CLKC2_CPHASE(39),
    .CLKC2_DIV(40),
    .CLKC2_DIV2_ENABLE("DISABLE"),
    .CLKC2_ENABLE("ENABLE"),
    .CLKC2_FPHASE(0),
    .CLKC3_CPHASE(124),
    .CLKC3_DIV(125),
    .CLKC3_DIV2_ENABLE("DISABLE"),
    .CLKC3_ENABLE("ENABLE"),
    .CLKC3_FPHASE(0),
    .CLKC4_CPHASE(1),
    .CLKC4_DIV(1),
    .CLKC4_DIV2_ENABLE("DISABLE"),
    .CLKC4_ENABLE("DISABLE"),
    .CLKC4_FPHASE(0),
    .CLKC5_CPHASE(1),
    .CLKC5_DIV(1),
    .CLKC5_DIV2_ENABLE("DISABLE"),
    .CLKC5_ENABLE("DISABLE"),
    .CLKC6_CPHASE(1),
    .CLKC6_DIV(1),
    .CLKC6_DIV2_ENABLE("DISABLE"),
    .CLKC6_ENABLE("DISABLE"),
    .DERIVE_PLL_CLOCKS("DISABLE"),
    .DPHASE_SOURCE("DISABLE"),
    .DYNCFG("DISABLE"),
    .FBCLK_DIV(40),
    .FEEDBK_MODE("NOCOMP"),
    .FEEDBK_PATH("VCO_PHASE_0"),
    .FIN("25.000"),
    .FREQ_LOCK_ACCURACY(2),
    .FREQ_OFFSET("0.000000"),
    .FREQ_OFFSET_INT("0"),
    .GEN_BASIC_CLOCK("DISABLE"),
    .GMC_GAIN(6),
    .GMC_TEST(14),
    .HIGH_SPEED_EN("ENABLE"),
    .ICP_CURRENT(3),
    .IF_ESCLKSTSW("DISABLE"),
    .INTFB_WAKE("DISABLE"),
    .INTPI(3),
    .KVCO(6),
    .LPF_CAPACITOR(3),
    .LPF_RESISTOR(2),
    .NORESET("DISABLE"),
    .ODIV_MUXC0("DIV"),
    .ODIV_MUXC1("DIV"),
    .ODIV_MUXC2("DIV"),
    .ODIV_MUXC3("DIV"),
    .ODIV_MUXC4("DIV"),
    .OFFSET_MODE("EXT"),
    .PLLC2RST_ENA("DISABLE"),
    .PLLC34RST_ENA("DISABLE"),
    .PLLMRST_ENA("DISABLE"),
    .PLLRST_ENA("ENABLE"),
    .PLL_LOCK_MODE(0),
    .PREDIV_MUXC0("VCO"),
    .PREDIV_MUXC1("VCO"),
    .PREDIV_MUXC2("VCO"),
    .PREDIV_MUXC3("VCO"),
    .PREDIV_MUXC4("VCO"),
    .PREDIV_MUXC5("VCO"),
    .PREDIV_MUXC6("VCO"),
    .PU_INTP("DISABLE"),
    .REFCLK_DIV(1),
    .REFCLK_SEL("INTERNAL"),
    .SSC_AMP("0.000000"),
    .SSC_ENABLE("DISABLE"),
    .SSC_FREQ_DIV(0),
    .SSC_MODE("Down"),
    .SSC_RNGE(0),
    .STDBY_ENABLE("DISABLE"),
    .STDBY_VCO_ENA("DISABLE"),
    .SYNC_ENABLE("DISABLE"),
    .VCO_NORESET("DISABLE"))
    \U_PLL/pll_inst  (
    .daddr(6'b000000),
    .dclk(1'b0),
    .dcs(1'b0),
    .di(8'b00000000),
    .dsm_refclk(1'b0),
    .dsm_rst(1'b0),
    .dwe(1'b0),
    .fbclk(1'b0),
    .frac_offset_valid(1'b0),
    .psclk(1'b0),
    .psclksel(3'b000),
    .psdown(1'b0),
    .psstep(1'b0),
    .refclk(clkin_pad),
    .reset(1'b0),
    .ssc_en(1'b0),
    .stdby(1'b0),
    .clkc({open_n34080,open_n34081,open_n34082,open_n34083,clk25m,clk100m_keep,open_n34084}),
    .extlock(rstn));  // al_ip/PLL.v(92)
  EF2_PHY_PAD #(
    //.LOCATION("P70"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u100 (
    .ipad(limit_r[5]),
    .di(limit_r_pad[5]));  // CPLD_SOC_AHB_TOP.v(6)
  EF2_PHY_PAD #(
    //.LOCATION("P59"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u101 (
    .ipad(limit_r[4]),
    .di(limit_r_pad[4]));  // CPLD_SOC_AHB_TOP.v(6)
  EF2_PHY_PAD #(
    //.LOCATION("P57"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u102 (
    .ipad(limit_r[3]),
    .di(limit_r_pad[3]));  // CPLD_SOC_AHB_TOP.v(6)
  EF2_PHY_PAD #(
    //.LOCATION("P55"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u103 (
    .ipad(limit_r[2]),
    .di(limit_r_pad[2]));  // CPLD_SOC_AHB_TOP.v(6)
  EF2_PHY_PAD #(
    //.LOCATION("P49"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u104 (
    .ipad(limit_r[1]),
    .di(limit_r_pad[1]));  // CPLD_SOC_AHB_TOP.v(6)
  EF2_PHY_PAD #(
    //.LOCATION("P40"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u105 (
    .ipad(limit_r[0]),
    .di(limit_r_pad[0]));  // CPLD_SOC_AHB_TOP.v(6)
  EF2_PHY_PAD #(
    //.LOCATION("P111"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u106 (
    .do({open_n34233,open_n34234,open_n34235,pwm_pad[15]}),
    .opad(pwm[15]));  // CPLD_SOC_AHB_TOP.v(7)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~D*~C*~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1067|PWM9/reg0_b23  (
    .a({\PWM9/FreCnt [23],open_n34255}),
    .b({\PWM9/FreCnt [24],\PWM9/n12 [23]}),
    .c({\PWM9/FreCnt [25],freq9[23]}),
    .clk(clk100m),
    .d({\PWM9/FreCnt [26],\PWM9/n0_lutinv }),
    .sr(\PWM9/n11 ),
    .f({_al_u1067_o,open_n34269}),
    .q({open_n34273,\PWM9/FreCnt [23]}));  // src/OnePWM.v(37)
  // src/AHB.v(54)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~D*~C*~B*A)"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(~D*~C*~B*A)"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b0000000000000010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1068|U_AHB/reg9_b9  (
    .a({_al_u1067_o,_al_u1068_o}),
    .b({\PWM9/FreCnt [3],\PWM9/FreCnt [7]}),
    .c({\PWM9/FreCnt [4],\PWM9/FreCnt [8]}),
    .ce(\U_AHB/n20 ),
    .clk(clk100m),
    .d({\PWM9/FreCnt [5],\PWM9/FreCnt [9]}),
    .e({\PWM9/FreCnt [6],open_n34274}),
    .mi({open_n34276,\U_AHB/h2h_hwdata [9]}),
    .f({_al_u1068_o,_al_u1069_o}),
    .q({open_n34292,freq8[9]}));  // src/AHB.v(54)
  EF2_PHY_PAD #(
    //.LOCATION("P112"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u107 (
    .do({open_n34294,open_n34295,open_n34296,pwm_pad[14]}),
    .opad(pwm[14]));  // CPLD_SOC_AHB_TOP.v(7)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1070|PWM9/reg0_b1  (
    .a({\PWM9/FreCnt [0],open_n34316}),
    .b({\PWM9/FreCnt [1],\PWM9/n12 [1]}),
    .c({\PWM9/FreCnt [10],freq9[1]}),
    .clk(clk100m),
    .d({\PWM9/FreCnt [11],\PWM9/n0_lutinv }),
    .sr(\PWM9/n11 ),
    .f({_al_u1070_o,open_n34334}),
    .q({open_n34338,\PWM9/FreCnt [1]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1071|PWM9/reg0_b15  (
    .a({_al_u1070_o,open_n34339}),
    .b({\PWM9/FreCnt [12],\PWM9/n12 [15]}),
    .c({\PWM9/FreCnt [13],freq9[15]}),
    .clk(clk100m),
    .d({\PWM9/FreCnt [14],\PWM9/n0_lutinv }),
    .e({\PWM9/FreCnt [15],open_n34341}),
    .sr(\PWM9/n11 ),
    .f({_al_u1071_o,open_n34356}),
    .q({open_n34360,\PWM9/FreCnt [15]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1072|PWM9/reg0_b19  (
    .a({\PWM9/FreCnt [16],open_n34361}),
    .b({\PWM9/FreCnt [17],\PWM9/n12 [19]}),
    .c({\PWM9/FreCnt [18],freq9[19]}),
    .clk(clk100m),
    .d({\PWM9/FreCnt [19],\PWM9/n0_lutinv }),
    .sr(\PWM9/n11 ),
    .f({_al_u1072_o,open_n34379}),
    .q({open_n34383,\PWM9/FreCnt [19]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1073|PWM9/reg0_b21  (
    .a({_al_u1072_o,open_n34384}),
    .b({\PWM9/FreCnt [2],\PWM9/n12 [21]}),
    .c({\PWM9/FreCnt [20],freq9[21]}),
    .clk(clk100m),
    .d({\PWM9/FreCnt [21],\PWM9/n0_lutinv }),
    .e({\PWM9/FreCnt [22],open_n34386}),
    .sr(\PWM9/n11 ),
    .f({_al_u1073_o,open_n34401}),
    .q({open_n34405,\PWM9/FreCnt [21]}));  // src/OnePWM.v(37)
  EF2_PHY_PAD #(
    //.LOCATION("P115"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u108 (
    .do({open_n34407,open_n34408,open_n34409,pwm_pad[13]}),
    .opad(pwm[13]));  // CPLD_SOC_AHB_TOP.v(7)
  EF2_PHY_PAD #(
    //.LOCATION("P117"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u109 (
    .do({open_n34430,open_n34431,open_n34432,pwm_pad[12]}),
    .opad(pwm[12]));  // CPLD_SOC_AHB_TOP.v(7)
  EF2_PHY_PAD #(
    //.LOCATION("P52"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u110 (
    .do({open_n34453,open_n34454,open_n34455,pwm_pad[11]}),
    .opad(pwm[11]));  // CPLD_SOC_AHB_TOP.v(7)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~D*~C*~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1104|PWMA/reg0_b23  (
    .a({\PWMA/FreCnt [23],open_n34475}),
    .b({\PWMA/FreCnt [24],\PWMA/n12 [23]}),
    .c({\PWMA/FreCnt [25],freqA[23]}),
    .clk(clk100m),
    .d({\PWMA/FreCnt [26],\PWMA/n0_lutinv }),
    .sr(\PWMA/n11 ),
    .f({_al_u1104_o,open_n34489}),
    .q({open_n34493,\PWMA/FreCnt [23]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*B*A*~(0@D))"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(C*B*A*~(1@D))"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1105|PWMA/reg1_b4  (
    .a({_al_u1104_o,_al_u1534_o}),
    .b({\PWMA/FreCnt [3],_al_u1536_o}),
    .c({\PWMA/FreCnt [4],_al_u1537_o}),
    .ce(\PWMA/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d(\PWMA/FreCnt [5:4]),
    .e({\PWMA/FreCnt [6],\PWMA/FreCntr [4]}),
    .mi({open_n34495,freqA[4]}),
    .f({_al_u1105_o,_al_u1538_o}),
    .q({open_n34511,\PWMA/FreCntr [4]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*B*A*~(0@D))"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(C*B*A*~(1@D))"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1107|PWMA/reg1_b2  (
    .a({\PWMA/FreCnt [0],_al_u2557_o}),
    .b({\PWMA/FreCnt [1],_al_u2559_o}),
    .c({\PWMA/FreCnt [10],_al_u2560_o}),
    .ce(\PWMA/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMA/FreCnt [11],\PWMA/FreCnt [1]}),
    .e({open_n34512,\PWMA/FreCntr [2]}),
    .mi({open_n34514,freqA[2]}),
    .f({_al_u1107_o,_al_u2561_o}),
    .q({open_n34530,\PWMA/FreCntr [2]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1108|PWMA/reg0_b12  (
    .a({_al_u1107_o,open_n34531}),
    .b({\PWMA/FreCnt [12],\PWMA/n12 [12]}),
    .c({\PWMA/FreCnt [13],freqA[12]}),
    .clk(clk100m),
    .d({\PWMA/FreCnt [14],\PWMA/n0_lutinv }),
    .e({\PWMA/FreCnt [15],open_n34533}),
    .sr(\PWMA/n11 ),
    .f({_al_u1108_o,open_n34548}),
    .q({open_n34552,\PWMA/FreCnt [12]}));  // src/OnePWM.v(37)
  // src/AHB.v(54)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1109|U_AHB/reg9_b8  (
    .a({\PWMA/FreCnt [16],_al_u1533_o}),
    .b({\PWMA/FreCnt [17],\PWMA/FreCnt [17]}),
    .c({\PWMA/FreCnt [18],\PWMA/FreCnt [8]}),
    .ce(\U_AHB/n20 ),
    .clk(clk100m),
    .d({\PWMA/FreCnt [19],\PWMA/FreCntr [17]}),
    .e({open_n34553,\PWMA/FreCntr [8]}),
    .mi({open_n34555,\U_AHB/h2h_hwdata [8]}),
    .f({_al_u1109_o,_al_u1534_o}),
    .q({open_n34571,freq8[8]}));  // src/AHB.v(54)
  EF2_PHY_PAD #(
    //.LOCATION("P47"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u111 (
    .do({open_n34573,open_n34574,open_n34575,pwm_pad[10]}),
    .opad(pwm[10]));  // CPLD_SOC_AHB_TOP.v(7)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1110|PWMA/reg1_b23  (
    .a({_al_u1109_o,open_n34595}),
    .b({\PWMA/FreCnt [2],_al_u1108_o}),
    .c({\PWMA/FreCnt [20],_al_u1110_o}),
    .ce(\PWMA/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMA/FreCnt [21],_al_u1106_o}),
    .e({\PWMA/FreCnt [22],open_n34596}),
    .mi({open_n34598,freqA[23]}),
    .f({_al_u1110_o,\PWMA/n0_lutinv }),
    .q({open_n34614,\PWMA/FreCntr [23]}));  // src/OnePWM.v(37)
  EF2_PHY_PAD #(
    //.LOCATION("P44"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u112 (
    .do({open_n34616,open_n34617,open_n34618,pwm_pad[9]}),
    .opad(pwm[9]));  // CPLD_SOC_AHB_TOP.v(7)
  EF2_PHY_SPAD #(
    //.LOCATION("P107"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("16"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u113 (
    .do({open_n34640,pwm_pad[8]}),
    .ts(1'b1),
    .opad(pwm[8]));  // CPLD_SOC_AHB_TOP.v(7)
  EF2_PHY_PAD #(
    //.LOCATION("P113"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u114 (
    .do({open_n34648,open_n34649,open_n34650,pwm_pad[7]}),
    .opad(pwm[7]));  // CPLD_SOC_AHB_TOP.v(7)
  // src/AHB.v(57)
  EF2_PHY_LSLICE #(
    //.LUTF0("(D*~(C@B))"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(D*~(C@B))"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100001100000000),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b1100001100000000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1144|U_AHB/reg12_b6  (
    .a({\PWMB/FreCnt [0],open_n34670}),
    .b({\PWMB/FreCnt [1],\PWMB/FreCnt [6]}),
    .c({\PWMB/FreCnt [10],\PWMB/FreCntr [6]}),
    .ce(\U_AHB/n26 ),
    .clk(clk100m),
    .d({\PWMB/FreCnt [11],_al_u1557_o}),
    .mi({open_n34674,\U_AHB/h2h_hwdata [6]}),
    .f({_al_u1144_o,_al_u1558_o}),
    .q({open_n34690,freqB[6]}));  // src/AHB.v(57)
  // src/OnePWM.v(15)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u1145|PWMB/stopreq_reg  (
    .a({_al_u1144_o,open_n34691}),
    .b({\PWMB/FreCnt [12],open_n34692}),
    .c({\PWMB/FreCnt [13],\PWMB/stopreq }),
    .clk(clk100m),
    .d({\PWMB/FreCnt [14],\PWMB/n0_lutinv }),
    .e({\PWMB/FreCnt [15],open_n34694}),
    .sr(pwm_start_stop[11]),
    .f({_al_u1145_o,open_n34709}),
    .q({open_n34713,\PWMB/stopreq_keep }));  // src/OnePWM.v(15)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~D*~C*~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1146|PWMB/reg0_b19  (
    .a({\PWMB/FreCnt [16],open_n34714}),
    .b({\PWMB/FreCnt [17],\PWMB/n12 [19]}),
    .c({\PWMB/FreCnt [18],freqB[19]}),
    .clk(clk100m),
    .d({\PWMB/FreCnt [19],\PWMB/n0_lutinv }),
    .sr(\PWMB/n11 ),
    .f({_al_u1146_o,open_n34728}),
    .q({open_n34732,\PWMB/FreCnt [19]}));  // src/OnePWM.v(37)
  EF2_PHY_PAD #(
    //.LOCATION("P121"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u115 (
    .do({open_n34734,open_n34735,open_n34736,pwm_pad[6]}),
    .opad(pwm[6]));  // CPLD_SOC_AHB_TOP.v(7)
  EF2_PHY_SPAD #(
    //.LOCATION("P25"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("16"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u116 (
    .do({open_n34758,pwm_pad[5]}),
    .ts(1'b1),
    .opad(pwm[5]));  // CPLD_SOC_AHB_TOP.v(7)
  EF2_PHY_PAD #(
    //.LOCATION("P125"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u117 (
    .do({open_n34766,open_n34767,open_n34768,pwm_pad[4]}),
    .opad(pwm[4]));  // CPLD_SOC_AHB_TOP.v(7)
  EF2_PHY_PAD #(
    //.LOCATION("P126"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u118 (
    .do({open_n34789,open_n34790,open_n34791,pwm_pad[3]}),
    .opad(pwm[3]));  // CPLD_SOC_AHB_TOP.v(7)
  // src/AHB.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(~C*D)"),
    //.LUT1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000111100000000),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1181|U_AHB/reg13_b25  (
    .a({\PWMC/FreCnt [0],open_n34811}),
    .b({\PWMC/FreCnt [1],open_n34812}),
    .c({\PWMC/FreCnt [10],\PWMC/FreCntr [26]}),
    .ce(\U_AHB/n28 ),
    .clk(clk100m),
    .d({\PWMC/FreCnt [11],\PWMC/FreCnt [25]}),
    .mi({open_n34823,\U_AHB/h2h_hwdata [25]}),
    .f({_al_u1181_o,_al_u2716_o}),
    .q({open_n34828,freqC[25]}));  // src/AHB.v(58)
  // src/AHB.v(58)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*B*A*~(0@D))"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(C*B*A*~(1@D))"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1182|U_AHB/reg13_b14  (
    .a({_al_u1181_o,_al_u1569_o}),
    .b({\PWMC/FreCnt [12],_al_u1571_o}),
    .c({\PWMC/FreCnt [13],_al_u1572_o}),
    .ce(\U_AHB/n28 ),
    .clk(clk100m),
    .d({\PWMC/FreCnt [14],\PWMC/FreCnt [14]}),
    .e({\PWMC/FreCnt [15],\PWMC/FreCntr [14]}),
    .mi({open_n34830,\U_AHB/h2h_hwdata [14]}),
    .f({_al_u1182_o,_al_u1573_o}),
    .q({open_n34846,freqC[14]}));  // src/AHB.v(58)
  EF2_PHY_PAD #(
    //.LOCATION("P127"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u119 (
    .do({open_n34848,open_n34849,open_n34850,pwm_pad[2]}),
    .opad(pwm[2]));  // CPLD_SOC_AHB_TOP.v(7)
  EF2_PHY_PAD #(
    //.LOCATION("P128"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u120 (
    .do({open_n34871,open_n34872,open_n34873,pwm_pad[1]}),
    .opad(pwm[1]));  // CPLD_SOC_AHB_TOP.v(7)
  EF2_PHY_PAD #(
    //.LOCATION("P141"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u121 (
    .do({open_n34894,open_n34895,open_n34896,pwm_pad[0]}),
    .opad(pwm[0]));  // CPLD_SOC_AHB_TOP.v(7)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1215|PWMD/reg0_b23  (
    .a({\PWMD/FreCnt [23],open_n34916}),
    .b({\PWMD/FreCnt [24],\PWMD/n12 [23]}),
    .c({\PWMD/FreCnt [25],freqD[23]}),
    .clk(clk100m),
    .d({\PWMD/FreCnt [26],\PWMD/n0_lutinv }),
    .sr(\PWMD/n11 ),
    .f({_al_u1215_o,open_n34934}),
    .q({open_n34938,\PWMD/FreCnt [23]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1216|PWMD/reg0_b6  (
    .a({_al_u1215_o,open_n34939}),
    .b({\PWMD/FreCnt [3],\PWMD/n12 [6]}),
    .c({\PWMD/FreCnt [4],freqD[6]}),
    .clk(clk100m),
    .d({\PWMD/FreCnt [5],\PWMD/n0_lutinv }),
    .e({\PWMD/FreCnt [6],open_n34941}),
    .sr(\PWMD/n11 ),
    .f({_al_u1216_o,open_n34956}),
    .q({open_n34960,\PWMD/FreCnt [6]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1218|PWMD/reg0_b1  (
    .a({\PWMD/FreCnt [0],open_n34961}),
    .b({\PWMD/FreCnt [1],\PWMD/n12 [1]}),
    .c({\PWMD/FreCnt [10],freqD[1]}),
    .clk(clk100m),
    .d({\PWMD/FreCnt [11],\PWMD/n0_lutinv }),
    .sr(\PWMD/n11 ),
    .f({_al_u1218_o,open_n34979}),
    .q({open_n34983,\PWMD/FreCnt [1]}));  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(~0*~D*~C*~B*A)"),
    //.LUT1("(~1*~D*~C*~B*A)"),
    .INIT_LUT0(16'b0000000000000010),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1219 (
    .a({_al_u1218_o,_al_u1218_o}),
    .b({\PWMD/FreCnt [12],\PWMD/FreCnt [12]}),
    .c({\PWMD/FreCnt [13],\PWMD/FreCnt [13]}),
    .d({\PWMD/FreCnt [14],\PWMD/FreCnt [14]}),
    .mi({open_n34996,\PWMD/FreCnt [15]}),
    .fx({open_n35001,_al_u1219_o}));
  EF2_PHY_PAD #(
    //.LOCATION("P38"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u122 (
    .ipad(rst_n),
    .di(rst_n_pad));  // CPLD_SOC_AHB_TOP.v(4)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1220|PWMD/reg0_b19  (
    .a({\PWMD/FreCnt [16],open_n35027}),
    .b({\PWMD/FreCnt [17],\PWMD/n12 [19]}),
    .c({\PWMD/FreCnt [18],freqD[19]}),
    .clk(clk100m),
    .d({\PWMD/FreCnt [19],\PWMD/n0_lutinv }),
    .sr(\PWMD/n11 ),
    .f({_al_u1220_o,open_n35045}),
    .q({open_n35049,\PWMD/FreCnt [19]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(D@B)*~(C@A))"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(~(D@B)*~(C@A))"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000010000100001),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b1000010000100001),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1221|PWMD/reg1_b23  (
    .a({_al_u1220_o,\PWMD/FreCnt [22]}),
    .b({\PWMD/FreCnt [2],\PWMD/FreCnt [23]}),
    .c({\PWMD/FreCnt [20],\PWMD/FreCntr [22]}),
    .ce(\PWMD/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMD/FreCnt [21],\PWMD/FreCntr [23]}),
    .e({\PWMD/FreCnt [22],open_n35050}),
    .mi({open_n35052,freqD[23]}),
    .f({_al_u1221_o,_al_u1587_o}),
    .q({open_n35068,\PWMD/FreCntr [23]}));  // src/OnePWM.v(37)
  // src/AHB.v(54)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(D@B)*~(C@A))"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(~(D@B)*~(C@A))"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000010000100001),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b1000010000100001),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1253|U_AHB/reg9_b6  (
    .a({_al_u1252_o,\PWME/FreCnt [6]}),
    .b({\PWME/FreCnt [3],\PWME/FreCnt [7]}),
    .c({\PWME/FreCnt [4],\PWME/FreCntr [6]}),
    .ce(\U_AHB/n20 ),
    .clk(clk100m),
    .d({\PWME/FreCnt [5],\PWME/FreCntr [7]}),
    .e({\PWME/FreCnt [6],open_n35069}),
    .mi({open_n35071,\U_AHB/h2h_hwdata [6]}),
    .f({_al_u1253_o,_al_u1604_o}),
    .q({open_n35087,freq8[6]}));  // src/AHB.v(54)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1255|PWME/reg0_b1  (
    .a({\PWME/FreCnt [0],open_n35088}),
    .b({\PWME/FreCnt [1],\PWME/n12 [1]}),
    .c({\PWME/FreCnt [10],freqE[1]}),
    .clk(clk100m),
    .d({\PWME/FreCnt [11],\PWME/n0_lutinv }),
    .sr(\PWME/n11 ),
    .f({_al_u1255_o,open_n35106}),
    .q({open_n35110,\PWME/FreCnt [1]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1256|PWME/reg0_b15  (
    .a({_al_u1255_o,open_n35111}),
    .b({\PWME/FreCnt [12],\PWME/n12 [15]}),
    .c({\PWME/FreCnt [13],freqE[15]}),
    .clk(clk100m),
    .d({\PWME/FreCnt [14],\PWME/n0_lutinv }),
    .e({\PWME/FreCnt [15],open_n35113}),
    .sr(\PWME/n11 ),
    .f({_al_u1256_o,open_n35128}),
    .q({open_n35132,\PWME/FreCnt [15]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~D*~C*~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1257|PWME/reg0_b19  (
    .a({\PWME/FreCnt [16],open_n35133}),
    .b({\PWME/FreCnt [17],\PWME/n12 [19]}),
    .c({\PWME/FreCnt [18],freqE[19]}),
    .clk(clk100m),
    .d({\PWME/FreCnt [19],\PWME/n0_lutinv }),
    .sr(\PWME/n11 ),
    .f({_al_u1257_o,open_n35147}),
    .q({open_n35151,\PWME/FreCnt [19]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1258|PWME/reg0_b21  (
    .a({_al_u1257_o,open_n35152}),
    .b({\PWME/FreCnt [2],\PWME/n12 [21]}),
    .c({\PWME/FreCnt [20],freqE[21]}),
    .clk(clk100m),
    .d({\PWME/FreCnt [21],\PWME/n0_lutinv }),
    .e({\PWME/FreCnt [22],open_n35154}),
    .sr(\PWME/n11 ),
    .f({_al_u1258_o,open_n35169}),
    .q({open_n35173,\PWME/FreCnt [21]}));  // src/OnePWM.v(37)
  // src/AHB.v(62)
  EF2_PHY_MSLICE #(
    //.LUT0("(~D*~C*~B*~A)"),
    //.LUT1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000001),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1292|U_AHB/reg16_b24  (
    .a({\PWMF/FreCnt [0],pnumcntB[18]}),
    .b({\PWMF/FreCnt [1],pnumcntB[19]}),
    .c({\PWMF/FreCnt [10],pnumcntB[1]}),
    .ce(\U_AHB/n34 ),
    .clk(clk100m),
    .d({\PWMF/FreCnt [11],pnumcntB[20]}),
    .mi({open_n35184,\U_AHB/h2h_hwdata [24]}),
    .f({_al_u1292_o,_al_u2579_o}),
    .q({open_n35189,freqF[24]}));  // src/AHB.v(62)
  // src/OnePWM.v(15)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u1293|PWMF/stopreq_reg  (
    .a({_al_u1292_o,open_n35190}),
    .b({\PWMF/FreCnt [12],open_n35191}),
    .c({\PWMF/FreCnt [13],\PWMF/stopreq }),
    .clk(clk100m),
    .d({\PWMF/FreCnt [14],\PWMF/n0_lutinv }),
    .e({\PWMF/FreCnt [15],open_n35193}),
    .sr(pwm_start_stop[15]),
    .f({_al_u1293_o,open_n35208}),
    .q({open_n35212,\PWMF/stopreq_keep }));  // src/OnePWM.v(15)
  // src/AHB.v(62)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1294|U_AHB/reg16_b21  (
    .a({\PWMF/FreCnt [16],_al_u1294_o}),
    .b({\PWMF/FreCnt [17],\PWMF/FreCnt [2]}),
    .c({\PWMF/FreCnt [18],\PWMF/FreCnt [20]}),
    .ce(\U_AHB/n34 ),
    .clk(clk100m),
    .d({\PWMF/FreCnt [19],\PWMF/FreCnt [21]}),
    .e({open_n35213,\PWMF/FreCnt [22]}),
    .mi({open_n35215,\U_AHB/h2h_hwdata [21]}),
    .f({_al_u1294_o,_al_u1295_o}),
    .q({open_n35231,freqF[21]}));  // src/AHB.v(62)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1369|PWM0/reg0_b1  (
    .b({open_n35234,\PWM0/n12 [1]}),
    .c({\PWM0/FreCntr [1],freq0[1]}),
    .clk(clk100m),
    .d({\PWM0/FreCnt [1],\PWM0/n0_lutinv }),
    .sr(\PWM0/n11 ),
    .f({_al_u1369_o,open_n35252}),
    .q({open_n35256,\PWM0/FreCnt [1]}));  // src/OnePWM.v(37)
  // src/AHB.v(46)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~A*~(0@C)*~(~D*B))"),
    //.LUTF1("(C*B*A*~(0@D))"),
    //.LUTG0("(~A*~(1@C)*~(~D*B))"),
    //.LUTG1("(C*B*A*~(1@D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010100000001),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b0101000000010000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1372|U_AHB/reg1_b12  (
    .a({_al_u1368_o,_al_u1369_o}),
    .b({_al_u1370_o,\PWM0/FreCnt [12]}),
    .c({_al_u1371_o,\PWM0/FreCnt [24]}),
    .ce(\U_AHB/n2 ),
    .clk(clk100m),
    .d({\PWM0/FreCnt [0],\PWM0/FreCntr [12]}),
    .e({\PWM0/FreCntr [0],\PWM0/FreCntr [24]}),
    .mi({open_n35258,\U_AHB/h2h_hwdata [12]}),
    .f({_al_u1372_o,_al_u1370_o}),
    .q({open_n35274,freq0[12]}));  // src/AHB.v(46)
  // src/AHB.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~D*B)*~(~C*A))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(~(~D*B)*~(~C*A))"),
    //.LUTG1("(C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111010100110001),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b1111010100110001),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1404|U_AHB/reg3_b1  (
    .a({open_n35275,\PWM2/FreCnt [1]}),
    .b({open_n35276,\PWM2/FreCnt [15]}),
    .c({\PWM2/FreCntr [1],\PWM2/FreCntr [1]}),
    .ce(\U_AHB/n8 ),
    .clk(clk100m),
    .d({\PWM2/FreCnt [1],\PWM2/FreCntr [15]}),
    .mi({open_n35280,\U_AHB/h2h_hwdata [1]}),
    .f({_al_u1404_o,_al_u1406_o}),
    .q({open_n35296,freq2[1]}));  // src/AHB.v(48)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*B*A*~(0@D))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*B*A*~(1@D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1407|PWM2/reg1_b0  (
    .a({_al_u1403_o,open_n35297}),
    .b({_al_u1405_o,open_n35298}),
    .c({_al_u1406_o,\PWM2/n11 }),
    .ce(\PWM2/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM2/FreCnt [0],\PWM2/n0_lutinv }),
    .e({\PWM2/FreCntr [0],open_n35299}),
    .mi({open_n35301,freq2[0]}),
    .f({_al_u1407_o,\PWM2/mux3_b0_sel_is_3_o }),
    .q({open_n35317,\PWM2/FreCntr [0]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(45)
  EF2_PHY_LSLICE #(
    //.LUTF0("~(~C*~D)"),
    //.LUTF1("(0*D*C*B*A)"),
    //.LUTG0("~(~C*~D)"),
    //.LUTG1("(1*D*C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111111111110000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1111111111110000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1478|PWM6/pwm_reg  (
    .a({_al_u1469_o,open_n35318}),
    .b({_al_u1471_o,open_n35319}),
    .c({_al_u1473_o,pwm_pad[6]}),
    .clk(clk100m),
    .d({_al_u1475_o,\PWM6/n18_lutinv }),
    .e({_al_u1477_o,open_n35321}),
    .sr(\PWM6/u14_sel_is_1_o ),
    .f({\PWM6/n18_lutinv ,open_n35336}),
    .q({open_n35340,\PWM6/pwm_keep }));  // src/OnePWM.v(45)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~(D@B)*~(C@A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1000010000100001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1516|PWM9/reg0_b3  (
    .a({\PWM9/FreCnt [16],open_n35341}),
    .b({\PWM9/FreCnt [3],\PWM9/n12 [3]}),
    .c({\PWM9/FreCntr [16],freq9[3]}),
    .clk(clk100m),
    .d({\PWM9/FreCntr [3],\PWM9/n0_lutinv }),
    .sr(\PWM9/n11 ),
    .f({_al_u1516_o,open_n35355}),
    .q({open_n35359,\PWM9/FreCnt [3]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(A*~(0@C)*~(D@B))"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(A*~(1@C)*~(D@B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b0000100000000010),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1000000000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1517|PWM9/reg0_b5  (
    .a({_al_u1516_o,open_n35360}),
    .b({\PWM9/FreCnt [18],\PWM9/n12 [5]}),
    .c({\PWM9/FreCnt [5],freq9[5]}),
    .clk(clk100m),
    .d({\PWM9/FreCntr [18],\PWM9/n0_lutinv }),
    .e({\PWM9/FreCntr [5],open_n35362}),
    .sr(\PWM9/n11 ),
    .f({_al_u1517_o,open_n35377}),
    .q({open_n35381,\PWM9/FreCnt [5]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~A*~(0*~C)*~(D@B))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(~A*~(1*~C)*~(D@B))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0100010000010001),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b0100000000010000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1518|PWM9/reg1_b23  (
    .a({\PWM9/FreCnt [22],_al_u2484_o}),
    .b(\PWM9/FreCnt [23:22]),
    .c({\PWM9/FreCntr [22],\PWM9/FreCnt [3]}),
    .ce(\PWM9/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM9/FreCntr [23],\PWM9/FreCntr [23]}),
    .e({open_n35382,\PWM9/FreCntr [4]}),
    .mi({open_n35384,freq9[23]}),
    .f({_al_u1518_o,_al_u2485_o}),
    .q({open_n35400,\PWM9/FreCntr [23]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(D*~(C@B))"),
    //.LUTF1("(A*~(0@C)*~(D@B))"),
    //.LUTG0("(D*~(C@B))"),
    //.LUTG1("(A*~(1@C)*~(D@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100001100000000),
    .INIT_LUTF1(16'b0000100000000010),
    .INIT_LUTG0(16'b1100001100000000),
    .INIT_LUTG1(16'b1000000000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1519|PWM9/reg1_b3  (
    .a({_al_u1518_o,open_n35401}),
    .b({\PWM9/FreCnt [17],\PWM9/FreCnt [2]}),
    .c({\PWM9/FreCnt [8],\PWM9/FreCntr [3]}),
    .ce(\PWM9/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM9/FreCntr [17],_al_u2491_o}),
    .e({\PWM9/FreCntr [8],open_n35402}),
    .mi({open_n35404,freq9[3]}),
    .f({_al_u1519_o,_al_u2492_o}),
    .q({open_n35420,\PWM9/FreCntr [3]}));  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(C*B*A*~(0@D))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(C*B*A*~(1@D))"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1521|_al_u1586  (
    .a({_al_u1517_o,_al_u1585_o}),
    .b({_al_u1519_o,\PWMD/FreCnt [18]}),
    .c({_al_u1520_o,\PWMD/FreCnt [5]}),
    .d({\PWM9/FreCnt [14],\PWMD/FreCntr [18]}),
    .e({\PWM9/FreCntr [14],\PWMD/FreCntr [5]}),
    .f({_al_u1521_o,_al_u1586_o}));
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~(D*~B)*~(C*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1000110010101111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1522|PWM9/reg0_b12  (
    .a({\PWM9/FreCnt [12],open_n35443}),
    .b({\PWM9/FreCnt [15],\PWM9/n12 [12]}),
    .c({\PWM9/FreCntr [12],freq9[12]}),
    .clk(clk100m),
    .d({\PWM9/FreCntr [15],\PWM9/n0_lutinv }),
    .sr(\PWM9/n11 ),
    .f({_al_u1522_o,open_n35457}),
    .q({open_n35461,\PWM9/FreCnt [12]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(D*~(C@B))"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(D*~(C@B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1100001100000000),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1100001100000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1523|PWM9/reg0_b6  (
    .b({\PWM9/FreCnt [6],\PWM9/n12 [6]}),
    .c({\PWM9/FreCntr [6],freq9[6]}),
    .clk(clk100m),
    .d({_al_u1522_o,\PWM9/n0_lutinv }),
    .sr(\PWM9/n11 ),
    .f({_al_u1523_o,open_n35481}),
    .q({open_n35485,\PWM9/FreCnt [6]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1000010000100001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1524|PWM9/reg1_b0  (
    .a({\PWM9/FreCnt [0],open_n35486}),
    .b({\PWM9/FreCnt [24],open_n35487}),
    .c({\PWM9/FreCntr [0],\PWM9/n11 }),
    .ce(\PWM9/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM9/FreCntr [24],\PWM9/n0_lutinv }),
    .mi({open_n35498,freq9[0]}),
    .f({_al_u1524_o,\PWM9/mux3_b0_sel_is_3_o }),
    .q({open_n35503,\PWM9/FreCntr [0]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(A*~(0@C)*~(D@B))"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(A*~(1@C)*~(D@B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b0000100000000010),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1000000000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1525|PWM9/reg0_b13  (
    .a({_al_u1524_o,open_n35504}),
    .b({\PWM9/FreCnt [13],\PWM9/n12 [13]}),
    .c({\PWM9/FreCnt [19],freq9[13]}),
    .clk(clk100m),
    .d({\PWM9/FreCntr [13],\PWM9/n0_lutinv }),
    .e({\PWM9/FreCntr [19],open_n35506}),
    .sr(\PWM9/n11 ),
    .f({_al_u1525_o,open_n35521}),
    .q({open_n35525,\PWM9/FreCnt [13]}));  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*B*A*~(0@D))"),
    //.LUT1("(C*B*A*~(1@D))"),
    .INIT_LUT0(16'b0000000010000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1527 (
    .a({_al_u1523_o,_al_u1523_o}),
    .b({_al_u1525_o,_al_u1525_o}),
    .c({_al_u1526_o,_al_u1526_o}),
    .d({\PWM9/FreCnt [21],\PWM9/FreCnt [21]}),
    .mi({open_n35538,\PWM9/FreCntr [21]}),
    .fx({open_n35543,_al_u1527_o}));
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(A*~(0@C)*~(D@B))"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(A*~(1@C)*~(D@B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b0000100000000010),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1000000000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1529|PWM9/reg0_b4  (
    .a({_al_u1528_o,open_n35546}),
    .b({\PWM9/FreCnt [11],\PWM9/n12 [4]}),
    .c({\PWM9/FreCnt [4],freq9[4]}),
    .clk(clk100m),
    .d({\PWM9/FreCntr [11],\PWM9/n0_lutinv }),
    .e({\PWM9/FreCntr [4],open_n35548}),
    .sr(\PWM9/n11 ),
    .f({_al_u1529_o,open_n35563}),
    .q({open_n35567,\PWM9/FreCnt [4]}));  // src/OnePWM.v(37)
  // src/AHB.v(55)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(C*B)*~(D*A))"),
    //.LUT1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0001010100111111),
    .INIT_LUT1(16'b1000010000100001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1530|U_AHB/reg10_b25  (
    .a({\PWM9/FreCnt [2],\U_AHB/n113_lutinv }),
    .b({\PWM9/FreCnt [25],\U_AHB/n111 }),
    .c({\PWM9/FreCntr [2],pnumcntA[18]}),
    .ce(\U_AHB/n22 ),
    .clk(clk100m),
    .d({\PWM9/FreCntr [25],\U_AHB/h2h_hrdata [18]}),
    .mi({open_n35578,\U_AHB/h2h_hwdata [25]}),
    .f({_al_u1530_o,_al_u3242_o}),
    .q({open_n35583,freq9[25]}));  // src/AHB.v(55)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(A*~(0@C)*~(D@B))"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(A*~(1@C)*~(D@B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b0000100000000010),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1000000000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1531|PWM9/reg0_b2  (
    .a({_al_u1530_o,open_n35584}),
    .b({\PWM9/FreCnt [1],\PWM9/n12 [2]}),
    .c({\PWM9/FreCnt [10],freq9[2]}),
    .clk(clk100m),
    .d({\PWM9/FreCntr [1],\PWM9/n0_lutinv }),
    .e({\PWM9/FreCntr [10],open_n35586}),
    .sr(\PWM9/n11 ),
    .f({_al_u1531_o,open_n35601}),
    .q({open_n35605,\PWM9/FreCnt [2]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~(D*~B)*~(C*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1000110010101111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1539|PWMA/reg0_b15  (
    .a({\PWMA/FreCnt [12],open_n35606}),
    .b({\PWMA/FreCnt [15],\PWMA/n12 [15]}),
    .c({\PWMA/FreCntr [12],freqA[15]}),
    .clk(clk100m),
    .d({\PWMA/FreCntr [15],\PWMA/n0_lutinv }),
    .sr(\PWMA/n11 ),
    .f({_al_u1539_o,open_n35620}),
    .q({open_n35624,\PWMA/FreCnt [15]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(~0*C)*~(D@B))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(A*~(~1*C)*~(D@B))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000100000100010),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1540|PWMA/reg1_b3  (
    .a({\PWMA/FreCnt [10],_al_u2556_o}),
    .b(\PWMA/FreCnt [3:2]),
    .c({\PWMA/FreCntr [10],\PWMA/FreCnt [8]}),
    .ce(\PWMA/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMA/FreCntr [3],\PWMA/FreCntr [3]}),
    .e({open_n35625,\PWMA/FreCntr [9]}),
    .mi({open_n35627,freqA[3]}),
    .f({_al_u1540_o,_al_u2557_o}),
    .q({open_n35643,\PWMA/FreCntr [3]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(D*~(C@B))"),
    //.LUT1("(B*A*~(D@C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100001100000000),
    .INIT_LUT1(16'b1000000000001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1541|PWMA/reg1_b21  (
    .a({_al_u1539_o,open_n35644}),
    .b({_al_u1540_o,\PWMA/FreCnt [20]}),
    .c({\PWMA/FreCnt [21],\PWMA/FreCntr [21]}),
    .ce(\PWMA/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMA/FreCntr [21],_al_u2569_o}),
    .mi({open_n35655,freqA[21]}),
    .f({_al_u1541_o,_al_u2570_o}),
    .q({open_n35660,\PWMA/FreCntr [21]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1542|PWMA/reg0_b1  (
    .b({open_n35663,\PWMA/n12 [1]}),
    .c({\PWMA/FreCntr [1],freqA[1]}),
    .clk(clk100m),
    .d({\PWMA/FreCnt [1],\PWMA/n0_lutinv }),
    .sr(\PWMA/n11 ),
    .f({_al_u1542_o,open_n35681}),
    .q({open_n35685,\PWMA/FreCnt [1]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(15)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(~A*~(0@C)*~(~D*B))"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(~A*~(1@C)*~(~D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000010100000001),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0101000000010000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u1543|PWM7/stopreq_reg  (
    .a({_al_u1542_o,open_n35686}),
    .b({\PWMA/FreCnt [12],open_n35687}),
    .c({\PWMA/FreCnt [24],\PWM7/stopreq }),
    .clk(clk100m),
    .d({\PWMA/FreCntr [12],\PWM7/n0_lutinv }),
    .e({\PWMA/FreCntr [24],open_n35689}),
    .sr(pwm_start_stop[7]),
    .f({_al_u1543_o,open_n35704}),
    .q({open_n35708,\PWM7/stopreq_keep }));  // src/OnePWM.v(15)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~(~D*B)*~(~C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111010100110001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1544|PWMA/reg0_b2  (
    .a({\PWMA/FreCnt [1],open_n35709}),
    .b({\PWMA/FreCnt [15],\PWMA/n12 [2]}),
    .c({\PWMA/FreCntr [1],freqA[2]}),
    .clk(clk100m),
    .d({\PWMA/FreCntr [15],\PWMA/n0_lutinv }),
    .sr(\PWMA/n11 ),
    .f({_al_u1544_o,open_n35723}),
    .q({open_n35727,\PWMA/FreCnt [2]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*B*A*~(0@D))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*B*A*~(1@D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1545|PWMA/reg1_b0  (
    .a({_al_u1541_o,open_n35728}),
    .b({_al_u1543_o,open_n35729}),
    .c({_al_u1544_o,\PWMA/n11 }),
    .ce(\PWMA/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMA/FreCnt [0],\PWMA/n0_lutinv }),
    .e({\PWMA/FreCntr [0],open_n35730}),
    .mi({open_n35732,freqA[0]}),
    .f({_al_u1545_o,\PWMA/mux3_b0_sel_is_3_o }),
    .q({open_n35748,\PWMA/FreCntr [0]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~A*~(~0*C)*~(D@B))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(~A*~(~1*C)*~(D@B))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010000000001),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b0100010000010001),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1546|PWMA/reg1_b25  (
    .a({\PWMA/FreCnt [14],_al_u2558_o}),
    .b(\PWMA/FreCnt [25:24]),
    .c({\PWMA/FreCntr [14],\PWMA/FreCnt [3]}),
    .ce(\PWMA/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMA/FreCntr [25],\PWMA/FreCntr [25]}),
    .e({open_n35749,\PWMA/FreCntr [4]}),
    .mi({open_n35751,freqA[25]}),
    .f({_al_u1546_o,_al_u2559_o}),
    .q({open_n35767,\PWMA/FreCntr [25]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*B*A*~(0@D))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(C*B*A*~(1@D))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1548|PWMA/reg1_b17  (
    .a({\PWMA/FreCnt [13],_al_u2564_o}),
    .b({\PWMA/FreCnt [16],_al_u2566_o}),
    .c({\PWMA/FreCntr [13],_al_u2567_o}),
    .ce(\PWMA/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMA/FreCntr [16],\PWMA/FreCnt [16]}),
    .e({open_n35768,\PWMA/FreCntr [17]}),
    .mi({open_n35770,freqA[17]}),
    .f({_al_u1548_o,_al_u2568_o}),
    .q({open_n35786,\PWMA/FreCntr [17]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(A*~(0@C)*~(D@B))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(A*~(1@C)*~(D@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b0000100000000010),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000000000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1549|PWMA/reg1_b19  (
    .a({_al_u1548_o,_al_u2571_o}),
    .b(\PWMA/FreCnt [19:18]),
    .c({\PWMA/FreCnt [2],\PWMA/FreCnt [22]}),
    .ce(\PWMA/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMA/FreCntr [19],\PWMA/FreCntr [19]}),
    .e({\PWMA/FreCntr [2],\PWMA/FreCntr [23]}),
    .mi({open_n35788,freqA[19]}),
    .f({_al_u1549_o,_al_u2572_o}),
    .q({open_n35804,\PWMA/FreCntr [19]}));  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*B*A*~(0@D))"),
    //.LUT1("(C*B*A*~(1@D))"),
    .INIT_LUT0(16'b0000000010000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1556 (
    .a({_al_u1552_o,_al_u1552_o}),
    .b({_al_u1554_o,_al_u1554_o}),
    .c({_al_u1555_o,_al_u1555_o}),
    .d({\PWMB/FreCnt [14],\PWMB/FreCnt [14]}),
    .mi({open_n35817,\PWMB/FreCntr [14]}),
    .fx({open_n35822,_al_u1556_o}));
  // src/AHB.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*A*~(D@C))"),
    //.LUTF1("(~(D*~B)*~(C*~A))"),
    //.LUTG0("(B*A*~(D@C))"),
    //.LUTG1("(~(D*~B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000000000001000),
    .INIT_LUTF1(16'b1000110010101111),
    .INIT_LUTG0(16'b1000000000001000),
    .INIT_LUTG1(16'b1000110010101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1557|U_AHB/reg3_b21  (
    .a({\PWMB/FreCnt [12],_al_u1401_o}),
    .b({\PWMB/FreCnt [15],_al_u1402_o}),
    .c({\PWMB/FreCntr [12],\PWM2/FreCnt [21]}),
    .ce(\U_AHB/n8 ),
    .clk(clk100m),
    .d({\PWMB/FreCntr [15],\PWM2/FreCntr [21]}),
    .mi({open_n35828,\U_AHB/h2h_hwdata [21]}),
    .f({_al_u1557_o,_al_u1403_o}),
    .q({open_n35844,freq2[21]}));  // src/AHB.v(48)
  // src/AHB.v(57)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(D@B)*~(C@A))"),
    //.LUTF1("(A*~(0@C)*~(D@B))"),
    //.LUTG0("(~(D@B)*~(C@A))"),
    //.LUTG1("(A*~(1@C)*~(D@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000010000100001),
    .INIT_LUTF1(16'b0000100000000010),
    .INIT_LUTG0(16'b1000010000100001),
    .INIT_LUTG1(16'b1000000000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1566|U_AHB/reg12_b25  (
    .a({_al_u1565_o,\PWMB/FreCnt [2]}),
    .b({\PWMB/FreCnt [1],\PWMB/FreCnt [25]}),
    .c({\PWMB/FreCnt [10],\PWMB/FreCntr [2]}),
    .ce(\U_AHB/n26 ),
    .clk(clk100m),
    .d({\PWMB/FreCntr [1],\PWMB/FreCntr [25]}),
    .e({\PWMB/FreCntr [10],open_n35845}),
    .mi({open_n35847,\U_AHB/h2h_hwdata [25]}),
    .f({_al_u1566_o,_al_u1565_o}),
    .q({open_n35863,freqB[25]}));  // src/AHB.v(57)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1589|PWMD/reg0_b26  (
    .a({\PWMD/FreCnt [20],open_n35864}),
    .b({\PWMD/FreCnt [26],\PWMD/n12 [26]}),
    .c({\PWMD/FreCntr [20],freqD[26]}),
    .clk(clk100m),
    .d({\PWMD/FreCntr [26],\PWMD/n0_lutinv }),
    .sr(\PWMD/n11 ),
    .f({_al_u1589_o,open_n35882}),
    .q({open_n35886,\PWMD/FreCnt [26]}));  // src/OnePWM.v(37)
  // src/AHB.v(52)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(C*B*A*~(0@D))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(C*B*A*~(1@D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1590|U_AHB/reg7_b8  (
    .a({_al_u1586_o,_al_u1587_o}),
    .b({_al_u1588_o,\PWMD/FreCnt [17]}),
    .c({_al_u1589_o,\PWMD/FreCnt [8]}),
    .ce(\U_AHB/n16 ),
    .clk(clk100m),
    .d({\PWMD/FreCnt [14],\PWMD/FreCntr [17]}),
    .e({\PWMD/FreCntr [14],\PWMD/FreCntr [8]}),
    .mi({open_n35888,\U_AHB/h2h_hwdata [8]}),
    .f({_al_u1590_o,_al_u1588_o}),
    .q({open_n35904,freq6[8]}));  // src/AHB.v(52)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~(D*~B)*~(C*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1000110010101111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1591|PWMD/reg0_b15  (
    .a({\PWMD/FreCnt [12],open_n35905}),
    .b({\PWMD/FreCnt [15],\PWMD/n12 [15]}),
    .c({\PWMD/FreCntr [12],freqD[15]}),
    .clk(clk100m),
    .d({\PWMD/FreCntr [15],\PWMD/n0_lutinv }),
    .sr(\PWMD/n11 ),
    .f({_al_u1591_o,open_n35919}),
    .q({open_n35923,\PWMD/FreCnt [15]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*D)"),
    //.LUT1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000000000000),
    .INIT_LUT1(16'b1000010000100001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1593|PWMD/reg1_b0  (
    .a({\PWMD/FreCnt [0],open_n35924}),
    .b({\PWMD/FreCnt [24],open_n35925}),
    .c({\PWMD/FreCntr [0],\PWMD/n11 }),
    .ce(\PWMD/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMD/FreCntr [24],\PWMD/n0_lutinv }),
    .mi({open_n35936,freqD[0]}),
    .f({_al_u1593_o,\PWMD/mux3_b0_sel_is_3_o }),
    .q({open_n35941,\PWMD/FreCntr [0]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~(~D*B)*~(~C*A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1111010100110001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1595|PWMD/reg0_b12  (
    .a({\PWMD/FreCnt [12],open_n35942}),
    .b({\PWMD/FreCnt [15],\PWMD/n12 [12]}),
    .c({\PWMD/FreCntr [12],freqD[12]}),
    .clk(clk100m),
    .d({\PWMD/FreCntr [15],\PWMD/n0_lutinv }),
    .sr(\PWMD/n11 ),
    .f({_al_u1595_o,open_n35956}),
    .q({open_n35960,\PWMD/FreCnt [12]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*A*~(D@C))"),
    //.LUTF1("(C*B*A*~(0@D))"),
    //.LUTG0("(B*A*~(D@C))"),
    //.LUTG1("(C*B*A*~(1@D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000000000001000),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b1000000000001000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1596|PWMD/reg1_b21  (
    .a({_al_u1592_o,_al_u2810_o}),
    .b({_al_u1594_o,_al_u2811_o}),
    .c({_al_u1595_o,\PWMD/FreCnt [20]}),
    .ce(\PWMD/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMD/FreCnt [21],\PWMD/FreCntr [21]}),
    .e({\PWMD/FreCntr [21],open_n35961}),
    .mi({open_n35963,freqD[21]}),
    .f({_al_u1596_o,_al_u2812_o}),
    .q({open_n35979,\PWMD/FreCntr [21]}));  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(A*~(0@C)*~(D@B))"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(A*~(1@C)*~(D@B))"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000100000000010),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b1000000000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1598|_al_u2741  (
    .a({_al_u1597_o,_al_u2740_o}),
    .b({\PWMD/FreCnt [11],pnumcntD[21]}),
    .c({\PWMD/FreCnt [25],pnumcntD[22]}),
    .d({\PWMD/FreCntr [11],pnumcntD[23]}),
    .e({\PWMD/FreCntr [25],pnumcntD[2]}),
    .f({_al_u1598_o,_al_u2741_o}));
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(D@B)*~(C@A))"),
    //.LUTF1("(A*~(0@C)*~(D@B))"),
    //.LUTG0("(~(D@B)*~(C@A))"),
    //.LUTG1("(A*~(1@C)*~(D@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000010000100001),
    .INIT_LUTF1(16'b0000100000000010),
    .INIT_LUTG0(16'b1000010000100001),
    .INIT_LUTG1(16'b1000000000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1600|PWMD/reg1_b3  (
    .a({_al_u1599_o,\PWMD/FreCnt [2]}),
    .b({\PWMD/FreCnt [1],\PWMD/FreCnt [3]}),
    .c({\PWMD/FreCnt [10],\PWMD/FreCntr [2]}),
    .ce(\PWMD/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWMD/FreCntr [1],\PWMD/FreCntr [3]}),
    .e({\PWMD/FreCntr [10],open_n36002}),
    .mi({open_n36004,freqD[3]}),
    .f({_al_u1600_o,_al_u1599_o}),
    .q({open_n36020,\PWMD/FreCntr [3]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1602|PWME/reg1_b8  (
    .a({\PWME/FreCnt [22],_al_u1602_o}),
    .b({\PWME/FreCnt [23],\PWME/FreCnt [17]}),
    .c({\PWME/FreCntr [22],\PWME/FreCnt [8]}),
    .ce(\PWME/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWME/FreCntr [23],\PWME/FreCntr [17]}),
    .e({open_n36021,\PWME/FreCntr [8]}),
    .mi({open_n36023,freqE[8]}),
    .f({_al_u1602_o,_al_u1603_o}),
    .q({open_n36039,\PWME/FreCntr [8]}));  // src/OnePWM.v(37)
  // src/AHB.v(61)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(C*B*A*~(0@D))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(C*B*A*~(1@D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1607|U_AHB/reg15_b9  (
    .a({_al_u1603_o,_al_u1604_o}),
    .b({_al_u1605_o,\PWME/FreCnt [11]}),
    .c({_al_u1606_o,\PWME/FreCnt [9]}),
    .ce(\U_AHB/n32 ),
    .clk(clk100m),
    .d({\PWME/FreCnt [4],\PWME/FreCntr [11]}),
    .e({\PWME/FreCntr [4],\PWME/FreCntr [9]}),
    .mi({open_n36041,\U_AHB/h2h_hwdata [9]}),
    .f({_al_u1607_o,_al_u1605_o}),
    .q({open_n36057,freqE[9]}));  // src/AHB.v(61)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*B*A*~(0@D))"),
    //.LUTF1("(~(D*~B)*~(C*~A))"),
    //.LUTG0("(C*B*A*~(1@D))"),
    //.LUTG1("(~(D*~B)*~(C*~A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b1000110010101111),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b1000110010101111),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1608|PWME/reg1_b12  (
    .a({\PWME/FreCnt [12],_al_u2884_o}),
    .b({\PWME/FreCnt [15],_al_u2886_o}),
    .c({\PWME/FreCntr [12],_al_u2887_o}),
    .ce(\PWME/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWME/FreCntr [15],\PWME/FreCnt [11]}),
    .e({open_n36058,\PWME/FreCntr [12]}),
    .mi({open_n36060,freqE[12]}),
    .f({_al_u1608_o,_al_u2888_o}),
    .q({open_n36076,\PWME/FreCntr [12]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(B*A*~(D@C))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1000000000001000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1610|PWME/reg0_b2  (
    .a({_al_u1608_o,open_n36077}),
    .b({_al_u1609_o,\PWME/n12 [2]}),
    .c({\PWME/FreCnt [21],freqE[2]}),
    .clk(clk100m),
    .d({\PWME/FreCntr [21],\PWME/n0_lutinv }),
    .sr(\PWME/n11 ),
    .f({_al_u1610_o,open_n36091}),
    .q({open_n36095,\PWME/FreCnt [2]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(D@B)*~(C@A))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(~(D@B)*~(C@A))"),
    //.LUTG1("(C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000010000100001),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b1000010000100001),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1611|PWME/reg1_b1  (
    .a({open_n36096,\PWME/FreCnt [0]}),
    .b({open_n36097,\PWME/FreCnt [14]}),
    .c({\PWME/FreCntr [1],\PWME/FreCntr [1]}),
    .ce(\PWME/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWME/FreCnt [1],\PWME/FreCntr [15]}),
    .mi({open_n36101,freqE[1]}),
    .f({_al_u1611_o,_al_u2879_o}),
    .q({open_n36117,\PWME/FreCntr [1]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*D)"),
    //.LUTF1("(C*B*A*~(0@D))"),
    //.LUTG0("(C*D)"),
    //.LUTG1("(C*B*A*~(1@D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000000000000),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b1111000000000000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1614|PWME/reg1_b0  (
    .a({_al_u1610_o,open_n36118}),
    .b({_al_u1612_o,open_n36119}),
    .c({_al_u1613_o,\PWME/n11 }),
    .ce(\PWME/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWME/FreCnt [0],\PWME/n0_lutinv }),
    .e({\PWME/FreCntr [0],open_n36120}),
    .mi({open_n36122,freqE[0]}),
    .f({_al_u1614_o,\PWME/mux3_b0_sel_is_3_o }),
    .q({open_n36138,\PWME/FreCntr [0]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1615|PWME/reg1_b20  (
    .a({\PWME/FreCnt [14],_al_u1615_o}),
    .b({\PWME/FreCnt [25],\PWME/FreCnt [20]}),
    .c({\PWME/FreCntr [14],\PWME/FreCnt [26]}),
    .ce(\PWME/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWME/FreCntr [25],\PWME/FreCntr [20]}),
    .e({open_n36139,\PWME/FreCntr [26]}),
    .mi({open_n36141,freqE[20]}),
    .f({_al_u1615_o,_al_u1616_o}),
    .q({open_n36157,\PWME/FreCntr [20]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~(D@B)*~(C@A))"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~(D@B)*~(C@A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1000010000100001),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1000010000100001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1617|PWME/reg0_b13  (
    .a({\PWME/FreCnt [13],open_n36158}),
    .b({\PWME/FreCnt [16],\PWME/n12 [13]}),
    .c({\PWME/FreCntr [13],freqE[13]}),
    .clk(clk100m),
    .d({\PWME/FreCntr [16],\PWME/n0_lutinv }),
    .sr(\PWME/n11 ),
    .f({_al_u1617_o,open_n36176}),
    .q({open_n36180,\PWME/FreCnt [13]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(A*~(0@C)*~(D@B))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(A*~(1@C)*~(D@B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b0000100000000010),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000000000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1618|PWME/reg1_b19  (
    .a({_al_u1617_o,_al_u2891_o}),
    .b(\PWME/FreCnt [19:18]),
    .c({\PWME/FreCnt [2],\PWME/FreCnt [25]}),
    .ce(\PWME/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWME/FreCntr [19],\PWME/FreCntr [19]}),
    .e({\PWME/FreCntr [2],\PWME/FreCntr [26]}),
    .mi({open_n36182,freqE[19]}),
    .f({_al_u1618_o,_al_u2892_o}),
    .q({open_n36198,\PWME/FreCntr [19]}));  // src/OnePWM.v(37)
  // src/AHB.v(62)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~D*B)*~(~C*A))"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(~(~D*B)*~(~C*A))"),
    //.LUTG1("(C*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111010100110001),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b1111010100110001),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1629|U_AHB/reg16_b1  (
    .a({open_n36199,\PWMF/FreCnt [1]}),
    .b({open_n36200,\PWMF/FreCnt [15]}),
    .c({\PWMF/FreCntr [1],\PWMF/FreCntr [1]}),
    .ce(\U_AHB/n34 ),
    .clk(clk100m),
    .d({\PWMF/FreCnt [1],\PWMF/FreCntr [15]}),
    .mi({open_n36204,\U_AHB/h2h_hwdata [1]}),
    .f({_al_u1629_o,_al_u1631_o}),
    .q({open_n36220,freqF[1]}));  // src/AHB.v(62)
  // src/AHB.v(62)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~A*~(0@C)*~(~D*B))"),
    //.LUTF1("(C*B*A*~(0@D))"),
    //.LUTG0("(~A*~(1@C)*~(~D*B))"),
    //.LUTG1("(C*B*A*~(1@D))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010100000001),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b0101000000010000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1632|U_AHB/reg16_b12  (
    .a({_al_u1628_o,_al_u1629_o}),
    .b({_al_u1630_o,\PWMF/FreCnt [12]}),
    .c({_al_u1631_o,\PWMF/FreCnt [24]}),
    .ce(\U_AHB/n34 ),
    .clk(clk100m),
    .d({\PWMF/FreCnt [0],\PWMF/FreCntr [12]}),
    .e({\PWMF/FreCntr [0],\PWMF/FreCntr [24]}),
    .mi({open_n36222,\U_AHB/h2h_hwdata [12]}),
    .f({_al_u1632_o,_al_u1630_o}),
    .q({open_n36238,freqF[12]}));  // src/AHB.v(62)
  // src/AHB.v(60)
  EF2_PHY_MSLICE #(
    //.LUT0("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    //.LUT1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101001101011111),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1686|U_AHB/reg14_b6  (
    .a({pnumcnt0[18],pnumcnt0[19]}),
    .b({pnumcnt0[19],pnumcnt1[19]}),
    .c({pnumcnt0[1],\U_AHB/h2h_haddr [2]}),
    .ce(\U_AHB/n30 ),
    .clk(clk100m),
    .d({pnumcnt0[20],\U_AHB/h2h_haddr [3]}),
    .mi({open_n36249,\U_AHB/h2h_hwdata [6]}),
    .f({_al_u1686_o,_al_u3222_o}),
    .q({open_n36254,freqD[6]}));  // src/AHB.v(60)
  EF2_PHY_MSLICE #(
    //.LUT0("(~0*~D*~C*~B*A)"),
    //.LUT1("(~1*~D*~C*~B*A)"),
    .INIT_LUT0(16'b0000000000000010),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1687 (
    .a({_al_u1686_o,_al_u1686_o}),
    .b({pnumcnt0[21],pnumcnt0[21]}),
    .c({pnumcnt0[22],pnumcnt0[22]}),
    .d({pnumcnt0[23],pnumcnt0[23]}),
    .mi({open_n36267,pnumcnt0[2]}),
    .fx({open_n36272,_al_u1687_o}));
  EF2_PHY_MSLICE #(
    //.LUT0("(~0*~D*~C*~B*A)"),
    //.LUT1("(~1*~D*~C*~B*A)"),
    .INIT_LUT0(16'b0000000000000010),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1688 (
    .a({_al_u1687_o,_al_u1687_o}),
    .b({pnumcnt0[6],pnumcnt0[6]}),
    .c({pnumcnt0[7],pnumcnt0[7]}),
    .d({pnumcnt0[8],pnumcnt0[8]}),
    .mi({open_n36287,pnumcnt0[9]}),
    .fx({open_n36292,_al_u1688_o}));
  // src/AHB.v(60)
  EF2_PHY_MSLICE #(
    //.LUT0("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    //.LUT1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101001101011111),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1689|U_AHB/reg14_b2  (
    .a({pnumcnt0[10],pnumcnt0[13]}),
    .b({pnumcnt0[11],pnumcnt1[13]}),
    .c({pnumcnt0[12],\U_AHB/h2h_haddr [2]}),
    .ce(\U_AHB/n30 ),
    .clk(clk100m),
    .d({pnumcnt0[13],\U_AHB/h2h_haddr [3]}),
    .mi({open_n36305,\U_AHB/h2h_hwdata [2]}),
    .f({_al_u1689_o,_al_u3288_o}),
    .q({open_n36310,freqD[2]}));  // src/AHB.v(60)
  // src/OnePWM.v(15)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u1690|PWM0/stopreq_reg  (
    .a({_al_u1689_o,open_n36311}),
    .b({pnumcnt0[14],open_n36312}),
    .c({pnumcnt0[15],\PWM0/stopreq }),
    .clk(clk100m),
    .d({pnumcnt0[16],\PWM0/n0_lutinv }),
    .e({pnumcnt0[17],open_n36314}),
    .sr(pwm_start_stop[0]),
    .f({_al_u1690_o,open_n36329}),
    .q({open_n36333,\PWM0/stopreq_keep }));  // src/OnePWM.v(15)
  // src/AHB.v(61)
  EF2_PHY_MSLICE #(
    //.LUT0("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    //.LUT1("(~C*~B*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101001101011111),
    .INIT_LUT1(16'b0000000000000011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1691|U_AHB/reg15_b20  (
    .a({open_n36334,pnumcnt0[5]}),
    .b({pnumcnt0[4],pnumcnt1[5]}),
    .c({pnumcnt0[5],\U_AHB/h2h_haddr [2]}),
    .ce(\U_AHB/n32 ),
    .clk(clk100m),
    .d({pnumcnt0[3],\U_AHB/h2h_haddr [3]}),
    .mi({open_n36345,\U_AHB/h2h_hwdata [20]}),
    .f({_al_u1691_o,_al_u3133_o}),
    .q({open_n36350,freqE[20]}));  // src/AHB.v(61)
  // src/AHB.v(80)
  EF2_PHY_LSLICE #(
    //.LUTF0("(D*~C*B*A)"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(D*~C*B*A)"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000000),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0000100000000000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1756|U_AHB/reg31_b31  (
    .a({_al_u1750_o,timer[22]}),
    .b({_al_u1752_o,timer[23]}),
    .c({_al_u1754_o,timer[26]}),
    .clk(clk100m),
    .d({_al_u1755_o,timer[27]}),
    .mi({open_n36355,\U_AHB/h2h_hwdata [31]}),
    .sr(\U_AHB/n73 ),
    .f({_al_u1756_o,_al_u1649_o}),
    .q({open_n36370,pnumD[31]}));  // src/AHB.v(80)
  // src/AHB.v(81)
  EF2_PHY_LSLICE #(
    //.LUTF0("(D*~C*B*A)"),
    //.LUTF1("(0*D*C*B*A)"),
    //.LUTG0("(D*~C*B*A)"),
    //.LUTG1("(1*D*C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000100000000000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1765|U_AHB/reg32_b31  (
    .a({_al_u1748_o,timer[12]}),
    .b({_al_u1756_o,timer[13]}),
    .c({_al_u1760_o,timer[16]}),
    .clk(clk100m),
    .d({_al_u1762_o,timer[17]}),
    .e({_al_u1764_o,open_n36372}),
    .mi({open_n36374,\U_AHB/h2h_hwdata [31]}),
    .sr(\U_AHB/n75 ),
    .f({_al_u1765_o,_al_u1643_o}),
    .q({open_n36389,pnumE[31]}));  // src/AHB.v(81)
  // CPLD_SOC_AHB_TOP.v(49)
  EF2_PHY_MSLICE #(
    //.LUT0("~(C*~(~B*~(~D*A)))"),
    //.LUT1("(~D*~C*~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0011111100011111),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \_al_u1768|reg1_b1  (
    .a({pnumcnt1[18],_al_u3055_o}),
    .b({pnumcnt1[19],_al_u2983_o}),
    .c({pnumcnt1[1],n4_neg}),
    .clk(clk25m),
    .d({pnumcnt1[20],ledout_pad[1]}),
    .sr(rst_n_pad),
    .f({_al_u1768_o,open_n36403}),
    .q({open_n36407,ledout_pad[1]}));  // CPLD_SOC_AHB_TOP.v(49)
  EF2_PHY_MSLICE #(
    //.LUT0("(~0*~D*~C*~B*A)"),
    //.LUT1("(~1*~D*~C*~B*A)"),
    .INIT_LUT0(16'b0000000000000010),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1769 (
    .a({_al_u1768_o,_al_u1768_o}),
    .b({pnumcnt1[21],pnumcnt1[21]}),
    .c({pnumcnt1[22],pnumcnt1[22]}),
    .d({pnumcnt1[23],pnumcnt1[23]}),
    .mi({open_n36420,pnumcnt1[2]}),
    .fx({open_n36425,_al_u1769_o}));
  // src/AHB.v(84)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~(D*C*B*A))"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(~1*~(D*C*B*A))"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111111111111111),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1770|U_AHB/reg34_b1  (
    .a({_al_u1769_o,_al_u1770_o}),
    .b({pnumcnt1[6],_al_u1772_o}),
    .c({pnumcnt1[7],_al_u1773_o}),
    .clk(clk100m),
    .d({pnumcnt1[8],pnumcnt1[0]}),
    .e({pnumcnt1[9],\PWM1/stopreq }),
    .mi({open_n36430,\U_AHB/h2h_hwdata [1]}),
    .sr(\U_AHB/n79 ),
    .f({_al_u1770_o,_al_u3010_o}),
    .q({open_n36445,pwm_start_stop[1]}));  // src/AHB.v(84)
  // src/AHB.v(68)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUT1("(~D*~C*~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1010100000100000),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1771|U_AHB/reg19_b2  (
    .a({pnumcnt1[10],\PWM1/n24 }),
    .b({pnumcnt1[11],\PWM1/n25_neg_lutinv }),
    .c({pnumcnt1[12],\PWM1/n26 [2]}),
    .clk(clk100m),
    .d({pnumcnt1[13],\PWM1/pnumr [2]}),
    .mi({open_n36457,\U_AHB/h2h_hwdata [2]}),
    .sr(\U_AHB/n47 ),
    .f({_al_u1771_o,_al_u1797_o}),
    .q({open_n36461,pnum1[2]}));  // src/AHB.v(68)
  EF2_PHY_MSLICE #(
    //.LUT0("(~0*~D*~C*~B*A)"),
    //.LUT1("(~1*~D*~C*~B*A)"),
    .INIT_LUT0(16'b0000000000000010),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1772 (
    .a({_al_u1771_o,_al_u1771_o}),
    .b({pnumcnt1[14],pnumcnt1[14]}),
    .c({pnumcnt1[15],pnumcnt1[15]}),
    .d({pnumcnt1[16],pnumcnt1[16]}),
    .mi({open_n36474,pnumcnt1[17]}),
    .fx({open_n36479,_al_u1772_o}));
  // src/AHB.v(61)
  EF2_PHY_MSLICE #(
    //.LUT0("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    //.LUT1("(~C*~B*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101001101011111),
    .INIT_LUT1(16'b0000000000000011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1773|U_AHB/reg15_b19  (
    .a({open_n36482,pnumcnt0[4]}),
    .b({pnumcnt1[4],pnumcnt1[4]}),
    .c({pnumcnt1[5],\U_AHB/h2h_haddr [2]}),
    .ce(\U_AHB/n32 ),
    .clk(clk100m),
    .d({pnumcnt1[3],\U_AHB/h2h_haddr [3]}),
    .mi({open_n36493,\U_AHB/h2h_hwdata [19]}),
    .f({_al_u1773_o,_al_u3145_o}),
    .q({open_n36498,freqE[19]}));  // src/AHB.v(61)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~A*~(0@C)*~(~D*B))"),
    //.LUTF1("(0*D*C*B*A)"),
    //.LUTG0("(~A*~(1@C)*~(~D*B))"),
    //.LUTG1("(1*D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000010100000001),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0101000000010000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1838|PWM1/reg1_b21  (
    .a({_al_u1829_o,_al_u1836_o}),
    .b({_al_u1831_o,\PWM1/FreCnt [15]}),
    .c({_al_u1833_o,\PWM1/FreCnt [20]}),
    .ce(\PWM1/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({_al_u1835_o,\PWM1/FreCntr [16]}),
    .e({_al_u1837_o,\PWM1/FreCntr [21]}),
    .mi({open_n36500,freq1[21]}),
    .f({_al_u1838_o,_al_u1837_o}),
    .q({open_n36516,\PWM1/FreCntr [21]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(D*~(C@B))"),
    //.LUTF1("(0*D*C*B*A)"),
    //.LUTG0("(D*~(C@B))"),
    //.LUTG1("(1*D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100001100000000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1100001100000000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1847|PWM1/reg1_b3  (
    .a({_al_u1838_o,open_n36517}),
    .b({_al_u1840_o,\PWM1/FreCnt [2]}),
    .c({_al_u1842_o,\PWM1/FreCntr [3]}),
    .ce(\PWM1/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({_al_u1844_o,_al_u1841_o}),
    .e({_al_u1846_o,open_n36518}),
    .mi({open_n36520,freq1[3]}),
    .f({_al_u1847_o,_al_u1842_o}),
    .q({open_n36536,\PWM1/FreCntr [3]}));  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~D*~C*~B*~A)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(~D*~C*~B*~A)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .INIT_LUTF0(16'b0000000000000001),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000000000000001),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1850|_al_u1930  (
    .a({pnumcnt2[18],pnumcnt3[18]}),
    .b({pnumcnt2[19],pnumcnt3[19]}),
    .c({pnumcnt2[1],pnumcnt3[1]}),
    .d({pnumcnt2[20],pnumcnt3[20]}),
    .f({_al_u1850_o,_al_u1930_o}));
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1851|_al_u1852  (
    .a({_al_u1850_o,_al_u1851_o}),
    .b({pnumcnt2[21],pnumcnt2[6]}),
    .c({pnumcnt2[22],pnumcnt2[7]}),
    .d({pnumcnt2[23],pnumcnt2[8]}),
    .e({pnumcnt2[2],pnumcnt2[9]}),
    .f({_al_u1851_o,_al_u1852_o}));
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1853|_al_u1854  (
    .a({pnumcnt2[10],_al_u1853_o}),
    .b({pnumcnt2[11],pnumcnt2[14]}),
    .c({pnumcnt2[12],pnumcnt2[15]}),
    .d({pnumcnt2[13],pnumcnt2[16]}),
    .e({open_n36585,pnumcnt2[17]}),
    .f({_al_u1853_o,_al_u1854_o}));
  // src/OnePWM.v(15)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(~C*~B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000000000000011),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u1855|PWM2/stopreq_reg  (
    .b({pnumcnt2[4],open_n36608}),
    .c({pnumcnt2[5],\PWM2/stopreq }),
    .clk(clk100m),
    .d({pnumcnt2[3],\PWM2/n0_lutinv }),
    .sr(pwm_start_stop[2]),
    .f({_al_u1855_o,open_n36622}),
    .q({open_n36626,\PWM2/stopreq_keep }));  // src/OnePWM.v(15)
  // src/AHB.v(78)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~(D*C*B*A))"),
    //.LUTF1("(~D*C*B*A)"),
    //.LUTG0("(~1*~(D*C*B*A))"),
    //.LUTG1("(~D*C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111111111111111),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1856|U_AHB/reg29_b27  (
    .a({_al_u1852_o,_al_u1852_o}),
    .b({_al_u1854_o,_al_u1854_o}),
    .c({_al_u1855_o,_al_u1855_o}),
    .clk(clk100m),
    .d({pnumcnt2[0],pnumcnt2[0]}),
    .e({open_n36628,\PWM2/stopreq }),
    .mi({open_n36630,\U_AHB/h2h_hwdata [27]}),
    .sr(\U_AHB/n69 ),
    .f({\PWM2/n25_neg_lutinv ,_al_u3013_o}),
    .q({open_n36645,pnumB[27]}));  // src/AHB.v(78)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1903|PWM2/reg2_b27  (
    .a({\PWM2/n24 ,\PWM2/pnumr [27]}),
    .b({\PWM2/n25_neg_lutinv ,pnum2[27]}),
    .c({\PWM2/n26 [0],pnum2[32]}),
    .clk(clk100m),
    .d({\PWM2/pnumr [0],pwm_start_stop[18]}),
    .f({_al_u1903_o,open_n36660}),
    .q({open_n36664,\PWM2/pnumr[27]_keep }));  // src/OnePWM.v(48)
  // src/AHB.v(64)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1101110011110000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1927|U_AHB/reg17_b29  (
    .a({_al_u1921_o,\U_AHB/n38 }),
    .b({_al_u1923_o,\U_AHB/n36 }),
    .c({_al_u1925_o,gpio_out_pad[29]}),
    .clk(clk100m),
    .d({_al_u1926_o,\U_AHB/h2h_hwdata [29]}),
    .f({_al_u1927_o,open_n36679}),
    .q({open_n36683,gpio_out_pad[29]}));  // src/AHB.v(64)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1931|_al_u2095  (
    .a({_al_u1930_o,_al_u2094_o}),
    .b({pnumcnt3[21],pnumcnt5[21]}),
    .c({pnumcnt3[22],pnumcnt5[22]}),
    .d({pnumcnt3[23],pnumcnt5[23]}),
    .e({pnumcnt3[2],pnumcnt5[2]}),
    .f({_al_u1931_o,_al_u2095_o}));
  EF2_PHY_MSLICE #(
    //.LUT0("(~0*~D*~C*~B*A)"),
    //.LUT1("(~1*~D*~C*~B*A)"),
    .INIT_LUT0(16'b0000000000000010),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1932 (
    .a({_al_u1931_o,_al_u1931_o}),
    .b({pnumcnt3[6],pnumcnt3[6]}),
    .c({pnumcnt3[7],pnumcnt3[7]}),
    .d({pnumcnt3[8],pnumcnt3[8]}),
    .mi({open_n36718,pnumcnt3[9]}),
    .fx({open_n36723,_al_u1932_o}));
  EF2_PHY_LSLICE #(
    //.LUTF0("(~D*~C*~B*~A)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(~D*~C*~B*~A)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .INIT_LUTF0(16'b0000000000000001),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000000000000001),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u1933|_al_u2097  (
    .a({pnumcnt3[10],pnumcnt5[10]}),
    .b({pnumcnt3[11],pnumcnt5[11]}),
    .c({pnumcnt3[12],pnumcnt5[12]}),
    .d({pnumcnt3[13],pnumcnt5[13]}),
    .f({_al_u1933_o,_al_u2097_o}));
  EF2_PHY_MSLICE #(
    //.LUT0("(~0*~D*~C*~B*A)"),
    //.LUT1("(~1*~D*~C*~B*A)"),
    .INIT_LUT0(16'b0000000000000010),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u1934 (
    .a({_al_u1933_o,_al_u1933_o}),
    .b({pnumcnt3[14],pnumcnt3[14]}),
    .c({pnumcnt3[15],pnumcnt3[15]}),
    .d({pnumcnt3[16],pnumcnt3[16]}),
    .mi({open_n36762,pnumcnt3[17]}),
    .fx({open_n36767,_al_u1934_o}));
  // src/OnePWM.v(15)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(~C*~B*~D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(~C*~B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000000000000011),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000000000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u1935|PWM3/stopreq_reg  (
    .b({pnumcnt3[4],open_n36772}),
    .c({pnumcnt3[5],\PWM3/stopreq }),
    .clk(clk100m),
    .d({pnumcnt3[3],\PWM3/n0_lutinv }),
    .sr(pwm_start_stop[3]),
    .f({_al_u1935_o,open_n36790}),
    .q({open_n36794,\PWM3/stopreq_keep }));  // src/OnePWM.v(15)
  // src/AHB.v(78)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~(D*C*B*A))"),
    //.LUTF1("(~D*C*B*A)"),
    //.LUTG0("(~1*~(D*C*B*A))"),
    //.LUTG1("(~D*C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111111111111111),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u1936|U_AHB/reg29_b25  (
    .a({_al_u1932_o,_al_u1932_o}),
    .b({_al_u1934_o,_al_u1934_o}),
    .c({_al_u1935_o,_al_u1935_o}),
    .clk(clk100m),
    .d({pnumcnt3[0],pnumcnt3[0]}),
    .e({open_n36796,\PWM3/stopreq }),
    .mi({open_n36798,\U_AHB/h2h_hwdata [25]}),
    .sr(\U_AHB/n69 ),
    .f({\PWM3/n25_neg_lutinv ,_al_u3016_o}),
    .q({open_n36813,pnumB[25]}));  // src/AHB.v(78)
  // src/OnePWM.v(58)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1010100000100000),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1010100000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1983|PWM3/reg3_b0  (
    .a({\PWM3/n24 ,_al_u1983_o}),
    .b({\PWM3/n25_neg_lutinv ,\PWM3/n24 }),
    .c({\PWM3/n26 [0],pnumcnt3[0]}),
    .clk(clk100m),
    .d({\PWM3/pnumr [0],\PWM3/pnumr [0]}),
    .e({open_n36815,pwm_start_stop[19]}),
    .f({_al_u1983_o,open_n36831}),
    .q({open_n36835,\PWM3/RemaTxNum[0]_keep }));  // src/OnePWM.v(58)
  // src/AHB.v(49)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(~0*C)*~(D*~B))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(A*~(~1*C)*~(D*~B))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000001010),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b1000100010101010),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u1992|U_AHB/reg4_b13  (
    .a({_al_u1986_o,_al_u1989_o}),
    .b({_al_u1988_o,\PWM3/FreCnt [12]}),
    .c({_al_u1990_o,\PWM3/FreCnt [25]}),
    .ce(\U_AHB/n10 ),
    .clk(clk100m),
    .d({_al_u1991_o,\PWM3/FreCntr [13]}),
    .e({open_n36836,\PWM3/FreCntr [26]}),
    .mi({open_n36838,\U_AHB/h2h_hwdata [13]}),
    .f({_al_u1992_o,_al_u1990_o}),
    .q({open_n36854,freq3[13]}));  // src/AHB.v(49)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(D*~(C@B))"),
    //.LUT1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100001100000000),
    .INIT_LUT1(16'b1100000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2000|PWM3/reg1_b3  (
    .b({_al_u1997_o,\PWM3/FreCnt [2]}),
    .c({_al_u1999_o,\PWM3/FreCntr [3]}),
    .ce(\PWM3/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({_al_u1995_o,_al_u1985_o}),
    .mi({open_n36867,freq3[3]}),
    .f({_al_u2000_o,_al_u1986_o}),
    .q({open_n36872,\PWM3/FreCntr [3]}));  // src/OnePWM.v(37)
  // src/AHB.v(78)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(0*D*C*B*A)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(1*D*C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2009|U_AHB/reg29_b26  (
    .a({_al_u1992_o,open_n36873}),
    .b({_al_u2000_o,open_n36874}),
    .c({_al_u2004_o,pwm_state_read[3]}),
    .clk(clk100m),
    .d({_al_u2006_o,_al_u2009_o}),
    .e({_al_u2008_o,open_n36876}),
    .mi({open_n36878,\U_AHB/h2h_hwdata [26]}),
    .sr(\U_AHB/n69 ),
    .f({_al_u2009_o,\PWM3/u14_sel_is_1_o }),
    .q({open_n36893,pnumB[26]}));  // src/AHB.v(78)
  // src/AHB.v(50)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2012|U_AHB/reg5_b24  (
    .a({pnumcnt4[18],_al_u3234_o}),
    .b({pnumcnt4[19],\U_AHB/n96 }),
    .c({pnumcnt4[1],\U_AHB/n93 }),
    .ce(\U_AHB/n12 ),
    .clk(clk100m),
    .d({pnumcnt4[20],pnumcnt4[18]}),
    .e({open_n36894,pnumcnt5[18]}),
    .mi({open_n36896,\U_AHB/h2h_hwdata [24]}),
    .f({_al_u2012_o,_al_u3235_o}),
    .q({open_n36912,freq4[24]}));  // src/AHB.v(50)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2013|_al_u2014  (
    .a({_al_u2012_o,_al_u2013_o}),
    .b({pnumcnt4[21],pnumcnt4[6]}),
    .c({pnumcnt4[22],pnumcnt4[7]}),
    .d({pnumcnt4[23],pnumcnt4[8]}),
    .e({pnumcnt4[2],pnumcnt4[9]}),
    .f({_al_u2013_o,_al_u2014_o}));
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2015|_al_u2016  (
    .a({pnumcnt4[10],_al_u2015_o}),
    .b({pnumcnt4[11],pnumcnt4[14]}),
    .c({pnumcnt4[12],pnumcnt4[15]}),
    .d({pnumcnt4[13],pnumcnt4[16]}),
    .e({open_n36937,pnumcnt4[17]}),
    .f({_al_u2015_o,_al_u2016_o}));
  // src/OnePWM.v(15)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(~C*~B*~D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(~C*~B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000000000000011),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000000000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2017|PWM4/stopreq_reg  (
    .b({pnumcnt4[4],open_n36960}),
    .c({pnumcnt4[5],\PWM4/stopreq }),
    .clk(clk100m),
    .d({pnumcnt4[3],\PWM4/n0_lutinv }),
    .sr(pwm_start_stop[4]),
    .f({_al_u2017_o,open_n36978}),
    .q({open_n36982,\PWM4/stopreq_keep }));  // src/OnePWM.v(15)
  // src/AHB.v(77)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~(D*C*B*A))"),
    //.LUTF1("(~D*C*B*A)"),
    //.LUTG0("(~1*~(D*C*B*A))"),
    //.LUTG1("(~D*C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111111111111111),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2018|U_AHB/reg28_b9  (
    .a({_al_u2014_o,_al_u2014_o}),
    .b({_al_u2016_o,_al_u2016_o}),
    .c({_al_u2017_o,_al_u2017_o}),
    .clk(clk100m),
    .d({pnumcnt4[0],pnumcnt4[0]}),
    .e({open_n36984,\PWM4/stopreq }),
    .mi({open_n36986,\U_AHB/h2h_hwdata [9]}),
    .sr(\U_AHB/n67 ),
    .f({\PWM4/n25_neg_lutinv ,_al_u3019_o}),
    .q({open_n37001,pnumA[9]}));  // src/AHB.v(77)
  // src/AHB.v(50)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~D*~C*~B*A)"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(~D*~C*~B*A)"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b0000000000000010),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2075|U_AHB/reg5_b8  (
    .a({open_n37002,_al_u883_o}),
    .b({_al_u2072_o,\PWM4/FreCnt [7]}),
    .c({_al_u2074_o,\PWM4/FreCnt [8]}),
    .ce(\U_AHB/n12 ),
    .clk(clk100m),
    .d({_al_u2070_o,\PWM4/FreCnt [9]}),
    .mi({open_n37006,\U_AHB/h2h_hwdata [8]}),
    .f({_al_u2075_o,_al_u884_o}),
    .q({open_n37022,freq4[8]}));  // src/AHB.v(50)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~C*~(0*~B)*~(D@A))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~C*~(1*~B)*~(D@A))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101000000101),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0000100000000100),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2083|PWM4/reg1_b11  (
    .a({_al_u2077_o,\PWM4/FreCnt [10]}),
    .b({_al_u2079_o,\PWM4/FreCnt [25]}),
    .c({_al_u2081_o,\PWM4/FreCnt [26]}),
    .ce(\PWM4/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({_al_u2082_o,\PWM4/FreCntr [11]}),
    .e({open_n37023,\PWM4/FreCntr [26]}),
    .mi({open_n37025,freq4[11]}),
    .f({_al_u2083_o,_al_u2082_o}),
    .q({open_n37041,\PWM4/FreCntr [11]}));  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(0*D*C*B*A)"),
    //.LUT1("(1*D*C*B*A)"),
    .INIT_LUT0(16'b0000000000000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2091 (
    .a({_al_u2075_o,_al_u2075_o}),
    .b({_al_u2083_o,_al_u2083_o}),
    .c({_al_u2086_o,_al_u2086_o}),
    .d({_al_u2088_o,_al_u2088_o}),
    .mi({open_n37054,_al_u2090_o}),
    .fx({open_n37059,_al_u2091_o}));
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*A*~(D*~C))"),
    //.LUT1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000000010001000),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2094|PWM0/reg1_b24  (
    .a({pnumcnt5[18],_al_u1758_o}),
    .b({pnumcnt5[19],_al_u1759_o}),
    .c({pnumcnt5[1],\PWM0/FreCnt [23]}),
    .ce(\PWM0/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({pnumcnt5[20],\PWM0/FreCntr [24]}),
    .mi({open_n37072,freq0[24]}),
    .f({_al_u2094_o,_al_u1760_o}),
    .q({open_n37077,\PWM0/FreCntr [24]}));  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(~0*~D*~C*~B*A)"),
    //.LUT1("(~1*~D*~C*~B*A)"),
    .INIT_LUT0(16'b0000000000000010),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2096 (
    .a({_al_u2095_o,_al_u2095_o}),
    .b({pnumcnt5[6],pnumcnt5[6]}),
    .c({pnumcnt5[7],pnumcnt5[7]}),
    .d({pnumcnt5[8],pnumcnt5[8]}),
    .mi({open_n37090,pnumcnt5[9]}),
    .fx({open_n37095,_al_u2096_o}));
  EF2_PHY_MSLICE #(
    //.LUT0("(~0*~D*~C*~B*A)"),
    //.LUT1("(~1*~D*~C*~B*A)"),
    .INIT_LUT0(16'b0000000000000010),
    .INIT_LUT1(16'b0000000000000000),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u2098 (
    .a({_al_u2097_o,_al_u2097_o}),
    .b({pnumcnt5[14],pnumcnt5[14]}),
    .c({pnumcnt5[15],pnumcnt5[15]}),
    .d({pnumcnt5[16],pnumcnt5[16]}),
    .mi({open_n37110,pnumcnt5[17]}),
    .fx({open_n37115,_al_u2098_o}));
  // src/OnePWM.v(15)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(~C*~B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000000000000011),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2099|PWM5/stopreq_reg  (
    .b({pnumcnt5[4],open_n37120}),
    .c({pnumcnt5[5],\PWM5/stopreq }),
    .clk(clk100m),
    .d({pnumcnt5[3],\PWM5/n0_lutinv }),
    .sr(pwm_start_stop[5]),
    .f({_al_u2099_o,open_n37134}),
    .q({open_n37138,\PWM5/stopreq_keep }));  // src/OnePWM.v(15)
  // src/AHB.v(77)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~(D*C*B*A))"),
    //.LUTF1("(~D*C*B*A)"),
    //.LUTG0("(~1*~(D*C*B*A))"),
    //.LUTG1("(~D*C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111111111111111),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2100|U_AHB/reg28_b30  (
    .a({_al_u2096_o,_al_u2096_o}),
    .b({_al_u2098_o,_al_u2098_o}),
    .c({_al_u2099_o,_al_u2099_o}),
    .clk(clk100m),
    .d({pnumcnt5[0],pnumcnt5[0]}),
    .e({open_n37140,\PWM5/stopreq }),
    .mi({open_n37142,\U_AHB/h2h_hwdata [30]}),
    .sr(\U_AHB/n67 ),
    .f({\PWM5/n25_neg_lutinv ,_al_u3022_o}),
    .q({open_n37157,pnumA[30]}));  // src/AHB.v(77)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*A*~(~D*C))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000100000001000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2157|PWM5/reg1_b9  (
    .a({_al_u2150_o,_al_u2166_o}),
    .b({_al_u2152_o,_al_u2167_o}),
    .c({_al_u2154_o,\PWM5/FreCnt [8]}),
    .ce(\PWM5/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({_al_u2156_o,\PWM5/FreCntr [9]}),
    .mi({open_n37168,freq5[9]}),
    .f({_al_u2157_o,_al_u2168_o}),
    .q({open_n37173,\PWM5/FreCntr [9]}));  // src/OnePWM.v(37)
  // src/AHB.v(51)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(~D*C)*~(0*~B))"),
    //.LUTF1("(C*B*D)"),
    //.LUTG0("(A*~(~D*C)*~(1*~B))"),
    //.LUTG1("(C*B*D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1010101000001010),
    .INIT_LUTF1(16'b1100000000000000),
    .INIT_LUTG0(16'b1000100000001000),
    .INIT_LUTG1(16'b1100000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2164|U_AHB/reg6_b16  (
    .a({open_n37174,_al_u2158_o}),
    .b({_al_u2161_o,\PWM5/FreCnt [1]}),
    .c({_al_u2163_o,\PWM5/FreCnt [15]}),
    .ce(\U_AHB/n14 ),
    .clk(clk100m),
    .d({_al_u2159_o,\PWM5/FreCntr [16]}),
    .e({open_n37175,\PWM5/FreCntr [2]}),
    .mi({open_n37177,\U_AHB/h2h_hwdata [16]}),
    .f({_al_u2164_o,_al_u2159_o}),
    .q({open_n37193,freq5[16]}));  // src/AHB.v(51)
  // src/AHB.v(68)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2176|U_AHB/reg19_b26  (
    .a({pnumcnt6[18],_al_u3235_o}),
    .b({pnumcnt6[19],\U_AHB/n102 }),
    .c({pnumcnt6[1],\U_AHB/n99 }),
    .clk(clk100m),
    .d({pnumcnt6[20],pnumcnt6[18]}),
    .e({open_n37195,pnumcnt7[18]}),
    .mi({open_n37197,\U_AHB/h2h_hwdata [26]}),
    .sr(\U_AHB/n47 ),
    .f({_al_u2176_o,_al_u3236_o}),
    .q({open_n37212,pnum1[26]}));  // src/AHB.v(68)
  // src/AHB.v(68)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2177|U_AHB/reg19_b9  (
    .a({_al_u2176_o,_al_u3169_o}),
    .b({pnumcnt6[21],\U_AHB/n102 }),
    .c({pnumcnt6[22],\U_AHB/n99 }),
    .clk(clk100m),
    .d({pnumcnt6[23],pnumcnt6[23]}),
    .e({pnumcnt6[2],pnumcnt7[23]}),
    .mi({open_n37215,\U_AHB/h2h_hwdata [9]}),
    .sr(\U_AHB/n47 ),
    .f({_al_u2177_o,_al_u3170_o}),
    .q({open_n37230,pnum1[9]}));  // src/AHB.v(68)
  // src/AHB.v(69)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2178|U_AHB/reg20_b30  (
    .a({_al_u2177_o,_al_u3087_o}),
    .b({pnumcnt6[6],\U_AHB/n102 }),
    .c({pnumcnt6[7],\U_AHB/n99 }),
    .clk(clk100m),
    .d({pnumcnt6[8],pnumcnt6[9]}),
    .e({pnumcnt6[9],pnumcnt7[9]}),
    .mi({open_n37233,\U_AHB/h2h_hwdata [30]}),
    .sr(\U_AHB/n51 ),
    .f({_al_u2178_o,_al_u3089_o}),
    .q({open_n37248,pnum2[30]}));  // src/AHB.v(69)
  // src/AHB.v(67)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2179|U_AHB/reg18_b30  (
    .a({pnumcnt6[10],_al_u3290_o}),
    .b({pnumcnt6[11],\U_AHB/n102 }),
    .c({pnumcnt6[12],\U_AHB/n99 }),
    .clk(clk100m),
    .d({pnumcnt6[13],pnumcnt6[13]}),
    .e({open_n37250,pnumcnt7[13]}),
    .mi({open_n37252,\U_AHB/h2h_hwdata [30]}),
    .sr(\U_AHB/n45 ),
    .f({_al_u2179_o,_al_u3291_o}),
    .q({open_n37267,pnum0[30]}));  // src/AHB.v(67)
  // src/AHB.v(68)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2180|U_AHB/reg19_b25  (
    .a({_al_u2179_o,_al_u3246_o}),
    .b({pnumcnt6[14],\U_AHB/n102 }),
    .c({pnumcnt6[15],\U_AHB/n99 }),
    .clk(clk100m),
    .d({pnumcnt6[16],pnumcnt6[17]}),
    .e({pnumcnt6[17],pnumcnt7[17]}),
    .mi({open_n37270,\U_AHB/h2h_hwdata [25]}),
    .sr(\U_AHB/n47 ),
    .f({_al_u2180_o,_al_u3247_o}),
    .q({open_n37285,pnum1[25]}));  // src/AHB.v(68)
  // src/AHB.v(69)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(~C*~B*~D)"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(~C*~B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000000000000011),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000000000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2181|U_AHB/reg20_b26  (
    .a({open_n37286,_al_u3135_o}),
    .b({pnumcnt6[4],\U_AHB/n102 }),
    .c({pnumcnt6[5],\U_AHB/n99 }),
    .clk(clk100m),
    .d({pnumcnt6[3],pnumcnt6[5]}),
    .e({open_n37288,pnumcnt7[5]}),
    .mi({open_n37290,\U_AHB/h2h_hwdata [26]}),
    .sr(\U_AHB/n51 ),
    .f({_al_u2181_o,_al_u3136_o}),
    .q({open_n37305,pnum2[26]}));  // src/AHB.v(69)
  // src/AHB.v(67)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(~D*C*B*A)"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(~D*C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2182|U_AHB/reg18_b25  (
    .a({_al_u2178_o,_al_u3345_o}),
    .b({_al_u2180_o,\U_AHB/n102 }),
    .c({_al_u2181_o,\U_AHB/n99 }),
    .clk(clk100m),
    .d({pnumcnt6[0],pnumcnt6[0]}),
    .e({open_n37307,pnumcnt7[0]}),
    .mi({open_n37309,\U_AHB/h2h_hwdata [25]}),
    .sr(\U_AHB/n45 ),
    .f({\PWM6/n25_neg_lutinv ,_al_u3346_o}),
    .q({open_n37324,pnum0[25]}));  // src/AHB.v(67)
  EF2_PHY_SPAD #(
    //.LOCATION("P28"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u22 (
    .ipad(clkin),
    .ts(1'b1),
    .di(clkin_pad));  // CPLD_SOC_AHB_TOP.v(3)
  // src/AHB.v(73)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b1010100000100000),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b1010100000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2229|U_AHB/reg24_b26  (
    .a({\PWM6/n24 ,open_n37334}),
    .b({\PWM6/n25_neg_lutinv ,limit_l_pad[9]}),
    .c({\PWM6/n26 [0],limit_r_pad[9]}),
    .clk(clk100m),
    .d({\PWM6/pnumr [0],\PWM9/n11 }),
    .mi({open_n37339,\U_AHB/h2h_hwdata [26]}),
    .sr(\U_AHB/n59 ),
    .f({_al_u2229_o,_al_u3035_o}),
    .q({open_n37354,pnum6[26]}));  // src/AHB.v(73)
  // src/AHB.v(72)
  EF2_PHY_MSLICE #(
    //.LUT0("(~D*~C*~B*~A)"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000000000001),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2247|U_AHB/reg23_b29  (
    .a({_al_u2240_o,pnumcntA[10]}),
    .b({_al_u2242_o,pnumcntA[11]}),
    .c({_al_u2244_o,pnumcntA[12]}),
    .clk(clk100m),
    .d({_al_u2246_o,pnumcntA[13]}),
    .mi({open_n37366,\U_AHB/h2h_hwdata [29]}),
    .sr(\U_AHB/n57 ),
    .f({_al_u2247_o,_al_u2503_o}),
    .q({open_n37370,pnum5[29]}));  // src/AHB.v(72)
  // src/AHB.v(68)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2256|U_AHB/reg19_b29  (
    .a({pnumcnt7[18],_al_u3202_o}),
    .b({pnumcnt7[19],\U_AHB/n102 }),
    .c({pnumcnt7[1],\U_AHB/n99 }),
    .clk(clk100m),
    .d({pnumcnt7[20],pnumcnt6[20]}),
    .e({open_n37372,pnumcnt7[20]}),
    .mi({open_n37374,\U_AHB/h2h_hwdata [29]}),
    .sr(\U_AHB/n47 ),
    .f({_al_u2256_o,_al_u3203_o}),
    .q({open_n37389,pnum1[29]}));  // src/AHB.v(68)
  // src/AHB.v(68)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2257|U_AHB/reg19_b31  (
    .a({_al_u2256_o,_al_u3180_o}),
    .b({pnumcnt7[21],\U_AHB/n102 }),
    .c({pnumcnt7[22],\U_AHB/n99 }),
    .clk(clk100m),
    .d({pnumcnt7[23],pnumcnt6[22]}),
    .e({pnumcnt7[2],pnumcnt7[22]}),
    .mi({open_n37392,\U_AHB/h2h_hwdata [31]}),
    .sr(\U_AHB/n47 ),
    .f({_al_u2257_o,_al_u3181_o}),
    .q({open_n37407,pnum1[31]}));  // src/AHB.v(68)
  // src/AHB.v(69)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2258|U_AHB/reg20_b29  (
    .a({_al_u2257_o,_al_u3102_o}),
    .b({pnumcnt7[6],\U_AHB/n102 }),
    .c({pnumcnt7[7],\U_AHB/n99 }),
    .clk(clk100m),
    .d({pnumcnt7[8],pnumcnt6[8]}),
    .e(pnumcnt7[9:8]),
    .mi({open_n37410,\U_AHB/h2h_hwdata [29]}),
    .sr(\U_AHB/n51 ),
    .f({_al_u2258_o,_al_u3103_o}),
    .q({open_n37425,pnum2[29]}));  // src/AHB.v(69)
  // src/AHB.v(67)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2259|U_AHB/reg18_b29  (
    .a({pnumcnt7[10],_al_u3301_o}),
    .b({pnumcnt7[11],\U_AHB/n102 }),
    .c({pnumcnt7[12],\U_AHB/n99 }),
    .clk(clk100m),
    .d({pnumcnt7[13],pnumcnt6[12]}),
    .e({open_n37427,pnumcnt7[12]}),
    .mi({open_n37429,\U_AHB/h2h_hwdata [29]}),
    .sr(\U_AHB/n45 ),
    .f({_al_u2259_o,_al_u3302_o}),
    .q({open_n37444,pnum0[29]}));  // src/AHB.v(67)
  // src/AHB.v(68)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2260|U_AHB/reg19_b24  (
    .a({_al_u2259_o,_al_u3257_o}),
    .b({pnumcnt7[14],\U_AHB/n102 }),
    .c({pnumcnt7[15],\U_AHB/n99 }),
    .clk(clk100m),
    .d({pnumcnt7[16],pnumcnt6[16]}),
    .e(pnumcnt7[17:16]),
    .mi({open_n37447,\U_AHB/h2h_hwdata [24]}),
    .sr(\U_AHB/n47 ),
    .f({_al_u2260_o,_al_u3258_o}),
    .q({open_n37462,pnum1[24]}));  // src/AHB.v(68)
  // src/AHB.v(69)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(~C*~B*~D)"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(~C*~B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000000000000011),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000000000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2261|U_AHB/reg20_b25  (
    .a({open_n37463,_al_u3147_o}),
    .b({pnumcnt7[4],\U_AHB/n102 }),
    .c({pnumcnt7[5],\U_AHB/n99 }),
    .clk(clk100m),
    .d({pnumcnt7[3],pnumcnt6[4]}),
    .e({open_n37465,pnumcnt7[4]}),
    .mi({open_n37467,\U_AHB/h2h_hwdata [25]}),
    .sr(\U_AHB/n51 ),
    .f({_al_u2261_o,_al_u3148_o}),
    .q({open_n37482,pnum2[25]}));  // src/AHB.v(69)
  // src/AHB.v(77)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~(D*C*B*A))"),
    //.LUTF1("(~D*C*B*A)"),
    //.LUTG0("(~1*~(D*C*B*A))"),
    //.LUTG1("(~D*C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111111111111111),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2262|U_AHB/reg28_b26  (
    .a({_al_u2258_o,_al_u2258_o}),
    .b({_al_u2260_o,_al_u2260_o}),
    .c({_al_u2261_o,_al_u2261_o}),
    .clk(clk100m),
    .d({pnumcnt7[0],pnumcnt7[0]}),
    .e({open_n37484,\PWM7/stopreq }),
    .mi({open_n37486,\U_AHB/h2h_hwdata [26]}),
    .sr(\U_AHB/n67 ),
    .f({\PWM7/n25_neg_lutinv ,_al_u3028_o}),
    .q({open_n37501,pnumA[26]}));  // src/AHB.v(77)
  EF2_PHY_PAD #(
    //.LOCATION("P142"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u23 (
    .do({open_n37503,open_n37504,open_n37505,dir_pad[15]}),
    .opad(dir[15]));  // CPLD_SOC_AHB_TOP.v(7)
  // src/OnePWM.v(48)
  EF2_PHY_MSLICE #(
    //.LUT0("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    //.LUT1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100000011001010),
    .INIT_LUT1(16'b1010100000100000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2307|PWM7/reg2_b1  (
    .a({\PWM7/n24 ,\PWM7/pnumr [1]}),
    .b({\PWM7/n25_neg_lutinv ,pnum7[1]}),
    .c({\PWM7/n26 [1],pnum7[32]}),
    .clk(clk100m),
    .d({\PWM7/pnumr [1],pwm_start_stop[23]}),
    .f({_al_u2307_o,open_n37539}),
    .q({open_n37543,\PWM7/pnumr[1]_keep }));  // src/OnePWM.v(48)
  // src/OnePWM.v(58)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~A*~(C*~B))*~(D)*~(0)+~(~A*~(C*~B))*D*~(0)+~(~(~A*~(C*~B)))*D*0+~(~A*~(C*~B))*D*0)"),
    //.LUTF1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    //.LUTG0("(~(~A*~(C*~B))*~(D)*~(1)+~(~A*~(C*~B))*D*~(1)+~(~(~A*~(C*~B)))*D*1+~(~A*~(C*~B))*D*1)"),
    //.LUTG1("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1011101010111010),
    .INIT_LUTF1(16'b1010100000100000),
    .INIT_LUTG0(16'b1111111100000000),
    .INIT_LUTG1(16'b1010100000100000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2309|PWM7/reg3_b0  (
    .a({\PWM7/n24 ,_al_u2309_o}),
    .b({\PWM7/n25_neg_lutinv ,\PWM7/n24 }),
    .c({\PWM7/n26 [0],pnumcnt7[0]}),
    .clk(clk100m),
    .d({\PWM7/pnumr [0],\PWM7/pnumr [0]}),
    .e({open_n37545,pwm_start_stop[23]}),
    .f({_al_u2309_o,open_n37561}),
    .q({open_n37565,\PWM7/RemaTxNum[0]_keep }));  // src/OnePWM.v(58)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*B*D)"),
    .INIT_LUT0(16'b1100000000000000),
    .MODE("LOGIC"))
    _al_u2319 (
    .b({open_n37568,_al_u2316_o}),
    .c({open_n37569,_al_u2318_o}),
    .d({open_n37572,_al_u2314_o}),
    .f({open_n37586,_al_u2319_o}));
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2327|PWM7/reg0_b26  (
    .a({_al_u2321_o,open_n37592}),
    .b({_al_u2323_o,\PWM7/n12 [26]}),
    .c({_al_u2325_o,freq7[26]}),
    .clk(clk100m),
    .d({_al_u2326_o,\PWM7/n0_lutinv }),
    .sr(\PWM7/n11 ),
    .f({_al_u2327_o,open_n37606}),
    .q({open_n37610,\PWM7/FreCnt [26]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0*~C)*~(D@B))"),
    //.LUTF1("(0*D*C*B*A)"),
    //.LUTG0("(A*~(1*~C)*~(D@B))"),
    //.LUTG1("(1*D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000100000100010),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2335|PWM7/reg1_b17  (
    .a({_al_u2319_o,_al_u2329_o}),
    .b({_al_u2327_o,\PWM7/FreCnt [16]}),
    .c({_al_u2330_o,\PWM7/FreCnt [2]}),
    .ce(\PWM7/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({_al_u2332_o,\PWM7/FreCntr [17]}),
    .e({_al_u2334_o,\PWM7/FreCntr [3]}),
    .mi({open_n37612,freq7[17]}),
    .f({_al_u2335_o,_al_u2330_o}),
    .q({open_n37628,\PWM7/FreCntr [17]}));  // src/OnePWM.v(37)
  // src/AHB.v(71)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2338|U_AHB/reg22_b24  (
    .a({pnumcnt8[18],_al_u3236_o}),
    .b({pnumcnt8[19],\U_AHB/n108 }),
    .c({pnumcnt8[1],\U_AHB/n105 }),
    .clk(clk100m),
    .d({pnumcnt8[20],pnumcnt8[18]}),
    .e({open_n37630,pnumcnt9[18]}),
    .mi({open_n37632,\U_AHB/h2h_hwdata [24]}),
    .sr(\U_AHB/n55 ),
    .f({_al_u2338_o,_al_u3237_o}),
    .q({open_n37647,pnum4[24]}));  // src/AHB.v(71)
  // src/AHB.v(70)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2339|U_AHB/reg21_b25  (
    .a({_al_u2338_o,_al_u3181_o}),
    .b({pnumcnt8[21],\U_AHB/n108 }),
    .c({pnumcnt8[22],\U_AHB/n105 }),
    .clk(clk100m),
    .d(pnumcnt8[23:22]),
    .e({pnumcnt8[2],pnumcnt9[22]}),
    .mi({open_n37650,\U_AHB/h2h_hwdata [25]}),
    .sr(\U_AHB/n53 ),
    .f({_al_u2339_o,_al_u3182_o}),
    .q({open_n37665,pnum3[25]}));  // src/AHB.v(70)
  // src/AHB.v(72)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2341|U_AHB/reg23_b31  (
    .a({pnumcnt8[10],_al_u3313_o}),
    .b({pnumcnt8[11],\U_AHB/n108 }),
    .c({pnumcnt8[12],\U_AHB/n105 }),
    .clk(clk100m),
    .d({pnumcnt8[13],pnumcnt8[11]}),
    .e({open_n37667,pnumcnt9[11]}),
    .mi({open_n37669,\U_AHB/h2h_hwdata [31]}),
    .sr(\U_AHB/n57 ),
    .f({_al_u2341_o,_al_u3314_o}),
    .q({open_n37684,pnum5[31]}));  // src/AHB.v(72)
  // src/AHB.v(72)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2342|U_AHB/reg23_b25  (
    .a({_al_u2341_o,_al_u3280_o}),
    .b({pnumcnt8[14],\U_AHB/n108 }),
    .c({pnumcnt8[15],\U_AHB/n105 }),
    .clk(clk100m),
    .d({pnumcnt8[16],pnumcnt8[14]}),
    .e({pnumcnt8[17],pnumcnt9[14]}),
    .mi({open_n37687,\U_AHB/h2h_hwdata [25]}),
    .sr(\U_AHB/n57 ),
    .f({_al_u2342_o,_al_u3281_o}),
    .q({open_n37702,pnum5[25]}));  // src/AHB.v(72)
  // src/AHB.v(74)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(~C*~B*~D)"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(~C*~B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000000000000011),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000000000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2343|U_AHB/reg25_b9  (
    .a({open_n37703,_al_u3159_o}),
    .b({pnumcnt8[4],\U_AHB/n108 }),
    .c({pnumcnt8[5],\U_AHB/n105 }),
    .clk(clk100m),
    .d({pnumcnt8[3],pnumcnt8[3]}),
    .e({open_n37705,pnumcnt9[3]}),
    .mi({open_n37707,\U_AHB/h2h_hwdata [9]}),
    .sr(\U_AHB/n61 ),
    .f({_al_u2343_o,_al_u3160_o}),
    .q({open_n37722,pnum7[9]}));  // src/AHB.v(74)
  // src/AHB.v(75)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(~D*C*B*A)"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(~D*C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2344|U_AHB/reg26_b27  (
    .a({_al_u2340_o,_al_u3346_o}),
    .b({_al_u2342_o,\U_AHB/n108 }),
    .c({_al_u2343_o,\U_AHB/n105 }),
    .clk(clk100m),
    .d({pnumcnt8[0],pnumcnt8[0]}),
    .e({open_n37724,pnumcnt9[0]}),
    .mi({open_n37726,\U_AHB/h2h_hwdata [27]}),
    .sr(\U_AHB/n63 ),
    .f({\PWM8/n25_neg_lutinv ,_al_u3347_o}),
    .q({open_n37741,pnum8[27]}));  // src/AHB.v(75)
  EF2_PHY_PAD #(
    //.LOCATION("P54"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u24 (
    .do({open_n37743,open_n37744,open_n37745,dir_pad[14]}),
    .opad(dir[14]));  // CPLD_SOC_AHB_TOP.v(7)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2407|PWM8/reg0_b2  (
    .a({_al_u2400_o,open_n37765}),
    .b({_al_u2402_o,\PWM8/n12 [2]}),
    .c({_al_u2404_o,freq8[2]}),
    .clk(clk100m),
    .d({_al_u2406_o,\PWM8/n0_lutinv }),
    .sr(\PWM8/n11 ),
    .f({_al_u2407_o,open_n37783}),
    .q({open_n37787,\PWM8/FreCnt [2]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~C*D)"),
    //.LUTF1("(0*D*C*B*A)"),
    //.LUTG0("(~C*D)"),
    //.LUTG1("(1*D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000111100000000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000111100000000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2415|PWM8/reg1_b2  (
    .a({_al_u2398_o,open_n37788}),
    .b({_al_u2407_o,open_n37789}),
    .c({_al_u2410_o,\PWM8/FreCntr [2]}),
    .ce(\PWM8/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({_al_u2412_o,\PWM8/FreCnt [1]}),
    .e({_al_u2414_o,open_n37790}),
    .mi({open_n37792,freq8[2]}),
    .f({_al_u2415_o,_al_u2413_o}),
    .q({open_n37808,\PWM8/FreCntr [2]}));  // src/OnePWM.v(37)
  // src/AHB.v(70)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2418|U_AHB/reg21_b9  (
    .a({pnumcnt9[18],_al_u3225_o}),
    .b({pnumcnt9[19],\U_AHB/n108 }),
    .c({pnumcnt9[1],\U_AHB/n105 }),
    .clk(clk100m),
    .d({pnumcnt9[20],pnumcnt8[19]}),
    .e({open_n37810,pnumcnt9[19]}),
    .mi({open_n37812,\U_AHB/h2h_hwdata [9]}),
    .sr(\U_AHB/n53 ),
    .f({_al_u2418_o,_al_u3226_o}),
    .q({open_n37827,pnum3[9]}));  // src/AHB.v(70)
  // src/AHB.v(69)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2419|U_AHB/reg20_b31  (
    .a({_al_u2418_o,_al_u3170_o}),
    .b({pnumcnt9[21],\U_AHB/n108 }),
    .c({pnumcnt9[22],\U_AHB/n105 }),
    .clk(clk100m),
    .d({pnumcnt9[23],pnumcnt8[23]}),
    .e({pnumcnt9[2],pnumcnt9[23]}),
    .mi({open_n37830,\U_AHB/h2h_hwdata [31]}),
    .sr(\U_AHB/n51 ),
    .f({_al_u2419_o,_al_u3171_o}),
    .q({open_n37845,pnum2[31]}));  // src/AHB.v(69)
  // src/AHB.v(72)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2421|U_AHB/reg23_b30  (
    .a({pnumcnt9[10],_al_u3302_o}),
    .b({pnumcnt9[11],\U_AHB/n108 }),
    .c({pnumcnt9[12],\U_AHB/n105 }),
    .clk(clk100m),
    .d({pnumcnt9[13],pnumcnt8[12]}),
    .e({open_n37847,pnumcnt9[12]}),
    .mi({open_n37849,\U_AHB/h2h_hwdata [30]}),
    .sr(\U_AHB/n57 ),
    .f({_al_u2421_o,_al_u3303_o}),
    .q({open_n37864,pnum5[30]}));  // src/AHB.v(72)
  // src/AHB.v(71)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2422|U_AHB/reg22_b26  (
    .a({_al_u2421_o,_al_u3247_o}),
    .b({pnumcnt9[14],\U_AHB/n108 }),
    .c({pnumcnt9[15],\U_AHB/n105 }),
    .clk(clk100m),
    .d({pnumcnt9[16],pnumcnt8[17]}),
    .e({pnumcnt9[17],pnumcnt9[17]}),
    .mi({open_n37867,\U_AHB/h2h_hwdata [26]}),
    .sr(\U_AHB/n55 ),
    .f({_al_u2422_o,_al_u3248_o}),
    .q({open_n37882,pnum4[26]}));  // src/AHB.v(71)
  // src/AHB.v(74)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(~C*~B*~D)"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(~C*~B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000000000000011),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000000000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2423|U_AHB/reg25_b30  (
    .a({open_n37883,_al_u3148_o}),
    .b({pnumcnt9[4],\U_AHB/n108 }),
    .c({pnumcnt9[5],\U_AHB/n105 }),
    .clk(clk100m),
    .d({pnumcnt9[3],pnumcnt8[4]}),
    .e({open_n37885,pnumcnt9[4]}),
    .mi({open_n37887,\U_AHB/h2h_hwdata [30]}),
    .sr(\U_AHB/n61 ),
    .f({_al_u2423_o,_al_u3149_o}),
    .q({open_n37902,pnum7[30]}));  // src/AHB.v(74)
  // src/AHB.v(82)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(~D*C*B*A)"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(~D*C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2424|U_AHB/reg33_b25  (
    .a({_al_u2420_o,_al_u2419_o}),
    .b({_al_u2422_o,pnumcnt9[6]}),
    .c({_al_u2423_o,pnumcnt9[7]}),
    .clk(clk100m),
    .d({pnumcnt9[0],pnumcnt9[8]}),
    .e({open_n37904,pnumcnt9[9]}),
    .mi({open_n37906,\U_AHB/h2h_hwdata [25]}),
    .sr(\U_AHB/n77 ),
    .f({\PWM9/n25_neg_lutinv ,_al_u2420_o}),
    .q({open_n37921,pnumF[25]}));  // src/AHB.v(82)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~(D*~B)*~(C*~A))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b1000110010101111),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2478|PWM9/reg0_b17  (
    .a({\PWM9/FreCnt [13],open_n37922}),
    .b({\PWM9/FreCnt [17],\PWM9/n12 [17]}),
    .c({\PWM9/FreCntr [14],freq9[17]}),
    .clk(clk100m),
    .d({\PWM9/FreCntr [18],\PWM9/n0_lutinv }),
    .sr(\PWM9/n11 ),
    .f({_al_u2478_o,open_n37936}),
    .q({open_n37940,\PWM9/FreCnt [17]}));  // src/OnePWM.v(37)
  // src/AHB.v(79)
  EF2_PHY_LSLICE #(
    //.LUTF0("~(D*C*B*A)"),
    //.LUTF1("(0*D*C*B*A)"),
    //.LUTG0("~(D*C*B*A)"),
    //.LUTG1("(1*D*C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111111111111111),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0111111111111111),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2488|U_AHB/reg30_b28  (
    .a({_al_u2479_o,_al_u1640_o}),
    .b({_al_u2481_o,_al_u1642_o}),
    .c({_al_u2483_o,_al_u1644_o}),
    .clk(clk100m),
    .d({_al_u2485_o,_al_u1645_o}),
    .e({_al_u2487_o,open_n37942}),
    .mi({open_n37944,\U_AHB/h2h_hwdata [28]}),
    .sr(\U_AHB/n71 ),
    .f({_al_u2488_o,n4_neg}),
    .q({open_n37959,pnumC[28]}));  // src/AHB.v(79)
  // src/AHB.v(74)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~C*~B*~D)"),
    //.LUTF1("(0*D*C*B*A)"),
    //.LUTG0("(~C*~B*~D)"),
    //.LUTG1("(1*D*C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000011),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000000000000011),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2497|U_AHB/reg25_b28  (
    .a({_al_u2488_o,open_n37960}),
    .b({_al_u2490_o,pnumcntA[4]}),
    .c({_al_u2492_o,pnumcntA[5]}),
    .clk(clk100m),
    .d({_al_u2494_o,pnumcntA[3]}),
    .e({_al_u2496_o,open_n37962}),
    .mi({open_n37964,\U_AHB/h2h_hwdata [28]}),
    .sr(\U_AHB/n61 ),
    .f({_al_u2497_o,_al_u2505_o}),
    .q({open_n37979,pnum7[28]}));  // src/AHB.v(74)
  EF2_PHY_PAD #(
    //.LOCATION("P48"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u25 (
    .do({open_n37981,open_n37982,open_n37983,dir_pad[13]}),
    .opad(dir[13]));  // CPLD_SOC_AHB_TOP.v(7)
  // src/AHB.v(53)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*~C)*~(~0*B))"),
    //.LUTF1("(~(~D*B)*~(~C*A))"),
    //.LUTG0("(A*~(D*~C)*~(~1*B))"),
    //.LUTG1("(~(~D*B)*~(~C*A))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010000000100010),
    .INIT_LUTF1(16'b1111010100110001),
    .INIT_LUTG0(16'b1010000010101010),
    .INIT_LUTG1(16'b1111010100110001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2555|U_AHB/reg8_b8  (
    .a({\PWMA/FreCnt [10],_al_u2555_o}),
    .b({\PWMA/FreCnt [15],\PWMA/FreCnt [7]}),
    .c({\PWMA/FreCntr [11],\PWMA/FreCnt [9]}),
    .ce(\U_AHB/n18 ),
    .clk(clk100m),
    .d({\PWMA/FreCntr [16],\PWMA/FreCntr [10]}),
    .e({open_n38003,\PWMA/FreCntr [8]}),
    .mi({open_n38005,\U_AHB/h2h_hwdata [8]}),
    .f({_al_u2555_o,_al_u2556_o}),
    .q({open_n38021,freq7[8]}));  // src/AHB.v(53)
  // src/OnePWM.v(15)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(A*~(~0*C)*~(~D*B))"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(A*~(~1*C)*~(~D*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000101000000010),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1010101000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2563|PWM8/stopreq_reg  (
    .a({_al_u2562_o,open_n38022}),
    .b({\PWMA/FreCnt [12],open_n38023}),
    .c({\PWMA/FreCnt [19],\PWM8/stopreq }),
    .clk(clk100m),
    .d({\PWMA/FreCntr [13],\PWM8/n0_lutinv }),
    .e({\PWMA/FreCntr [20],open_n38025}),
    .sr(pwm_start_stop[8]),
    .f({_al_u2563_o,open_n38040}),
    .q({open_n38044,\PWM8/stopreq_keep }));  // src/OnePWM.v(15)
  // src/AHB.v(76)
  EF2_PHY_MSLICE #(
    //.LUT0("(D*~(C*B*A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0111111100000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2576|U_AHB/reg27_b30  (
    .a({_al_u2570_o,_al_u2561_o}),
    .b({_al_u2572_o,_al_u2568_o}),
    .c({_al_u2574_o,_al_u2576_o}),
    .clk(clk100m),
    .d({_al_u2575_o,pwm_state_read[10]}),
    .mi({open_n38056,\U_AHB/h2h_hwdata [30]}),
    .sr(\U_AHB/n65 ),
    .f({_al_u2576_o,\PWMA/u14_sel_is_1_o }),
    .q({open_n38060,pnum9[30]}));  // src/AHB.v(76)
  // src/AHB.v(82)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2580|U_AHB/reg33_b27  (
    .a({_al_u2579_o,_al_u2580_o}),
    .b({pnumcntB[21],pnumcntB[6]}),
    .c({pnumcntB[22],pnumcntB[7]}),
    .clk(clk100m),
    .d({pnumcntB[23],pnumcntB[8]}),
    .e({pnumcntB[2],pnumcntB[9]}),
    .mi({open_n38063,\U_AHB/h2h_hwdata [27]}),
    .sr(\U_AHB/n77 ),
    .f({_al_u2580_o,_al_u2581_o}),
    .q({open_n38078,pnumF[27]}));  // src/AHB.v(82)
  // src/OnePWM.v(15)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(~D*~C*~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2582|PWM1/stopreq_reg  (
    .a({pnumcntB[10],open_n38079}),
    .b({pnumcntB[11],open_n38080}),
    .c({pnumcntB[12],\PWM1/stopreq }),
    .clk(clk100m),
    .d({pnumcntB[13],\PWM1/n0_lutinv }),
    .sr(pwm_start_stop[1]),
    .f({_al_u2582_o,open_n38094}),
    .q({open_n38098,\PWM1/stopreq_keep }));  // src/OnePWM.v(15)
  // src/AHB.v(84)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~(D*C*B*A))"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(~1*~(D*C*B*A))"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111111111111111),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2583|U_AHB/reg34_b11  (
    .a({_al_u2582_o,_al_u2581_o}),
    .b({pnumcntB[14],_al_u2583_o}),
    .c({pnumcntB[15],_al_u2584_o}),
    .clk(clk100m),
    .d({pnumcntB[16],pnumcntB[0]}),
    .e({pnumcntB[17],\PWMB/stopreq }),
    .mi({open_n38101,\U_AHB/h2h_hwdata [11]}),
    .sr(\U_AHB/n79 ),
    .f({_al_u2583_o,_al_u3040_o}),
    .q({open_n38116,pwm_start_stop[11]}));  // src/AHB.v(84)
  // src/AHB.v(61)
  EF2_PHY_MSLICE #(
    //.LUT0("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    //.LUT1("(~C*~B*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0101001101011111),
    .INIT_LUT1(16'b0000000000000011),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2584|U_AHB/reg15_b2  (
    .a({open_n38117,pnumcntB[5]}),
    .b({pnumcntB[4],pnumcntC[5]}),
    .c({pnumcntB[5],\U_AHB/h2h_haddr [2]}),
    .ce(\U_AHB/n32 ),
    .clk(clk100m),
    .d({pnumcntB[3],\U_AHB/h2h_haddr [3]}),
    .mi({open_n38128,\U_AHB/h2h_hwdata [2]}),
    .f({_al_u2584_o,_al_u3140_o}),
    .q({open_n38133,freqE[2]}));  // src/AHB.v(61)
  EF2_PHY_PAD #(
    //.LOCATION("P45"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u26 (
    .do({open_n38135,open_n38136,open_n38137,dir_pad[12]}),
    .opad(dir[12]));  // CPLD_SOC_AHB_TOP.v(7)
  // src/AHB.v(57)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(B*A*~(~D*C))"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(B*A*~(~D*C))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b1000100000001000),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000100000001000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2637|U_AHB/reg12_b4  (
    .a({_al_u2635_o,_al_u1563_o}),
    .b({_al_u2636_o,\PWMB/FreCnt [11]}),
    .c({\PWMB/FreCnt [10],\PWMB/FreCnt [4]}),
    .ce(\U_AHB/n26 ),
    .clk(clk100m),
    .d({\PWMB/FreCntr [11],\PWMB/FreCntr [11]}),
    .e({open_n38157,\PWMB/FreCntr [4]}),
    .mi({open_n38159,\U_AHB/h2h_hwdata [4]}),
    .f({_al_u2637_o,_al_u1564_o}),
    .q({open_n38175,freqB[4]}));  // src/AHB.v(57)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2650|PWMB/reg1_b22  (
    .a({_al_u2643_o,open_n38176}),
    .b({_al_u2645_o,open_n38177}),
    .c({_al_u2647_o,\PWMB/FreCntr [22]}),
    .ce(\PWMB/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({_al_u2649_o,\PWMB/FreCnt [21]}),
    .mi({open_n38181,freqB[22]}),
    .f({_al_u2650_o,_al_u2651_o}),
    .q({open_n38197,\PWMB/FreCntr [22]}));  // src/OnePWM.v(37)
  // src/AHB.v(76)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(0*D*C*B*A)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(1*D*C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2658|U_AHB/reg27_b29  (
    .a({_al_u2641_o,open_n38198}),
    .b({_al_u2650_o,open_n38199}),
    .c({_al_u2653_o,pwm_state_read[11]}),
    .clk(clk100m),
    .d({_al_u2655_o,_al_u2658_o}),
    .e({_al_u2657_o,open_n38201}),
    .mi({open_n38203,\U_AHB/h2h_hwdata [29]}),
    .sr(\U_AHB/n65 ),
    .f({_al_u2658_o,\PWMB/u14_sel_is_1_o }),
    .q({open_n38218,pnum9[29]}));  // src/AHB.v(76)
  // src/AHB.v(82)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2662|U_AHB/reg33_b28  (
    .a({_al_u2661_o,_al_u2662_o}),
    .b({pnumcntC[21],pnumcntC[6]}),
    .c({pnumcntC[22],pnumcntC[7]}),
    .clk(clk100m),
    .d({pnumcntC[23],pnumcntC[8]}),
    .e({pnumcntC[2],pnumcntC[9]}),
    .mi({open_n38221,\U_AHB/h2h_hwdata [28]}),
    .sr(\U_AHB/n77 ),
    .f({_al_u2662_o,_al_u2663_o}),
    .q({open_n38236,pnumF[28]}));  // src/AHB.v(82)
  // src/OnePWM.v(15)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2664|PWMC/stopreq_reg  (
    .a({pnumcntC[10],open_n38237}),
    .b({pnumcntC[11],open_n38238}),
    .c({pnumcntC[12],\PWMC/stopreq }),
    .clk(clk100m),
    .d({pnumcntC[13],\PWMC/n0_lutinv }),
    .sr(pwm_start_stop[12]),
    .f({_al_u2664_o,open_n38256}),
    .q({open_n38260,\PWMC/stopreq_keep }));  // src/OnePWM.v(15)
  // src/AHB.v(84)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~(D*C*B*A))"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(~1*~(D*C*B*A))"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111111111111111),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2665|U_AHB/reg34_b12  (
    .a({_al_u2664_o,_al_u2663_o}),
    .b({pnumcntC[14],_al_u2665_o}),
    .c({pnumcntC[15],_al_u2666_o}),
    .clk(clk100m),
    .d({pnumcntC[16],pnumcntC[0]}),
    .e({pnumcntC[17],\PWMC/stopreq }),
    .mi({open_n38263,\U_AHB/h2h_hwdata [12]}),
    .sr(\U_AHB/n79 ),
    .f({_al_u2665_o,_al_u3043_o}),
    .q({open_n38278,pwm_start_stop[12]}));  // src/AHB.v(84)
  // src/AHB.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~D*C*B*A)"),
    //.LUTF1("(~C*~B*~D)"),
    //.LUTG0("(~D*C*B*A)"),
    //.LUTG1("(~C*~B*~D)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000010000000),
    .INIT_LUTF1(16'b0000000000000011),
    .INIT_LUTG0(16'b0000000010000000),
    .INIT_LUTG1(16'b0000000000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2666|U_AHB/reg3_b5  (
    .a({open_n38279,_al_u2663_o}),
    .b({pnumcntC[4],_al_u2665_o}),
    .c({pnumcntC[5],_al_u2666_o}),
    .ce(\U_AHB/n8 ),
    .clk(clk100m),
    .d({pnumcntC[3],pnumcntC[0]}),
    .mi({open_n38283,\U_AHB/h2h_hwdata [5]}),
    .f({_al_u2666_o,\PWMC/n25_neg_lutinv }),
    .q({open_n38299,freq2[5]}));  // src/AHB.v(48)
  EF2_PHY_PAD #(
    //.LOCATION("P43"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u27 (
    .do({open_n38301,open_n38302,open_n38303,dir_pad[11]}),
    .opad(dir[11]));  // CPLD_SOC_AHB_TOP.v(7)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(D@B)*~(C@A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000010000100001),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2731|PWMC/reg1_b19  (
    .a({_al_u2725_o,\PWMC/FreCnt [18]}),
    .b({_al_u2727_o,\PWMC/FreCnt [2]}),
    .c({_al_u2729_o,\PWMC/FreCntr [19]}),
    .ce(\PWMC/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({_al_u2730_o,\PWMC/FreCntr [3]}),
    .mi({open_n38333,freqC[19]}),
    .f({_al_u2731_o,_al_u2726_o}),
    .q({open_n38338,\PWMC/FreCntr [19]}));  // src/OnePWM.v(37)
  // src/AHB.v(62)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2740|U_AHB/reg16_b5  (
    .a({pnumcntD[18],_al_u3238_o}),
    .b({pnumcntD[19],\U_AHB/n90 }),
    .c({pnumcntD[1],\U_AHB/n87 }),
    .ce(\U_AHB/n34 ),
    .clk(clk100m),
    .d({pnumcntD[20],pnumcntD[18]}),
    .e({open_n38339,pnumcntE[18]}),
    .mi({open_n38341,\U_AHB/h2h_hwdata [5]}),
    .f({_al_u2740_o,_al_u3239_o}),
    .q({open_n38357,freqF[5]}));  // src/AHB.v(62)
  // src/AHB.v(76)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~(D*C*B*A))"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(~1*~(D*C*B*A))"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111111111111111),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2742|U_AHB/reg27_b26  (
    .a({_al_u2741_o,_al_u2742_o}),
    .b({pnumcntD[6],_al_u2744_o}),
    .c({pnumcntD[7],_al_u2745_o}),
    .clk(clk100m),
    .d({pnumcntD[8],pnumcntD[0]}),
    .e({pnumcntD[9],\PWMD/stopreq }),
    .mi({open_n38360,\U_AHB/h2h_hwdata [26]}),
    .sr(\U_AHB/n65 ),
    .f({_al_u2742_o,_al_u3046_o}),
    .q({open_n38375,pnum9[26]}));  // src/AHB.v(76)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2743|_al_u2744  (
    .a({pnumcntD[10],_al_u2743_o}),
    .b({pnumcntD[11],pnumcntD[14]}),
    .c({pnumcntD[12],pnumcntD[15]}),
    .d({pnumcntD[13],pnumcntD[16]}),
    .e({open_n38378,pnumcntD[17]}),
    .f({_al_u2743_o,_al_u2744_o}));
  // src/OnePWM.v(15)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(~C*~B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000000000000011),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2745|PWMD/stopreq_reg  (
    .b({pnumcntD[4],open_n38401}),
    .c({pnumcntD[5],\PWMD/stopreq }),
    .clk(clk100m),
    .d({pnumcntD[3],\PWMD/n0_lutinv }),
    .sr(pwm_start_stop[13]),
    .f({_al_u2745_o,open_n38415}),
    .q({open_n38419,\PWMD/stopreq_keep }));  // src/OnePWM.v(15)
  // src/AHB.v(49)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(~D*C*B*A)"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(~D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2746|U_AHB/reg4_b24  (
    .a({_al_u2742_o,_al_u3349_o}),
    .b({_al_u2744_o,\U_AHB/n90 }),
    .c({_al_u2745_o,\U_AHB/n87 }),
    .ce(\U_AHB/n10 ),
    .clk(clk100m),
    .d({pnumcntD[0],pnumcntD[0]}),
    .e({open_n38420,pnumcntE[0]}),
    .mi({open_n38422,\U_AHB/h2h_hwdata [24]}),
    .f({\PWMD/n25_neg_lutinv ,_al_u3350_o}),
    .q({open_n38438,freq3[24]}));  // src/AHB.v(49)
  EF2_PHY_SPAD #(
    //.LOCATION("P106"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("16"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u28 (
    .do({open_n38441,dir_pad[10]}),
    .ts(1'b1),
    .opad(dir[10]));  // CPLD_SOC_AHB_TOP.v(7)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(D*~(C@B))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1100001100000000),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2808|PWMD/reg1_b25  (
    .a({_al_u2802_o,open_n38448}),
    .b({_al_u2804_o,\PWMD/FreCnt [24]}),
    .c({_al_u2806_o,\PWMD/FreCntr [25]}),
    .ce(\PWMD/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({_al_u2807_o,_al_u2801_o}),
    .mi({open_n38459,freqD[25]}),
    .f({_al_u2808_o,_al_u2802_o}),
    .q({open_n38464,\PWMD/FreCntr [25]}));  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(0*D*C*B*A)"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(1*D*C*B*A)"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b0000000000000000),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2817|_al_u1594  (
    .a({_al_u2800_o,_al_u1593_o}),
    .b({_al_u2808_o,\PWMD/FreCnt [13]}),
    .c({_al_u2812_o,\PWMD/FreCnt [19]}),
    .d({_al_u2814_o,\PWMD/FreCntr [13]}),
    .e({_al_u2816_o,\PWMD/FreCntr [19]}),
    .f({_al_u2817_o,_al_u1594_o}));
  // src/OnePWM.v(15)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(~D*~C*~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2820|PWM6/stopreq_reg  (
    .a({pnumcntE[18],open_n38487}),
    .b({pnumcntE[19],open_n38488}),
    .c({pnumcntE[1],\PWM6/stopreq }),
    .clk(clk100m),
    .d({pnumcntE[20],\PWM6/n0_lutinv }),
    .sr(pwm_start_stop[6]),
    .f({_al_u2820_o,open_n38502}),
    .q({open_n38506,\PWM6/stopreq_keep }));  // src/OnePWM.v(15)
  // src/AHB.v(70)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~D*~C*~B*~A)"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(~D*~C*~B*~A)"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000001),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b0000000000000001),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2821|U_AHB/reg21_b30  (
    .a({_al_u2820_o,pnumcntA[18]}),
    .b({pnumcntE[21],pnumcntA[19]}),
    .c({pnumcntE[22],pnumcntA[1]}),
    .clk(clk100m),
    .d({pnumcntE[23],pnumcntA[20]}),
    .e({pnumcntE[2],open_n38508}),
    .mi({open_n38510,\U_AHB/h2h_hwdata [30]}),
    .sr(\U_AHB/n53 ),
    .f({_al_u2821_o,_al_u2500_o}),
    .q({open_n38525,pnum3[30]}));  // src/AHB.v(70)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"))
    \_al_u2823|_al_u2824  (
    .a({pnumcntE[10],_al_u2823_o}),
    .b({pnumcntE[11],pnumcntE[14]}),
    .c({pnumcntE[12],pnumcntE[15]}),
    .d({pnumcntE[13],pnumcntE[16]}),
    .e({open_n38528,pnumcntE[17]}),
    .f({_al_u2823_o,_al_u2824_o}));
  // src/OnePWM.v(15)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(~C*~B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000000000000011),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \_al_u2825|PWME/stopreq_reg  (
    .b({pnumcntE[4],open_n38551}),
    .c({pnumcntE[5],\PWME/stopreq }),
    .clk(clk100m),
    .d({pnumcntE[3],\PWME/n0_lutinv }),
    .sr(pwm_start_stop[14]),
    .f({_al_u2825_o,open_n38565}),
    .q({open_n38569,\PWME/stopreq_keep }));  // src/OnePWM.v(15)
  // src/AHB.v(75)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~(D*C*B*A))"),
    //.LUTF1("(~D*C*B*A)"),
    //.LUTG0("(~1*~(D*C*B*A))"),
    //.LUTG1("(~D*C*B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0111111111111111),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2826|U_AHB/reg26_b9  (
    .a({_al_u2822_o,_al_u2822_o}),
    .b({_al_u2824_o,_al_u2824_o}),
    .c({_al_u2825_o,_al_u2825_o}),
    .clk(clk100m),
    .d({pnumcntE[0],pnumcntE[0]}),
    .e({open_n38571,\PWME/stopreq }),
    .mi({open_n38573,\U_AHB/h2h_hwdata [9]}),
    .sr(\U_AHB/n63 ),
    .f({\PWME/n25_neg_lutinv ,_al_u3049_o}),
    .q({open_n38588,pnum8[9]}));  // src/AHB.v(75)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2881|PWME/reg0_b17  (
    .b({open_n38591,\PWME/n12 [17]}),
    .c({\PWME/FreCntr [18],freqE[17]}),
    .clk(clk100m),
    .d({\PWME/FreCnt [17],\PWME/n0_lutinv }),
    .sr(\PWME/n11 ),
    .f({_al_u2881_o,open_n38605}),
    .q({open_n38609,\PWME/FreCnt [17]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(C@B)*~(D@A))"),
    //.LUT1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000001001000001),
    .INIT_LUT1(16'b1000000000000000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2896|PWME/reg1_b21  (
    .a({_al_u2890_o,\PWME/FreCnt [2]}),
    .b({_al_u2892_o,\PWME/FreCnt [20]}),
    .c({_al_u2894_o,\PWME/FreCntr [21]}),
    .ce(\PWME/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({_al_u2895_o,\PWME/FreCntr [3]}),
    .mi({open_n38620,freqE[21]}),
    .f({_al_u2896_o,_al_u2891_o}),
    .q({open_n38625,\PWME/FreCntr [21]}));  // src/OnePWM.v(37)
  // src/AHB.v(62)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2899|U_AHB/reg16_b9  (
    .a({pnumcntF[18],_al_u3339_o}),
    .b({pnumcntF[19],\U_AHB/n96 }),
    .c({pnumcntF[1],\U_AHB/n93 }),
    .ce(\U_AHB/n34 ),
    .clk(clk100m),
    .d({pnumcntF[20],pnumcntF[1]}),
    .e({open_n38626,pwm_state_read[1]}),
    .mi({open_n38628,\U_AHB/h2h_hwdata [9]}),
    .f({_al_u2899_o,_al_u3340_o}),
    .q({open_n38644,freqF[9]}));  // src/AHB.v(62)
  EF2_PHY_PAD #(
    //.LOCATION("P42"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u29 (
    .do({open_n38646,open_n38647,open_n38648,dir_pad[9]}),
    .opad(dir[9]));  // CPLD_SOC_AHB_TOP.v(7)
  // src/AHB.v(70)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2900|U_AHB/reg21_b24  (
    .a({_al_u2899_o,_al_u3185_o}),
    .b({pnumcntF[21],\U_AHB/n96 }),
    .c({pnumcntF[22],\U_AHB/n93 }),
    .clk(clk100m),
    .d(pnumcntF[23:22]),
    .e({pnumcntF[2],pwm_state_read[6]}),
    .mi({open_n38670,\U_AHB/h2h_hwdata [24]}),
    .sr(\U_AHB/n53 ),
    .f({_al_u2900_o,_al_u3186_o}),
    .q({open_n38685,pnum3[24]}));  // src/AHB.v(70)
  // src/AHB.v(72)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2902|U_AHB/reg23_b26  (
    .a({pnumcntF[10],_al_u3295_o}),
    .b({pnumcntF[11],\U_AHB/n96 }),
    .c({pnumcntF[12],\U_AHB/n93 }),
    .clk(clk100m),
    .d({pnumcntF[13],pnumcntF[13]}),
    .e({open_n38687,pwm_state_read[13]}),
    .mi({open_n38689,\U_AHB/h2h_hwdata [26]}),
    .sr(\U_AHB/n57 ),
    .f({_al_u2902_o,_al_u3296_o}),
    .q({open_n38704,pnum5[26]}));  // src/AHB.v(72)
  // src/AHB.v(71)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2903|U_AHB/reg22_b9  (
    .a({_al_u2902_o,_al_u3284_o}),
    .b({pnumcntF[14],\U_AHB/n96 }),
    .c({pnumcntF[15],\U_AHB/n93 }),
    .clk(clk100m),
    .d({pnumcntF[16],pnumcntF[14]}),
    .e({pnumcntF[17],pwm_state_read[14]}),
    .mi({open_n38707,\U_AHB/h2h_hwdata [9]}),
    .sr(\U_AHB/n55 ),
    .f({_al_u2903_o,_al_u3285_o}),
    .q({open_n38722,pnum4[9]}));  // src/AHB.v(71)
  // src/AHB.v(74)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(~C*~B*~D)"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(~C*~B*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000000000000011),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000000000000011),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u2904|U_AHB/reg25_b31  (
    .a({open_n38723,_al_u3163_o}),
    .b({pnumcntF[4],\U_AHB/n96 }),
    .c({pnumcntF[5],\U_AHB/n93 }),
    .clk(clk100m),
    .d({pnumcntF[3],pnumcntF[3]}),
    .e({open_n38725,pwm_state_read[3]}),
    .mi({open_n38727,\U_AHB/h2h_hwdata [31]}),
    .sr(\U_AHB/n61 ),
    .f({_al_u2904_o,_al_u3164_o}),
    .q({open_n38742,pnum7[31]}));  // src/AHB.v(74)
  // src/AHB.v(62)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(~D*C*B*A)"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(~D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000000010000000),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000000010000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2905|U_AHB/reg16_b6  (
    .a({_al_u2901_o,_al_u3350_o}),
    .b({_al_u2903_o,\U_AHB/n96 }),
    .c({_al_u2904_o,\U_AHB/n93 }),
    .ce(\U_AHB/n34 ),
    .clk(clk100m),
    .d({pnumcntF[0],pnumcntF[0]}),
    .e({open_n38743,pwm_state_read[0]}),
    .mi({open_n38745,\U_AHB/h2h_hwdata [6]}),
    .f({\PWMF/n25_neg_lutinv ,_al_u3351_o}),
    .q({open_n38761,freqF[6]}));  // src/AHB.v(62)
  // src/AHB.v(62)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~D*B*A*~(~0*C))"),
    //.LUTF1("(D*C*B*A)"),
    //.LUTG0("(~D*B*A*~(~1*C))"),
    //.LUTG1("(D*C*B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000001000),
    .INIT_LUTF1(16'b1000000000000000),
    .INIT_LUTG0(16'b0000000010001000),
    .INIT_LUTG1(16'b1000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u2963|U_AHB/reg16_b11  (
    .a({_al_u2956_o,_al_u2954_o}),
    .b({_al_u2958_o,_al_u2955_o}),
    .c({_al_u2960_o,\PWMF/FreCnt [10]}),
    .ce(\U_AHB/n34 ),
    .clk(clk100m),
    .d({_al_u2962_o,\PWMF/FreCnt [26]}),
    .e({open_n38762,\PWMF/FreCntr [11]}),
    .mi({open_n38764,\U_AHB/h2h_hwdata [11]}),
    .f({_al_u2963_o,_al_u2956_o}),
    .q({open_n38780,freqF[11]}));  // src/AHB.v(62)
  EF2_PHY_PAD #(
    //.LOCATION("P114"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u30 (
    .do({open_n38782,open_n38783,open_n38784,dir_pad[8]}),
    .opad(dir[8]));  // CPLD_SOC_AHB_TOP.v(7)
  // src/AHB.v(52)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3085|U_AHB/reg7_b26  (
    .a({_al_u3082_o,_al_u3085_o}),
    .b({\U_AHB/n90 ,\U_AHB/n96 }),
    .c({\U_AHB/n87 ,\U_AHB/n93 }),
    .ce(\U_AHB/n16 ),
    .clk(clk100m),
    .d({pnumcnt2[9],pnumcnt4[9]}),
    .e({pnumcnt3[9],pnumcnt5[9]}),
    .mi({open_n38805,\U_AHB/h2h_hwdata [26]}),
    .f({_al_u3085_o,_al_u3087_o}),
    .q({open_n38821,freq6[26]}));  // src/AHB.v(52)
  EF2_PHY_PAD #(
    //.LOCATION("P122"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u31 (
    .do({open_n38823,open_n38824,open_n38825,dir_pad[7]}),
    .opad(dir[7]));  // CPLD_SOC_AHB_TOP.v(7)
  // src/AHB.v(52)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3101|U_AHB/reg7_b24  (
    .a({_al_u3100_o,_al_u3101_o}),
    .b({\U_AHB/n90 ,\U_AHB/n96 }),
    .c({\U_AHB/n87 ,\U_AHB/n93 }),
    .ce(\U_AHB/n16 ),
    .clk(clk100m),
    .d({pnumcnt2[8],pnumcnt4[8]}),
    .e({pnumcnt3[8],pnumcnt5[8]}),
    .mi({open_n38846,\U_AHB/h2h_hwdata [24]}),
    .f({_al_u3101_o,_al_u3102_o}),
    .q({open_n38862,freq6[24]}));  // src/AHB.v(52)
  // src/AHB.v(61)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~((0*C)*~(B)*~(D)+(0*C)*B*~(D)+~((0*C))*B*D+(0*C)*B*D))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~((1*C)*~(B)*~(D)+(1*C)*B*~(D)+~((1*C))*B*D+(1*C)*B*D))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0010001000001010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3107|U_AHB/reg15_b25  (
    .a({_al_u3106_o,_al_u3061_o}),
    .b({\U_AHB/n90 ,pnumcntB[8]}),
    .c({\U_AHB/n87 ,pnumcntC[8]}),
    .ce(\U_AHB/n32 ),
    .clk(clk100m),
    .d({pnumcntD[8],\U_AHB/h2h_haddr [2]}),
    .e({pnumcntE[8],\U_AHB/h2h_haddr [3]}),
    .mi({open_n38864,\U_AHB/h2h_hwdata [25]}),
    .f({_al_u3107_o,_al_u3106_o}),
    .q({open_n38880,freqE[25]}));  // src/AHB.v(61)
  // src/AHB.v(51)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3112|U_AHB/reg6_b9  (
    .a({_al_u3111_o,_al_u3112_o}),
    .b({\U_AHB/n90 ,\U_AHB/n96 }),
    .c({\U_AHB/n87 ,\U_AHB/n93 }),
    .ce(\U_AHB/n14 ),
    .clk(clk100m),
    .d({pnumcnt2[7],pnumcnt4[7]}),
    .e({pnumcnt3[7],pnumcnt5[7]}),
    .mi({open_n38882,\U_AHB/h2h_hwdata [9]}),
    .f({_al_u3112_o,_al_u3113_o}),
    .q({open_n38898,freq5[9]}));  // src/AHB.v(51)
  // src/AHB.v(61)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~((0*C)*~(B)*~(D)+(0*C)*B*~(D)+~((0*C))*B*D+(0*C)*B*D))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~((1*C)*~(B)*~(D)+(1*C)*B*~(D)+~((1*C))*B*D+(1*C)*B*D))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0010001000001010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3118|U_AHB/reg15_b23  (
    .a({_al_u3117_o,_al_u3061_o}),
    .b({\U_AHB/n90 ,pnumcntB[7]}),
    .c({\U_AHB/n87 ,pnumcntC[7]}),
    .ce(\U_AHB/n32 ),
    .clk(clk100m),
    .d({pnumcntD[7],\U_AHB/h2h_haddr [2]}),
    .e({pnumcntE[7],\U_AHB/h2h_haddr [3]}),
    .mi({open_n38900,\U_AHB/h2h_hwdata [23]}),
    .f({_al_u3118_o,_al_u3117_o}),
    .q({open_n38916,freqE[23]}));  // src/AHB.v(61)
  // src/AHB.v(51)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3123|U_AHB/reg6_b8  (
    .a({_al_u3122_o,_al_u3123_o}),
    .b({\U_AHB/n90 ,\U_AHB/n96 }),
    .c({\U_AHB/n87 ,\U_AHB/n93 }),
    .ce(\U_AHB/n14 ),
    .clk(clk100m),
    .d({pnumcnt2[6],pnumcnt4[6]}),
    .e({pnumcnt3[6],pnumcnt5[6]}),
    .mi({open_n38918,\U_AHB/h2h_hwdata [8]}),
    .f({_al_u3123_o,_al_u3124_o}),
    .q({open_n38934,freq5[8]}));  // src/AHB.v(51)
  // src/AHB.v(61)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~((0*C)*~(B)*~(D)+(0*C)*B*~(D)+~((0*C))*B*D+(0*C)*B*D))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~((1*C)*~(B)*~(D)+(1*C)*B*~(D)+~((1*C))*B*D+(1*C)*B*D))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0010001000001010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3129|U_AHB/reg15_b21  (
    .a({_al_u3128_o,_al_u3061_o}),
    .b({\U_AHB/n90 ,pnumcntB[6]}),
    .c({\U_AHB/n87 ,pnumcntC[6]}),
    .ce(\U_AHB/n32 ),
    .clk(clk100m),
    .d({pnumcntD[6],\U_AHB/h2h_haddr [2]}),
    .e({pnumcntE[6],\U_AHB/h2h_haddr [3]}),
    .mi({open_n38936,\U_AHB/h2h_hwdata [21]}),
    .f({_al_u3129_o,_al_u3128_o}),
    .q({open_n38952,freqE[21]}));  // src/AHB.v(61)
  // src/AHB.v(51)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3134|U_AHB/reg6_b5  (
    .a({_al_u3133_o,_al_u3134_o}),
    .b({\U_AHB/n90 ,\U_AHB/n96 }),
    .c({\U_AHB/n87 ,\U_AHB/n93 }),
    .ce(\U_AHB/n14 ),
    .clk(clk100m),
    .d({pnumcnt2[5],pnumcnt4[5]}),
    .e({pnumcnt3[5],pnumcnt5[5]}),
    .mi({open_n38954,\U_AHB/h2h_hwdata [5]}),
    .f({_al_u3134_o,_al_u3135_o}),
    .q({open_n38970,freq5[5]}));  // src/AHB.v(51)
  // src/AHB.v(74)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*A*~(D*C))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(B*A*~(D*C))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100010001000),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000100010001000),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u3141|U_AHB/reg25_b26  (
    .a({_al_u3140_o,_al_u3139_o}),
    .b({\U_AHB/n90 ,_al_u3141_o}),
    .c({\U_AHB/n87 ,\U_AHB/n93 }),
    .clk(clk100m),
    .d({pnumcntD[5],pnumcntF[5]}),
    .e({pnumcntE[5],open_n38972}),
    .mi({open_n38974,\U_AHB/h2h_hwdata [26]}),
    .sr(\U_AHB/n61 ),
    .f({_al_u3141_o,_al_u3142_o}),
    .q({open_n38989,pnum7[26]}));  // src/AHB.v(74)
  // src/AHB.v(51)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3146|U_AHB/reg6_b26  (
    .a({_al_u3145_o,_al_u3146_o}),
    .b({\U_AHB/n90 ,\U_AHB/n96 }),
    .c({\U_AHB/n87 ,\U_AHB/n93 }),
    .ce(\U_AHB/n14 ),
    .clk(clk100m),
    .d({pnumcnt2[4],pnumcnt4[4]}),
    .e({pnumcnt3[4],pnumcnt5[4]}),
    .mi({open_n38991,\U_AHB/h2h_hwdata [26]}),
    .f({_al_u3146_o,_al_u3147_o}),
    .q({open_n39007,freq5[26]}));  // src/AHB.v(51)
  // src/AHB.v(61)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~((0*C)*~(B)*~(D)+(0*C)*B*~(D)+~((0*C))*B*D+(0*C)*B*D))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~((1*C)*~(B)*~(D)+(1*C)*B*~(D)+~((1*C))*B*D+(1*C)*B*D))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0010001000001010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3152|U_AHB/reg15_b18  (
    .a({_al_u3151_o,_al_u3061_o}),
    .b({\U_AHB/n90 ,pnumcntB[4]}),
    .c({\U_AHB/n87 ,pnumcntC[4]}),
    .ce(\U_AHB/n32 ),
    .clk(clk100m),
    .d({pnumcntD[4],\U_AHB/h2h_haddr [2]}),
    .e({pnumcntE[4],\U_AHB/h2h_haddr [3]}),
    .mi({open_n39009,\U_AHB/h2h_hwdata [18]}),
    .f({_al_u3152_o,_al_u3151_o}),
    .q({open_n39025,freqE[18]}));  // src/AHB.v(61)
  // src/AHB.v(51)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3157|U_AHB/reg6_b25  (
    .a({_al_u3156_o,_al_u3157_o}),
    .b({\U_AHB/n90 ,\U_AHB/n96 }),
    .c({\U_AHB/n87 ,\U_AHB/n93 }),
    .ce(\U_AHB/n14 ),
    .clk(clk100m),
    .d({pnumcnt2[3],pnumcnt4[3]}),
    .e({pnumcnt3[3],pnumcnt5[3]}),
    .mi({open_n39027,\U_AHB/h2h_hwdata [25]}),
    .f({_al_u3157_o,_al_u3158_o}),
    .q({open_n39043,freq5[25]}));  // src/AHB.v(51)
  // src/AHB.v(61)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~((0*C)*~(B)*~(D)+(0*C)*B*~(D)+~((0*C))*B*D+(0*C)*B*D))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~((1*C)*~(B)*~(D)+(1*C)*B*~(D)+~((1*C))*B*D+(1*C)*B*D))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0010001000001010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3163|U_AHB/reg15_b16  (
    .a({_al_u3162_o,_al_u3061_o}),
    .b({\U_AHB/n90 ,pnumcntB[3]}),
    .c({\U_AHB/n87 ,pnumcntC[3]}),
    .ce(\U_AHB/n32 ),
    .clk(clk100m),
    .d({pnumcntD[3],\U_AHB/h2h_haddr [2]}),
    .e({pnumcntE[3],\U_AHB/h2h_haddr [3]}),
    .mi({open_n39045,\U_AHB/h2h_hwdata [16]}),
    .f({_al_u3163_o,_al_u3162_o}),
    .q({open_n39061,freqE[16]}));  // src/AHB.v(61)
  // src/AHB.v(51)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3168|U_AHB/reg6_b19  (
    .a({_al_u3167_o,_al_u3168_o}),
    .b({\U_AHB/n90 ,\U_AHB/n96 }),
    .c({\U_AHB/n87 ,\U_AHB/n93 }),
    .ce(\U_AHB/n14 ),
    .clk(clk100m),
    .d({pnumcnt2[23],pnumcnt4[23]}),
    .e({pnumcnt3[23],pnumcnt5[23]}),
    .mi({open_n39063,\U_AHB/h2h_hwdata [19]}),
    .f({_al_u3168_o,_al_u3169_o}),
    .q({open_n39079,freq5[19]}));  // src/AHB.v(51)
  // src/AHB.v(61)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~((0*C)*~(B)*~(D)+(0*C)*B*~(D)+~((0*C))*B*D+(0*C)*B*D))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~((1*C)*~(B)*~(D)+(1*C)*B*~(D)+~((1*C))*B*D+(1*C)*B*D))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0010001000001010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3174|U_AHB/reg15_b14  (
    .a({_al_u3173_o,_al_u3061_o}),
    .b({\U_AHB/n90 ,pnumcntB[23]}),
    .c({\U_AHB/n87 ,pnumcntC[23]}),
    .ce(\U_AHB/n32 ),
    .clk(clk100m),
    .d({pnumcntD[23],\U_AHB/h2h_haddr [2]}),
    .e({pnumcntE[23],\U_AHB/h2h_haddr [3]}),
    .mi({open_n39081,\U_AHB/h2h_hwdata [14]}),
    .f({_al_u3174_o,_al_u3173_o}),
    .q({open_n39097,freqE[14]}));  // src/AHB.v(61)
  // src/AHB.v(50)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3179|U_AHB/reg5_b9  (
    .a({_al_u3178_o,_al_u3179_o}),
    .b({\U_AHB/n90 ,\U_AHB/n96 }),
    .c({\U_AHB/n87 ,\U_AHB/n93 }),
    .ce(\U_AHB/n12 ),
    .clk(clk100m),
    .d({pnumcnt2[22],pnumcnt4[22]}),
    .e({pnumcnt3[22],pnumcnt5[22]}),
    .mi({open_n39099,\U_AHB/h2h_hwdata [9]}),
    .f({_al_u3179_o,_al_u3180_o}),
    .q({open_n39115,freq4[9]}));  // src/AHB.v(50)
  // src/AHB.v(61)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~((0*C)*~(B)*~(D)+(0*C)*B*~(D)+~((0*C))*B*D+(0*C)*B*D))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~((1*C)*~(B)*~(D)+(1*C)*B*~(D)+~((1*C))*B*D+(1*C)*B*D))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0010001000001010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3185|U_AHB/reg15_b12  (
    .a({_al_u3184_o,_al_u3061_o}),
    .b({\U_AHB/n90 ,pnumcntB[22]}),
    .c({\U_AHB/n87 ,pnumcntC[22]}),
    .ce(\U_AHB/n32 ),
    .clk(clk100m),
    .d({pnumcntD[22],\U_AHB/h2h_haddr [2]}),
    .e({pnumcntE[22],\U_AHB/h2h_haddr [3]}),
    .mi({open_n39117,\U_AHB/h2h_hwdata [12]}),
    .f({_al_u3185_o,_al_u3184_o}),
    .q({open_n39133,freqE[12]}));  // src/AHB.v(61)
  // src/AHB.v(50)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3190|U_AHB/reg5_b5  (
    .a({_al_u3189_o,_al_u3190_o}),
    .b({\U_AHB/n90 ,\U_AHB/n96 }),
    .c({\U_AHB/n87 ,\U_AHB/n93 }),
    .ce(\U_AHB/n12 ),
    .clk(clk100m),
    .d({pnumcnt2[21],pnumcnt4[21]}),
    .e({pnumcnt3[21],pnumcnt5[21]}),
    .mi({open_n39135,\U_AHB/h2h_hwdata [5]}),
    .f({_al_u3190_o,_al_u3191_o}),
    .q({open_n39151,freq4[5]}));  // src/AHB.v(50)
  // src/AHB.v(70)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*A*~(D*C))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(B*A*~(D*C))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100010001000),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000100010001000),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u3196|U_AHB/reg21_b26  (
    .a({_al_u3195_o,_al_u3139_o}),
    .b({\U_AHB/n90 ,_al_u3196_o}),
    .c({\U_AHB/n87 ,\U_AHB/n93 }),
    .clk(clk100m),
    .d({pnumcntD[21],pnumcntF[21]}),
    .e({pnumcntE[21],open_n39153}),
    .mi({open_n39155,\U_AHB/h2h_hwdata [26]}),
    .sr(\U_AHB/n53 ),
    .f({_al_u3196_o,_al_u3197_o}),
    .q({open_n39170,pnum3[26]}));  // src/AHB.v(70)
  EF2_PHY_SPAD #(
    //.LOCATION("P24"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("16"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u32 (
    .do({open_n39173,dir_pad[6]}),
    .ts(1'b1),
    .opad(dir[6]));  // CPLD_SOC_AHB_TOP.v(7)
  // src/AHB.v(50)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3201|U_AHB/reg5_b4  (
    .a({_al_u3200_o,_al_u3201_o}),
    .b({\U_AHB/n90 ,\U_AHB/n96 }),
    .c({\U_AHB/n87 ,\U_AHB/n93 }),
    .ce(\U_AHB/n12 ),
    .clk(clk100m),
    .d({pnumcnt2[20],pnumcnt4[20]}),
    .e({pnumcnt3[20],pnumcnt5[20]}),
    .mi({open_n39181,\U_AHB/h2h_hwdata [4]}),
    .f({_al_u3201_o,_al_u3202_o}),
    .q({open_n39197,freq4[4]}));  // src/AHB.v(50)
  // src/AHB.v(60)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~((0*C)*~(B)*~(D)+(0*C)*B*~(D)+~((0*C))*B*D+(0*C)*B*D))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~((1*C)*~(B)*~(D)+(1*C)*B*~(D)+~((1*C))*B*D+(1*C)*B*D))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0010001000001010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3207|U_AHB/reg14_b9  (
    .a({_al_u3206_o,_al_u3061_o}),
    .b({\U_AHB/n90 ,pnumcntB[20]}),
    .c({\U_AHB/n87 ,pnumcntC[20]}),
    .ce(\U_AHB/n30 ),
    .clk(clk100m),
    .d({pnumcntD[20],\U_AHB/h2h_haddr [2]}),
    .e({pnumcntE[20],\U_AHB/h2h_haddr [3]}),
    .mi({open_n39199,\U_AHB/h2h_hwdata [9]}),
    .f({_al_u3207_o,_al_u3206_o}),
    .q({open_n39215,freqD[9]}));  // src/AHB.v(60)
  // src/AHB.v(50)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3212|U_AHB/reg5_b26  (
    .a({_al_u3211_o,_al_u3212_o}),
    .b({\U_AHB/n90 ,\U_AHB/n96 }),
    .c({\U_AHB/n87 ,\U_AHB/n93 }),
    .ce(\U_AHB/n12 ),
    .clk(clk100m),
    .d({pnumcnt2[2],pnumcnt4[2]}),
    .e({pnumcnt3[2],pnumcnt5[2]}),
    .mi({open_n39217,\U_AHB/h2h_hwdata [26]}),
    .f({_al_u3212_o,_al_u3213_o}),
    .q({open_n39233,freq4[26]}));  // src/AHB.v(50)
  // src/AHB.v(60)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~((0*C)*~(B)*~(D)+(0*C)*B*~(D)+~((0*C))*B*D+(0*C)*B*D))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~((1*C)*~(B)*~(D)+(1*C)*B*~(D)+~((1*C))*B*D+(1*C)*B*D))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0010001000001010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3218|U_AHB/reg14_b7  (
    .a({_al_u3217_o,_al_u3061_o}),
    .b({\U_AHB/n90 ,pnumcntB[2]}),
    .c({\U_AHB/n87 ,pnumcntC[2]}),
    .ce(\U_AHB/n30 ),
    .clk(clk100m),
    .d({pnumcntD[2],\U_AHB/h2h_haddr [2]}),
    .e({pnumcntE[2],\U_AHB/h2h_haddr [3]}),
    .mi({open_n39235,\U_AHB/h2h_hwdata [7]}),
    .f({_al_u3218_o,_al_u3217_o}),
    .q({open_n39251,freqD[7]}));  // src/AHB.v(60)
  // src/AHB.v(50)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3223|U_AHB/reg5_b25  (
    .a({_al_u3222_o,_al_u3223_o}),
    .b({\U_AHB/n90 ,\U_AHB/n96 }),
    .c({\U_AHB/n87 ,\U_AHB/n93 }),
    .ce(\U_AHB/n12 ),
    .clk(clk100m),
    .d({pnumcnt2[19],pnumcnt4[19]}),
    .e({pnumcnt3[19],pnumcnt5[19]}),
    .mi({open_n39253,\U_AHB/h2h_hwdata [25]}),
    .f({_al_u3223_o,_al_u3224_o}),
    .q({open_n39269,freq4[25]}));  // src/AHB.v(50)
  // src/AHB.v(60)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~((0*C)*~(B)*~(D)+(0*C)*B*~(D)+~((0*C))*B*D+(0*C)*B*D))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~((1*C)*~(B)*~(D)+(1*C)*B*~(D)+~((1*C))*B*D+(1*C)*B*D))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0010001000001010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3229|U_AHB/reg14_b5  (
    .a({_al_u3228_o,_al_u3061_o}),
    .b({\U_AHB/n90 ,pnumcntB[19]}),
    .c({\U_AHB/n87 ,pnumcntC[19]}),
    .ce(\U_AHB/n30 ),
    .clk(clk100m),
    .d({pnumcntD[19],\U_AHB/h2h_haddr [2]}),
    .e({pnumcntE[19],\U_AHB/h2h_haddr [3]}),
    .mi({open_n39271,\U_AHB/h2h_hwdata [5]}),
    .f({_al_u3229_o,_al_u3228_o}),
    .q({open_n39287,freqD[5]}));  // src/AHB.v(60)
  // src/AHB.v(60)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~((0*C)*~(B)*~(D)+(0*C)*B*~(D)+~((0*C))*B*D+(0*C)*B*D))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~((1*C)*~(B)*~(D)+(1*C)*B*~(D)+~((1*C))*B*D+(1*C)*B*D))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0010001000001010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3234|U_AHB/reg14_b4  (
    .a({_al_u3233_o,\U_AHB/n82 }),
    .b({\U_AHB/n90 ,pnumcnt0[18]}),
    .c({\U_AHB/n87 ,pnumcnt1[18]}),
    .ce(\U_AHB/n30 ),
    .clk(clk100m),
    .d({pnumcnt2[18],\U_AHB/h2h_haddr [2]}),
    .e({pnumcnt3[18],\U_AHB/h2h_haddr [3]}),
    .mi({open_n39289,\U_AHB/h2h_hwdata [4]}),
    .f({_al_u3234_o,_al_u3233_o}),
    .q({open_n39305,freqD[4]}));  // src/AHB.v(60)
  // src/AHB.v(47)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3245|U_AHB/reg2_b9  (
    .a({_al_u3244_o,_al_u3245_o}),
    .b({\U_AHB/n90 ,\U_AHB/n96 }),
    .c({\U_AHB/n87 ,\U_AHB/n93 }),
    .ce(\U_AHB/n4 ),
    .clk(clk100m),
    .d({pnumcnt2[17],pnumcnt4[17]}),
    .e({pnumcnt3[17],pnumcnt5[17]}),
    .mi({open_n39307,\U_AHB/h2h_hwdata [9]}),
    .f({_al_u3245_o,_al_u3246_o}),
    .q({open_n39323,freq1[9]}));  // src/AHB.v(47)
  // src/AHB.v(60)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~((0*C)*~(B)*~(D)+(0*C)*B*~(D)+~((0*C))*B*D+(0*C)*B*D))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~((1*C)*~(B)*~(D)+(1*C)*B*~(D)+~((1*C))*B*D+(1*C)*B*D))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0010001000001010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3251|U_AHB/reg14_b26  (
    .a({_al_u3250_o,_al_u3061_o}),
    .b({\U_AHB/n90 ,pnumcntB[17]}),
    .c({\U_AHB/n87 ,pnumcntC[17]}),
    .ce(\U_AHB/n30 ),
    .clk(clk100m),
    .d({pnumcntD[17],\U_AHB/h2h_haddr [2]}),
    .e({pnumcntE[17],\U_AHB/h2h_haddr [3]}),
    .mi({open_n39325,\U_AHB/h2h_hwdata [26]}),
    .f({_al_u3251_o,_al_u3250_o}),
    .q({open_n39341,freqD[26]}));  // src/AHB.v(60)
  // src/AHB.v(47)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3256|U_AHB/reg2_b8  (
    .a({_al_u3255_o,_al_u3256_o}),
    .b({\U_AHB/n90 ,\U_AHB/n96 }),
    .c({\U_AHB/n87 ,\U_AHB/n93 }),
    .ce(\U_AHB/n4 ),
    .clk(clk100m),
    .d({pnumcnt2[16],pnumcnt4[16]}),
    .e({pnumcnt3[16],pnumcnt5[16]}),
    .mi({open_n39343,\U_AHB/h2h_hwdata [8]}),
    .f({_al_u3256_o,_al_u3257_o}),
    .q({open_n39359,freq1[8]}));  // src/AHB.v(47)
  // src/AHB.v(60)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~((0*C)*~(B)*~(D)+(0*C)*B*~(D)+~((0*C))*B*D+(0*C)*B*D))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~((1*C)*~(B)*~(D)+(1*C)*B*~(D)+~((1*C))*B*D+(1*C)*B*D))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0010001000001010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3262|U_AHB/reg14_b24  (
    .a({_al_u3261_o,_al_u3061_o}),
    .b({\U_AHB/n90 ,pnumcntB[16]}),
    .c({\U_AHB/n87 ,pnumcntC[16]}),
    .ce(\U_AHB/n30 ),
    .clk(clk100m),
    .d({pnumcntD[16],\U_AHB/h2h_haddr [2]}),
    .e({pnumcntE[16],\U_AHB/h2h_haddr [3]}),
    .mi({open_n39361,\U_AHB/h2h_hwdata [24]}),
    .f({_al_u3262_o,_al_u3261_o}),
    .q({open_n39377,freqD[24]}));  // src/AHB.v(60)
  // src/AHB.v(47)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3267|U_AHB/reg2_b5  (
    .a({_al_u3266_o,_al_u3267_o}),
    .b({\U_AHB/n90 ,\U_AHB/n96 }),
    .c({\U_AHB/n87 ,\U_AHB/n93 }),
    .ce(\U_AHB/n4 ),
    .clk(clk100m),
    .d({pnumcnt2[15],pnumcnt4[15]}),
    .e({pnumcnt3[15],pnumcnt5[15]}),
    .mi({open_n39379,\U_AHB/h2h_hwdata [5]}),
    .f({_al_u3267_o,_al_u3268_o}),
    .q({open_n39395,freq1[5]}));  // src/AHB.v(47)
  // src/AHB.v(60)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~((0*C)*~(B)*~(D)+(0*C)*B*~(D)+~((0*C))*B*D+(0*C)*B*D))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~((1*C)*~(B)*~(D)+(1*C)*B*~(D)+~((1*C))*B*D+(1*C)*B*D))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0010001000001010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3273|U_AHB/reg14_b22  (
    .a({_al_u3272_o,_al_u3061_o}),
    .b({\U_AHB/n90 ,pnumcntB[15]}),
    .c({\U_AHB/n87 ,pnumcntC[15]}),
    .ce(\U_AHB/n30 ),
    .clk(clk100m),
    .d({pnumcntD[15],\U_AHB/h2h_haddr [2]}),
    .e({pnumcntE[15],\U_AHB/h2h_haddr [3]}),
    .mi({open_n39397,\U_AHB/h2h_hwdata [22]}),
    .f({_al_u3273_o,_al_u3272_o}),
    .q({open_n39413,freqD[22]}));  // src/AHB.v(60)
  // src/AHB.v(47)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3278|U_AHB/reg2_b4  (
    .a({_al_u3277_o,_al_u3278_o}),
    .b({\U_AHB/n90 ,\U_AHB/n96 }),
    .c({\U_AHB/n87 ,\U_AHB/n93 }),
    .ce(\U_AHB/n4 ),
    .clk(clk100m),
    .d({pnumcnt2[14],pnumcnt4[14]}),
    .e({pnumcnt3[14],pnumcnt5[14]}),
    .mi({open_n39415,\U_AHB/h2h_hwdata [4]}),
    .f({_al_u3278_o,_al_u3279_o}),
    .q({open_n39431,freq1[4]}));  // src/AHB.v(47)
  // src/AHB.v(60)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~((0*C)*~(B)*~(D)+(0*C)*B*~(D)+~((0*C))*B*D+(0*C)*B*D))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~((1*C)*~(B)*~(D)+(1*C)*B*~(D)+~((1*C))*B*D+(1*C)*B*D))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0010001000001010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3284|U_AHB/reg14_b20  (
    .a({_al_u3283_o,_al_u3061_o}),
    .b({\U_AHB/n90 ,pnumcntB[14]}),
    .c({\U_AHB/n87 ,pnumcntC[14]}),
    .ce(\U_AHB/n30 ),
    .clk(clk100m),
    .d({pnumcntD[14],\U_AHB/h2h_haddr [2]}),
    .e({pnumcntE[14],\U_AHB/h2h_haddr [3]}),
    .mi({open_n39433,\U_AHB/h2h_hwdata [20]}),
    .f({_al_u3284_o,_al_u3283_o}),
    .q({open_n39449,freqD[20]}));  // src/AHB.v(60)
  // src/AHB.v(47)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3289|U_AHB/reg2_b26  (
    .a({_al_u3288_o,_al_u3289_o}),
    .b({\U_AHB/n90 ,\U_AHB/n96 }),
    .c({\U_AHB/n87 ,\U_AHB/n93 }),
    .ce(\U_AHB/n4 ),
    .clk(clk100m),
    .d({pnumcnt2[13],pnumcnt4[13]}),
    .e({pnumcnt3[13],pnumcnt5[13]}),
    .mi({open_n39451,\U_AHB/h2h_hwdata [26]}),
    .f({_al_u3289_o,_al_u3290_o}),
    .q({open_n39467,freq1[26]}));  // src/AHB.v(47)
  // src/AHB.v(60)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~((0*C)*~(B)*~(D)+(0*C)*B*~(D)+~((0*C))*B*D+(0*C)*B*D))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~((1*C)*~(B)*~(D)+(1*C)*B*~(D)+~((1*C))*B*D+(1*C)*B*D))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0010001000001010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3295|U_AHB/reg14_b19  (
    .a({_al_u3294_o,_al_u3061_o}),
    .b({\U_AHB/n90 ,pnumcntB[13]}),
    .c({\U_AHB/n87 ,pnumcntC[13]}),
    .ce(\U_AHB/n30 ),
    .clk(clk100m),
    .d({pnumcntD[13],\U_AHB/h2h_haddr [2]}),
    .e({pnumcntE[13],\U_AHB/h2h_haddr [3]}),
    .mi({open_n39469,\U_AHB/h2h_hwdata [19]}),
    .f({_al_u3295_o,_al_u3294_o}),
    .q({open_n39485,freqD[19]}));  // src/AHB.v(60)
  EF2_PHY_SPAD #(
    //.LOCATION("P23"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("16"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u33 (
    .do({open_n39488,dir_pad[5]}),
    .ts(1'b1),
    .opad(dir[5]));  // CPLD_SOC_AHB_TOP.v(7)
  // src/AHB.v(47)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3300|U_AHB/reg2_b25  (
    .a({_al_u3299_o,_al_u3300_o}),
    .b({\U_AHB/n90 ,\U_AHB/n96 }),
    .c({\U_AHB/n87 ,\U_AHB/n93 }),
    .ce(\U_AHB/n4 ),
    .clk(clk100m),
    .d({pnumcnt2[12],pnumcnt4[12]}),
    .e({pnumcnt3[12],pnumcnt5[12]}),
    .mi({open_n39496,\U_AHB/h2h_hwdata [25]}),
    .f({_al_u3300_o,_al_u3301_o}),
    .q({open_n39512,freq1[25]}));  // src/AHB.v(47)
  // src/AHB.v(60)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~((0*C)*~(B)*~(D)+(0*C)*B*~(D)+~((0*C))*B*D+(0*C)*B*D))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~((1*C)*~(B)*~(D)+(1*C)*B*~(D)+~((1*C))*B*D+(1*C)*B*D))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0010001000001010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3306|U_AHB/reg14_b17  (
    .a({_al_u3305_o,_al_u3061_o}),
    .b({\U_AHB/n90 ,pnumcntB[12]}),
    .c({\U_AHB/n87 ,pnumcntC[12]}),
    .ce(\U_AHB/n30 ),
    .clk(clk100m),
    .d({pnumcntD[12],\U_AHB/h2h_haddr [2]}),
    .e({pnumcntE[12],\U_AHB/h2h_haddr [3]}),
    .mi({open_n39514,\U_AHB/h2h_hwdata [17]}),
    .f({_al_u3306_o,_al_u3305_o}),
    .q({open_n39530,freqD[17]}));  // src/AHB.v(60)
  // src/AHB.v(46)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3311|U_AHB/reg1_b8  (
    .a({_al_u3310_o,_al_u3311_o}),
    .b({\U_AHB/n90 ,\U_AHB/n96 }),
    .c({\U_AHB/n87 ,\U_AHB/n93 }),
    .ce(\U_AHB/n2 ),
    .clk(clk100m),
    .d({pnumcnt2[11],pnumcnt4[11]}),
    .e({pnumcnt3[11],pnumcnt5[11]}),
    .mi({open_n39532,\U_AHB/h2h_hwdata [8]}),
    .f({_al_u3311_o,_al_u3312_o}),
    .q({open_n39548,freq0[8]}));  // src/AHB.v(46)
  // src/AHB.v(60)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~((0*C)*~(B)*~(D)+(0*C)*B*~(D)+~((0*C))*B*D+(0*C)*B*D))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~((1*C)*~(B)*~(D)+(1*C)*B*~(D)+~((1*C))*B*D+(1*C)*B*D))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0010001000001010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3317|U_AHB/reg14_b15  (
    .a({_al_u3316_o,_al_u3061_o}),
    .b({\U_AHB/n90 ,pnumcntB[11]}),
    .c({\U_AHB/n87 ,pnumcntC[11]}),
    .ce(\U_AHB/n30 ),
    .clk(clk100m),
    .d({pnumcntD[11],\U_AHB/h2h_haddr [2]}),
    .e({pnumcntE[11],\U_AHB/h2h_haddr [3]}),
    .mi({open_n39550,\U_AHB/h2h_hwdata [15]}),
    .f({_al_u3317_o,_al_u3316_o}),
    .q({open_n39566,freqD[15]}));  // src/AHB.v(60)
  // src/AHB.v(46)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3322|U_AHB/reg1_b26  (
    .a({_al_u3321_o,_al_u3322_o}),
    .b({\U_AHB/n90 ,\U_AHB/n96 }),
    .c({\U_AHB/n87 ,\U_AHB/n93 }),
    .ce(\U_AHB/n2 ),
    .clk(clk100m),
    .d({pnumcnt2[10],pnumcnt4[10]}),
    .e({pnumcnt3[10],pnumcnt5[10]}),
    .mi({open_n39568,\U_AHB/h2h_hwdata [26]}),
    .f({_al_u3322_o,_al_u3323_o}),
    .q({open_n39584,freq0[26]}));  // src/AHB.v(46)
  // src/AHB.v(60)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~((0*C)*~(B)*~(D)+(0*C)*B*~(D)+~((0*C))*B*D+(0*C)*B*D))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~((1*C)*~(B)*~(D)+(1*C)*B*~(D)+~((1*C))*B*D+(1*C)*B*D))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0010001000001010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3328|U_AHB/reg14_b13  (
    .a({_al_u3327_o,_al_u3061_o}),
    .b({\U_AHB/n90 ,pnumcntB[10]}),
    .c({\U_AHB/n87 ,pnumcntC[10]}),
    .ce(\U_AHB/n30 ),
    .clk(clk100m),
    .d({pnumcntD[10],\U_AHB/h2h_haddr [2]}),
    .e({pnumcntE[10],\U_AHB/h2h_haddr [3]}),
    .mi({open_n39586,\U_AHB/h2h_hwdata [13]}),
    .f({_al_u3328_o,_al_u3327_o}),
    .q({open_n39602,freqD[13]}));  // src/AHB.v(60)
  EF2_PHY_MSLICE #(
    //.LUT0("(A*~(D*C)*~(0*B))"),
    //.LUT1("(A*~(D*C)*~(1*B))"),
    .INIT_LUT0(16'b0000101010101010),
    .INIT_LUT1(16'b0000001000100010),
    .MODE("LOGIC"),
    .MSFXMUX("ON"))
    _al_u3333 (
    .a({_al_u3332_o,_al_u3332_o}),
    .b({\U_AHB/n90 ,\U_AHB/n90 }),
    .c({\U_AHB/n87 ,\U_AHB/n87 }),
    .d({pnumcnt2[1],pnumcnt2[1]}),
    .mi({open_n39615,pnumcnt3[1]}),
    .fx({open_n39620,_al_u3333_o}));
  // src/AHB.v(60)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~((0*C)*~(B)*~(D)+(0*C)*B*~(D)+~((0*C))*B*D+(0*C)*B*D))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~((1*C)*~(B)*~(D)+(1*C)*B*~(D)+~((1*C))*B*D+(1*C)*B*D))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0010001010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0010001000001010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3339|U_AHB/reg14_b11  (
    .a({_al_u3338_o,_al_u3061_o}),
    .b({\U_AHB/n90 ,pnumcntB[1]}),
    .c({\U_AHB/n87 ,pnumcntC[1]}),
    .ce(\U_AHB/n30 ),
    .clk(clk100m),
    .d({pnumcntD[1],\U_AHB/h2h_haddr [2]}),
    .e({pnumcntE[1],\U_AHB/h2h_haddr [3]}),
    .mi({open_n39624,\U_AHB/h2h_hwdata [11]}),
    .f({_al_u3339_o,_al_u3338_o}),
    .q({open_n39640,freqD[11]}));  // src/AHB.v(60)
  // src/AHB.v(62)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(D*C)*~(0*B))"),
    //.LUTF1("(A*~(D*C)*~(0*B))"),
    //.LUTG0("(A*~(D*C)*~(1*B))"),
    //.LUTG1("(A*~(D*C)*~(1*B))"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000101010101010),
    .INIT_LUTF1(16'b0000101010101010),
    .INIT_LUTG0(16'b0000001000100010),
    .INIT_LUTG1(16'b0000001000100010),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u3344|U_AHB/reg16_b8  (
    .a({_al_u3343_o,_al_u3344_o}),
    .b({\U_AHB/n90 ,\U_AHB/n96 }),
    .c({\U_AHB/n87 ,\U_AHB/n93 }),
    .ce(\U_AHB/n34 ),
    .clk(clk100m),
    .d({pnumcnt2[0],pnumcnt4[0]}),
    .e({pnumcnt3[0],pnumcnt5[0]}),
    .mi({open_n39642,\U_AHB/h2h_hwdata [8]}),
    .f({_al_u3344_o,_al_u3345_o}),
    .q({open_n39658,freqF[8]}));  // src/AHB.v(62)
  EF2_PHY_SPAD #(
    //.LOCATION("P22"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("16"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u34 (
    .do({open_n39661,dir_pad[4]}),
    .ts(1'b1),
    .opad(dir[4]));  // CPLD_SOC_AHB_TOP.v(7)
  EF2_PHY_PAD #(
    //.LOCATION("P132"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u35 (
    .do({open_n39669,open_n39670,open_n39671,dir_pad[3]}),
    .opad(dir[3]));  // CPLD_SOC_AHB_TOP.v(7)
  EF2_PHY_PAD #(
    //.LOCATION("P133"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u36 (
    .do({open_n39692,open_n39693,open_n39694,dir_pad[2]}),
    .opad(dir[2]));  // CPLD_SOC_AHB_TOP.v(7)
  EF2_PHY_SPAD #(
    //.LOCATION("P21"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("16"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u37 (
    .do({open_n39716,dir_pad[1]}),
    .ts(1'b1),
    .opad(dir[1]));  // CPLD_SOC_AHB_TOP.v(7)
  EF2_PHY_PAD #(
    //.LOCATION("P138"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u38 (
    .do({open_n39724,open_n39725,open_n39726,dir_pad[0]}),
    .opad(dir[0]));  // CPLD_SOC_AHB_TOP.v(7)
  EF2_PHY_SPAD #(
    //.LOCATION("p10"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u39 (
    .do({open_n39748,gpio_out_pad[31]}),
    .ts(1'b1),
    .opad(gpio_out[31]));  // CPLD_SOC_AHB_TOP.v(8)
  EF2_PHY_PAD #(
    //.LOCATION("p120"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u40 (
    .do({open_n39756,open_n39757,open_n39758,gpio_out_pad[30]}),
    .opad(gpio_out[30]));  // CPLD_SOC_AHB_TOP.v(8)
  EF2_PHY_SPAD #(
    //.LOCATION("p19"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u41 (
    .do({open_n39780,gpio_out_pad[29]}),
    .ts(1'b1),
    .opad(gpio_out[29]));  // CPLD_SOC_AHB_TOP.v(8)
  EF2_PHY_PAD #(
    //.LOCATION("p61"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u42 (
    .do({open_n39788,open_n39789,open_n39790,gpio_out_pad[28]}),
    .opad(gpio_out[28]));  // CPLD_SOC_AHB_TOP.v(8)
  EF2_PHY_PAD #(
    //.LOCATION("p62"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u43 (
    .do({open_n39811,open_n39812,open_n39813,gpio_out_pad[27]}),
    .opad(gpio_out[27]));  // CPLD_SOC_AHB_TOP.v(8)
  EF2_PHY_SPAD #(
    //.LOCATION("p91"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u44 (
    .do({open_n39835,gpio_out_pad[26]}),
    .ts(1'b1),
    .opad(gpio_out[26]));  // CPLD_SOC_AHB_TOP.v(8)
  EF2_PHY_PAD #(
    //.LOCATION("p109"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u45 (
    .do({open_n39843,open_n39844,open_n39845,gpio_out_pad[25]}),
    .opad(gpio_out[25]));  // CPLD_SOC_AHB_TOP.v(8)
  EF2_PHY_PAD #(
    //.LOCATION("p143"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u46 (
    .do({open_n39866,open_n39867,open_n39868,gpio_out_pad[24]}),
    .opad(gpio_out[24]));  // CPLD_SOC_AHB_TOP.v(8)
  EF2_PHY_PAD #(
    //.LOCATION("p71"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u47 (
    .do({open_n39889,open_n39890,open_n39891,gpio_out_pad[23]}),
    .opad(gpio_out[23]));  // CPLD_SOC_AHB_TOP.v(8)
  EF2_PHY_SPAD #(
    //.LOCATION("p73"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u48 (
    .do({open_n39913,gpio_out_pad[22]}),
    .ts(1'b1),
    .opad(gpio_out[22]));  // CPLD_SOC_AHB_TOP.v(8)
  EF2_PHY_SPAD #(
    //.LOCATION("p11"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u49 (
    .do({open_n39922,gpio_out_pad[21]}),
    .ts(1'b1),
    .opad(gpio_out[21]));  // CPLD_SOC_AHB_TOP.v(8)
  EF2_PHY_SPAD #(
    //.LOCATION("p13"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u50 (
    .do({open_n39931,gpio_out_pad[20]}),
    .ts(1'b1),
    .opad(gpio_out[20]));  // CPLD_SOC_AHB_TOP.v(8)
  EF2_PHY_PAD #(
    //.LOCATION("p39"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u51 (
    .do({open_n39939,open_n39940,open_n39941,gpio_out_pad[19]}),
    .opad(gpio_out[19]));  // CPLD_SOC_AHB_TOP.v(8)
  EF2_PHY_SPAD #(
    //.LOCATION("p74"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u52 (
    .do({open_n39963,gpio_out_pad[18]}),
    .ts(1'b1),
    .opad(gpio_out[18]));  // CPLD_SOC_AHB_TOP.v(8)
  EF2_PHY_PAD #(
    //.LOCATION("p110"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u53 (
    .do({open_n39971,open_n39972,open_n39973,gpio_out_pad[17]}),
    .opad(gpio_out[17]));  // CPLD_SOC_AHB_TOP.v(8)
  EF2_PHY_PAD #(
    //.LOCATION("p140"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u54 (
    .do({open_n39994,open_n39995,open_n39996,gpio_out_pad[16]}),
    .opad(gpio_out[16]));  // CPLD_SOC_AHB_TOP.v(8)
  EF2_PHY_SPAD #(
    //.LOCATION("p75"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u55 (
    .do({open_n40018,gpio_out_pad[15]}),
    .ts(1'b1),
    .opad(gpio_out[15]));  // CPLD_SOC_AHB_TOP.v(8)
  EF2_PHY_SPAD #(
    //.LOCATION("p9"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u56 (
    .do({open_n40027,gpio_out_pad[14]}),
    .ts(1'b1),
    .opad(gpio_out[14]));  // CPLD_SOC_AHB_TOP.v(8)
  EF2_PHY_PAD #(
    //.LOCATION("p139"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u57 (
    .do({open_n40035,open_n40036,open_n40037,gpio_out_pad[13]}),
    .opad(gpio_out[13]));  // CPLD_SOC_AHB_TOP.v(8)
  EF2_PHY_SPAD #(
    //.LOCATION("p76"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u58 (
    .do({open_n40059,gpio_out_pad[12]}),
    .ts(1'b1),
    .opad(gpio_out[12]));  // CPLD_SOC_AHB_TOP.v(8)
  EF2_PHY_SPAD #(
    //.LOCATION("p83"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u59 (
    .do({open_n40068,gpio_out_pad[11]}),
    .ts(1'b1),
    .opad(gpio_out[11]));  // CPLD_SOC_AHB_TOP.v(8)
  EF2_PHY_SPAD #(
    //.LOCATION("p12"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u60 (
    .do({open_n40077,gpio_out_pad[10]}),
    .ts(1'b1),
    .opad(gpio_out[10]));  // CPLD_SOC_AHB_TOP.v(8)
  EF2_PHY_SPAD #(
    //.LOCATION("p77"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u61 (
    .do({open_n40086,gpio_out_pad[9]}),
    .ts(1'b1),
    .opad(gpio_out[9]));  // CPLD_SOC_AHB_TOP.v(8)
  EF2_PHY_SPAD #(
    //.LOCATION("p84"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u62 (
    .do({open_n40095,gpio_out_pad[8]}),
    .ts(1'b1),
    .opad(gpio_out[8]));  // CPLD_SOC_AHB_TOP.v(8)
  EF2_PHY_SPAD #(
    //.LOCATION("p14"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u63 (
    .do({open_n40104,gpio_out_pad[7]}),
    .ts(1'b1),
    .opad(gpio_out[7]));  // CPLD_SOC_AHB_TOP.v(8)
  EF2_PHY_SPAD #(
    //.LOCATION("p78"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u64 (
    .do({open_n40113,gpio_out_pad[6]}),
    .ts(1'b1),
    .opad(gpio_out[6]));  // CPLD_SOC_AHB_TOP.v(8)
  EF2_PHY_SPAD #(
    //.LOCATION("p97"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u65 (
    .do({open_n40122,gpio_out_pad[5]}),
    .ts(1'b1),
    .opad(gpio_out[5]));  // CPLD_SOC_AHB_TOP.v(8)
  EF2_PHY_SPAD #(
    //.LOCATION("p15"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u66 (
    .do({open_n40131,gpio_out_pad[4]}),
    .ts(1'b1),
    .opad(gpio_out[4]));  // CPLD_SOC_AHB_TOP.v(8)
  EF2_PHY_SPAD #(
    //.LOCATION("p92"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u67 (
    .do({open_n40140,gpio_out_pad[3]}),
    .ts(1'b1),
    .opad(gpio_out[3]));  // CPLD_SOC_AHB_TOP.v(8)
  EF2_PHY_SPAD #(
    //.LOCATION("p17"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u68 (
    .do({open_n40149,gpio_out_pad[2]}),
    .ts(1'b1),
    .opad(gpio_out[2]));  // CPLD_SOC_AHB_TOP.v(8)
  EF2_PHY_SPAD #(
    //.LOCATION("p93"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u69 (
    .do({open_n40158,gpio_out_pad[1]}),
    .ts(1'b1),
    .opad(gpio_out[1]));  // CPLD_SOC_AHB_TOP.v(8)
  EF2_PHY_SPAD #(
    //.LOCATION("p98"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u70 (
    .do({open_n40167,gpio_out_pad[0]}),
    .ts(1'b1),
    .opad(gpio_out[0]));  // CPLD_SOC_AHB_TOP.v(8)
  EF2_PHY_SPAD #(
    //.LOCATION("P100"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("16"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u71 (
    .do({open_n40176,ledout_pad[3]}),
    .ts(1'b1),
    .opad(ledout[3]));  // CPLD_SOC_AHB_TOP.v(10)
  EF2_PHY_SPAD #(
    //.LOCATION("P103"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("16"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u72 (
    .do({open_n40185,ledout_pad[2]}),
    .ts(1'b1),
    .opad(ledout[2]));  // CPLD_SOC_AHB_TOP.v(10)
  EF2_PHY_SPAD #(
    //.LOCATION("P104"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("16"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u73 (
    .do({open_n40194,ledout_pad[1]}),
    .ts(1'b1),
    .opad(ledout[1]));  // CPLD_SOC_AHB_TOP.v(10)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u737|PWM0/reg0_b2  (
    .a({\PWM0/FreCnt [0],open_n40201}),
    .b({\PWM0/FreCnt [1],\PWM0/n12 [2]}),
    .c({\PWM0/FreCnt [10],freq0[2]}),
    .clk(clk100m),
    .d({\PWM0/FreCnt [11],\PWM0/n0_lutinv }),
    .sr(\PWM0/n11 ),
    .f({_al_u737_o,open_n40219}),
    .q({open_n40223,\PWM0/FreCnt [2]}));  // src/OnePWM.v(37)
  // src/AHB.v(46)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u738|U_AHB/reg1_b20  (
    .a({_al_u737_o,_al_u1373_o}),
    .b({\PWM0/FreCnt [12],\PWM0/FreCnt [14]}),
    .c({\PWM0/FreCnt [13],\PWM0/FreCnt [20]}),
    .ce(\U_AHB/n2 ),
    .clk(clk100m),
    .d({\PWM0/FreCnt [14],\PWM0/FreCntr [14]}),
    .e({\PWM0/FreCnt [15],\PWM0/FreCntr [20]}),
    .mi({open_n40225,\U_AHB/h2h_hwdata [20]}),
    .f({_al_u738_o,_al_u1374_o}),
    .q({open_n40241,freq0[20]}));  // src/AHB.v(46)
  // src/OnePWM.v(37)
  EF2_PHY_MSLICE #(
    //.LUT0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUT1("(~D*~C*~B*~A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111000011001100),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u739|PWM0/reg0_b19  (
    .a({\PWM0/FreCnt [16],open_n40242}),
    .b({\PWM0/FreCnt [17],\PWM0/n12 [19]}),
    .c({\PWM0/FreCnt [18],freq0[19]}),
    .clk(clk100m),
    .d({\PWM0/FreCnt [19],\PWM0/n0_lutinv }),
    .sr(\PWM0/n11 ),
    .f({_al_u739_o,open_n40256}),
    .q({open_n40260,\PWM0/FreCnt [19]}));  // src/OnePWM.v(37)
  EF2_PHY_SPAD #(
    //.LOCATION("P87"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u74 (
    .ipad(limit_l[15]),
    .ts(1'b1),
    .di(limit_l_pad[15]));  // CPLD_SOC_AHB_TOP.v(5)
  EF2_PHY_SPAD #(
    //.LOCATION("P85"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u75 (
    .ipad(limit_l[14]),
    .ts(1'b1),
    .di(limit_l_pad[14]));  // CPLD_SOC_AHB_TOP.v(5)
  EF2_PHY_SPAD #(
    //.LOCATION("P1"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u76 (
    .ipad(limit_l[13]),
    .ts(1'b1),
    .di(limit_l_pad[13]));  // CPLD_SOC_AHB_TOP.v(5)
  EF2_PHY_PAD #(
    //.LOCATION("P69"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u77 (
    .ipad(limit_l[12]),
    .di(limit_l_pad[12]));  // CPLD_SOC_AHB_TOP.v(5)
  // src/AHB.v(47)
  EF2_PHY_MSLICE #(
    //.LUT0("(~(D@B)*~(C@A))"),
    //.LUT1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1000010000100001),
    .INIT_LUT1(16'b0000000000000001),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u774|U_AHB/reg2_b22  (
    .a({\PWM1/FreCnt [0],\PWM1/FreCnt [22]}),
    .b({\PWM1/FreCnt [1],\PWM1/FreCnt [23]}),
    .c({\PWM1/FreCnt [10],\PWM1/FreCntr [22]}),
    .ce(\U_AHB/n4 ),
    .clk(clk100m),
    .d({\PWM1/FreCnt [11],\PWM1/FreCntr [23]}),
    .mi({open_n40321,\U_AHB/h2h_hwdata [22]}),
    .f({_al_u774_o,_al_u1378_o}),
    .q({open_n40326,freq1[22]}));  // src/AHB.v(47)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u775|PWM1/reg0_b15  (
    .a({_al_u774_o,open_n40327}),
    .b({\PWM1/FreCnt [12],\PWM1/n12 [15]}),
    .c({\PWM1/FreCnt [13],freq1[15]}),
    .clk(clk100m),
    .d({\PWM1/FreCnt [14],\PWM1/n0_lutinv }),
    .e({\PWM1/FreCnt [15],open_n40329}),
    .sr(\PWM1/n11 ),
    .f({_al_u775_o,open_n40344}),
    .q({open_n40348,\PWM1/FreCnt [15]}));  // src/OnePWM.v(37)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(D*~B)*~(C*~A))"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(~(D*~B)*~(C*~A))"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1000110010101111),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b1000110010101111),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u777|PWM1/reg1_b13  (
    .a({_al_u776_o,\PWM1/FreCnt [12]}),
    .b({\PWM1/FreCnt [2],\PWM1/FreCnt [21]}),
    .c({\PWM1/FreCnt [20],\PWM1/FreCntr [13]}),
    .ce(\PWM1/mux3_b0_sel_is_3_o ),
    .clk(clk100m),
    .d({\PWM1/FreCnt [21],\PWM1/FreCntr [22]}),
    .e({\PWM1/FreCnt [22],open_n40349}),
    .mi({open_n40351,freq1[13]}),
    .f({_al_u777_o,_al_u1826_o}),
    .q({open_n40367,\PWM1/FreCntr [13]}));  // src/OnePWM.v(37)
  EF2_PHY_PAD #(
    //.LOCATION("P67"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u78 (
    .ipad(limit_l[11]),
    .di(limit_l_pad[11]));  // CPLD_SOC_AHB_TOP.v(5)
  EF2_PHY_PAD #(
    //.LOCATION("P65"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u79 (
    .ipad(limit_l[10]),
    .di(limit_l_pad[10]));  // CPLD_SOC_AHB_TOP.v(5)
  EF2_PHY_SPAD #(
    //.LOCATION("P34"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u80 (
    .ipad(limit_l[9]),
    .ts(1'b1),
    .di(limit_l_pad[9]));  // CPLD_SOC_AHB_TOP.v(5)
  EF2_PHY_SPAD #(
    //.LOCATION("P33"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u81 (
    .ipad(limit_l[8]),
    .ts(1'b1),
    .di(limit_l_pad[8]));  // CPLD_SOC_AHB_TOP.v(5)
  // src/AHB.v(48)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u811|U_AHB/reg3_b15  (
    .a({\PWM2/FreCnt [0],_al_u811_o}),
    .b({\PWM2/FreCnt [1],\PWM2/FreCnt [12]}),
    .c({\PWM2/FreCnt [10],\PWM2/FreCnt [13]}),
    .ce(\U_AHB/n8 ),
    .clk(clk100m),
    .d({\PWM2/FreCnt [11],\PWM2/FreCnt [14]}),
    .e({open_n40432,\PWM2/FreCnt [15]}),
    .mi({open_n40434,\U_AHB/h2h_hwdata [15]}),
    .f({_al_u811_o,_al_u812_o}),
    .q({open_n40450,freq2[15]}));  // src/AHB.v(48)
  EF2_PHY_SPAD #(
    //.LOCATION("P89"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u82 (
    .ipad(limit_l[7]),
    .ts(1'b1),
    .di(limit_l_pad[7]));  // CPLD_SOC_AHB_TOP.v(5)
  EF2_PHY_SPAD #(
    //.LOCATION("P2"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u83 (
    .ipad(limit_l[6]),
    .ts(1'b1),
    .di(limit_l_pad[6]));  // CPLD_SOC_AHB_TOP.v(5)
  EF2_PHY_SPAD #(
    //.LOCATION("P6"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u84 (
    .ipad(limit_l[5]),
    .ts(1'b1),
    .di(limit_l_pad[5]));  // CPLD_SOC_AHB_TOP.v(5)
  // src/AHB.v(49)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u848|U_AHB/reg4_b1  (
    .a({\PWM3/FreCnt [0],_al_u1427_o}),
    .b({\PWM3/FreCnt [1],\PWM3/FreCnt [1]}),
    .c({\PWM3/FreCnt [10],\PWM3/FreCnt [10]}),
    .ce(\U_AHB/n10 ),
    .clk(clk100m),
    .d({\PWM3/FreCnt [11],\PWM3/FreCntr [1]}),
    .e({open_n40478,\PWM3/FreCntr [10]}),
    .mi({open_n40480,\U_AHB/h2h_hwdata [1]}),
    .f({_al_u848_o,_al_u1428_o}),
    .q({open_n40496,freq3[1]}));  // src/AHB.v(49)
  // src/OnePWM.v(37)
  EF2_PHY_LSLICE #(
    //.LUTF0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D)"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111000011001100),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b1111000011001100),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u849|PWM3/reg0_b15  (
    .a({_al_u848_o,open_n40497}),
    .b({\PWM3/FreCnt [12],\PWM3/n12 [15]}),
    .c({\PWM3/FreCnt [13],freq3[15]}),
    .clk(clk100m),
    .d({\PWM3/FreCnt [14],\PWM3/n0_lutinv }),
    .e({\PWM3/FreCnt [15],open_n40499}),
    .sr(\PWM3/n11 ),
    .f({_al_u849_o,open_n40514}),
    .q({open_n40518,\PWM3/FreCnt [15]}));  // src/OnePWM.v(37)
  EF2_PHY_PAD #(
    //.LOCATION("P60"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u85 (
    .ipad(limit_l[4]),
    .di(limit_l_pad[4]));  // CPLD_SOC_AHB_TOP.v(5)
  // src/AHB.v(49)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~0*~D*~C*~B*A)"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(~1*~D*~C*~B*A)"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000010),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b0000000000000000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u850|U_AHB/reg4_b22  (
    .a({\PWM3/FreCnt [16],_al_u850_o}),
    .b({\PWM3/FreCnt [17],\PWM3/FreCnt [2]}),
    .c({\PWM3/FreCnt [18],\PWM3/FreCnt [20]}),
    .ce(\U_AHB/n10 ),
    .clk(clk100m),
    .d({\PWM3/FreCnt [19],\PWM3/FreCnt [21]}),
    .e({open_n40542,\PWM3/FreCnt [22]}),
    .mi({open_n40544,\U_AHB/h2h_hwdata [22]}),
    .f({_al_u850_o,_al_u851_o}),
    .q({open_n40560,freq3[22]}));  // src/AHB.v(49)
  EF2_PHY_PAD #(
    //.LOCATION("P58"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u86 (
    .ipad(limit_l[3]),
    .di(limit_l_pad[3]));  // CPLD_SOC_AHB_TOP.v(5)
  EF2_PHY_PAD #(
    //.LOCATION("P56"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u87 (
    .ipad(limit_l[2]),
    .di(limit_l_pad[2]));  // CPLD_SOC_AHB_TOP.v(5)
  EF2_PHY_PAD #(
    //.LOCATION("P50"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u88 (
    .ipad(limit_l[1]),
    .di(limit_l_pad[1]));  // CPLD_SOC_AHB_TOP.v(5)
  // src/AHB.v(50)
  EF2_PHY_LSLICE #(
    //.LUTF0("(~(~C*B)*~(~D*A))"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(~(~C*B)*~(~D*A))"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1111001101010001),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b1111001101010001),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u885|U_AHB/reg5_b13  (
    .a({\PWM4/FreCnt [0],\PWM4/FreCnt [1]}),
    .b({\PWM4/FreCnt [1],\PWM4/FreCnt [12]}),
    .c({\PWM4/FreCnt [10],\PWM4/FreCntr [13]}),
    .ce(\U_AHB/n12 ),
    .clk(clk100m),
    .d({\PWM4/FreCnt [11],\PWM4/FreCntr [2]}),
    .mi({open_n40633,\U_AHB/h2h_hwdata [13]}),
    .f({_al_u885_o,_al_u2067_o}),
    .q({open_n40649,freq4[13]}));  // src/AHB.v(50)
  // src/AHB.v(84)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u886|U_AHB/reg34_b4  (
    .a({_al_u885_o,open_n40650}),
    .b({\PWM4/FreCnt [12],_al_u886_o}),
    .c({\PWM4/FreCnt [13],_al_u888_o}),
    .clk(clk100m),
    .d({\PWM4/FreCnt [14],_al_u884_o}),
    .e({\PWM4/FreCnt [15],open_n40652}),
    .mi({open_n40654,\U_AHB/h2h_hwdata [4]}),
    .sr(\U_AHB/n79 ),
    .f({_al_u886_o,\PWM4/n0_lutinv }),
    .q({open_n40669,pwm_start_stop[4]}));  // src/AHB.v(84)
  EF2_PHY_PAD #(
    //.LOCATION("P41"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u89 (
    .ipad(limit_l[0]),
    .di(limit_l_pad[0]));  // CPLD_SOC_AHB_TOP.v(5)
  EF2_PHY_SPAD #(
    //.LOCATION("P95"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u90 (
    .ipad(limit_r[15]),
    .ts(1'b1),
    .di(limit_r_pad[15]));  // CPLD_SOC_AHB_TOP.v(6)
  EF2_PHY_SPAD #(
    //.LOCATION("P81"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u91 (
    .ipad(limit_r[14]),
    .ts(1'b1),
    .di(limit_r_pad[14]));  // CPLD_SOC_AHB_TOP.v(6)
  EF2_PHY_SPAD #(
    //.LOCATION("P3"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u92 (
    .ipad(limit_r[13]),
    .ts(1'b1),
    .di(limit_r_pad[13]));  // CPLD_SOC_AHB_TOP.v(6)
  // src/AHB.v(51)
  EF2_PHY_LSLICE #(
    //.LUTF0("(A*~(0@C)*~(D@B))"),
    //.LUTF1("(~D*~C*~B*~A)"),
    //.LUTG0("(A*~(1@C)*~(D@B))"),
    //.LUTG1("(~D*~C*~B*~A)"),
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000100000000010),
    .INIT_LUTF1(16'b0000000000000001),
    .INIT_LUTG0(16'b1000000000100000),
    .INIT_LUTG1(16'b0000000000000001),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \_al_u922|U_AHB/reg6_b11  (
    .a({\PWM5/FreCnt [0],_al_u1459_o}),
    .b({\PWM5/FreCnt [1],\PWM5/FreCnt [11]}),
    .c({\PWM5/FreCnt [10],\PWM5/FreCnt [25]}),
    .ce(\U_AHB/n14 ),
    .clk(clk100m),
    .d({\PWM5/FreCnt [11],\PWM5/FreCntr [11]}),
    .e({open_n40720,\PWM5/FreCntr [25]}),
    .mi({open_n40722,\U_AHB/h2h_hwdata [11]}),
    .f({_al_u922_o,_al_u1460_o}),
    .q({open_n40738,freq5[11]}));  // src/AHB.v(51)
  // src/AHB.v(84)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*B*D)"),
    //.LUTF1("(~0*~D*~C*~B*A)"),
    //.LUTG0("(C*B*D)"),
    //.LUTG1("(~1*~D*~C*~B*A)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b1100000000000000),
    .INIT_LUTF1(16'b0000000000000010),
    .INIT_LUTG0(16'b1100000000000000),
    .INIT_LUTG1(16'b0000000000000000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \_al_u923|U_AHB/reg34_b5  (
    .a({_al_u922_o,open_n40739}),
    .b({\PWM5/FreCnt [12],_al_u923_o}),
    .c({\PWM5/FreCnt [13],_al_u925_o}),
    .clk(clk100m),
    .d({\PWM5/FreCnt [14],_al_u921_o}),
    .e({\PWM5/FreCnt [15],open_n40741}),
    .mi({open_n40743,\U_AHB/h2h_hwdata [5]}),
    .sr(\U_AHB/n79 ),
    .f({_al_u923_o,\PWM5/n0_lutinv }),
    .q({open_n40758,pwm_start_stop[5]}));  // src/AHB.v(84)
  EF2_PHY_SPAD #(
    //.LOCATION("P5"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u93 (
    .ipad(limit_r[12]),
    .ts(1'b1),
    .di(limit_r_pad[12]));  // CPLD_SOC_AHB_TOP.v(6)
  EF2_PHY_PAD #(
    //.LOCATION("P68"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u94 (
    .ipad(limit_r[11]),
    .di(limit_r_pad[11]));  // CPLD_SOC_AHB_TOP.v(6)
  EF2_PHY_SPAD #(
    //.LOCATION("P35"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u95 (
    .ipad(limit_r[10]),
    .ts(1'b1),
    .di(limit_r_pad[10]));  // CPLD_SOC_AHB_TOP.v(6)
  EF2_PHY_SPAD #(
    //.LOCATION("P94"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u96 (
    .ipad(limit_r[9]),
    .ts(1'b1),
    .di(limit_r_pad[9]));  // CPLD_SOC_AHB_TOP.v(6)
  EF2_PHY_SPAD #(
    //.LOCATION("P86"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u97 (
    .ipad(limit_r[8]),
    .ts(1'b1),
    .di(limit_r_pad[8]));  // CPLD_SOC_AHB_TOP.v(6)
  EF2_PHY_SPAD #(
    //.LOCATION("P82"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u98 (
    .ipad(limit_r[7]),
    .ts(1'b1),
    .di(limit_r_pad[7]));  // CPLD_SOC_AHB_TOP.v(6)
  EF2_PHY_SPAD #(
    //.LOCATION("P4"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u99 (
    .ipad(limit_r[6]),
    .ts(1'b1),
    .di(limit_r_pad[6]));  // CPLD_SOC_AHB_TOP.v(6)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    _bufkeep_clk100m (
    .i(clk100m_keep),
    .o(clk100m));  // CPLD_SOC_AHB_TOP.v(13)
  EF2_PHY_LSLICE #(
    //.MACRO("add0/ucin_al_u3354"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \add0/u11_al_u3357  (
    .a({timer[13],timer[11]}),
    .b({timer[14],timer[12]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\add0/c11 ),
    .f({n2[13],n2[11]}),
    .fco(\add0/c15 ),
    .fx({n2[14],n2[12]}));
  EF2_PHY_LSLICE #(
    //.MACRO("add0/ucin_al_u3354"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \add0/u15_al_u3358  (
    .a({timer[17],timer[15]}),
    .b({timer[18],timer[16]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\add0/c15 ),
    .f({n2[17],n2[15]}),
    .fco(\add0/c19 ),
    .fx({n2[18],n2[16]}));
  EF2_PHY_LSLICE #(
    //.MACRO("add0/ucin_al_u3354"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \add0/u19_al_u3359  (
    .a({timer[21],timer[19]}),
    .b({timer[22],timer[20]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\add0/c19 ),
    .f({n2[21],n2[19]}),
    .fco(\add0/c23 ),
    .fx({n2[22],n2[20]}));
  EF2_PHY_LSLICE #(
    //.MACRO("add0/ucin_al_u3354"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \add0/u23_al_u3360  (
    .a({timer[25],timer[23]}),
    .b({timer[26],timer[24]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\add0/c23 ),
    .f({n2[25],n2[23]}),
    .fco(\add0/c27 ),
    .fx({n2[26],n2[24]}));
  EF2_PHY_LSLICE #(
    //.MACRO("add0/ucin_al_u3354"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \add0/u27_al_u3361  (
    .a({timer[29],timer[27]}),
    .b({timer[30],timer[28]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\add0/c27 ),
    .f({n2[29],n2[27]}),
    .fco(\add0/c31 ),
    .fx({n2[30],n2[28]}));
  EF2_PHY_LSLICE #(
    //.MACRO("add0/ucin_al_u3354"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \add0/u31_al_u3362  (
    .a({open_n40926,timer[31]}),
    .c(2'b00),
    .d({open_n40931,1'b0}),
    .fci(\add0/c31 ),
    .f({open_n40948,n2[31]}));
  EF2_PHY_LSLICE #(
    //.MACRO("add0/ucin_al_u3354"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \add0/u3_al_u3355  (
    .a({timer[5],timer[3]}),
    .b({timer[6],timer[4]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\add0/c3 ),
    .f({n2[5],n2[3]}),
    .fco(\add0/c7 ),
    .fx({n2[6],n2[4]}));
  EF2_PHY_LSLICE #(
    //.MACRO("add0/ucin_al_u3354"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \add0/u7_al_u3356  (
    .a({timer[9],timer[7]}),
    .b({timer[10],timer[8]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\add0/c7 ),
    .f({n2[9],n2[7]}),
    .fco(\add0/c11 ),
    .fx({n2[10],n2[8]}));
  EF2_PHY_LSLICE #(
    //.MACRO("add0/ucin_al_u3354"),
    //.R_POSITION("X0Y0Z0"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"),
    .REG0_REGSET("RESET"),
    .REG0_SD("MI"),
    .REG1_REGSET("RESET"),
    .REG1_SD("MI"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \add0/ucin_al_u3354  (
    .a({timer[1],1'b0}),
    .b({timer[2],timer[0]}),
    .c(2'b00),
    .clk(clk100m),
    .d(2'b01),
    .e(2'b01),
    .mi(\U_AHB/h2h_hwdata [28:27]),
    .sr(\U_AHB/n73 ),
    .f({n2[1],open_n41003}),
    .fco(\add0/c3 ),
    .fx({n2[2],n2[0]}),
    .q(pnumD[28:27]));
  EF2_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  EF2_PHY_LSLICE #(
    //.LUTF0("(0*D*C*B*A)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(1*D*C*B*A)"),
    //.LUTG1("(C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \reg0_b0|_al_u2978  (
    .a({open_n41051,_al_u2963_o}),
    .b({open_n41052,_al_u2970_o}),
    .c({n2[0],_al_u2973_o}),
    .clk(clk25m),
    .d({_al_u1652_o,_al_u2975_o}),
    .e({open_n41054,_al_u2977_o}),
    .sr(rst_n_pad),
    .f({open_n41069,_al_u2978_o}),
    .q({timer[0],open_n41073}));  // CPLD_SOC_AHB_TOP.v(35)
  EF2_PHY_LSLICE #(
    //.LUTF0("(0*D*C*B*A)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(1*D*C*B*A)"),
    //.LUTG1("(C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000000000000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b1000000000000000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \reg0_b10|_al_u2173  (
    .a({open_n41074,_al_u2157_o}),
    .b({open_n41075,_al_u2164_o}),
    .c({n2[10],_al_u2168_o}),
    .clk(clk25m),
    .d({_al_u1652_o,_al_u2170_o}),
    .e({open_n41077,_al_u2172_o}),
    .sr(rst_n_pad),
    .f({open_n41092,_al_u2173_o}),
    .q({timer[10],open_n41096}));  // CPLD_SOC_AHB_TOP.v(35)
  // CPLD_SOC_AHB_TOP.v(35)
  // CPLD_SOC_AHB_TOP.v(35)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \reg0_b11|reg0_b27  (
    .c({n2[11],n2[27]}),
    .clk(clk25m),
    .d({_al_u1652_o,_al_u1652_o}),
    .sr(rst_n_pad),
    .q({timer[11],timer[27]}));  // CPLD_SOC_AHB_TOP.v(35)
  // CPLD_SOC_AHB_TOP.v(35)
  // CPLD_SOC_AHB_TOP.v(35)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \reg0_b12|reg0_b26  (
    .c({n2[12],n2[26]}),
    .clk(clk25m),
    .d({_al_u1652_o,_al_u1652_o}),
    .sr(rst_n_pad),
    .q({timer[12],timer[26]}));  // CPLD_SOC_AHB_TOP.v(35)
  // CPLD_SOC_AHB_TOP.v(35)
  // CPLD_SOC_AHB_TOP.v(35)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \reg0_b13|reg0_b25  (
    .c({n2[13],n2[25]}),
    .clk(clk25m),
    .d({_al_u1652_o,_al_u1652_o}),
    .sr(rst_n_pad),
    .q({timer[13],timer[25]}));  // CPLD_SOC_AHB_TOP.v(35)
  // CPLD_SOC_AHB_TOP.v(35)
  // CPLD_SOC_AHB_TOP.v(35)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \reg0_b14|reg0_b24  (
    .c({n2[14],n2[24]}),
    .clk(clk25m),
    .d({_al_u1652_o,_al_u1652_o}),
    .sr(rst_n_pad),
    .q({timer[14],timer[24]}));  // CPLD_SOC_AHB_TOP.v(35)
  // CPLD_SOC_AHB_TOP.v(35)
  // CPLD_SOC_AHB_TOP.v(35)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \reg0_b15|reg0_b17  (
    .c({n2[15],n2[17]}),
    .clk(clk25m),
    .d({_al_u1652_o,_al_u1652_o}),
    .sr(rst_n_pad),
    .q({timer[15],timer[17]}));  // CPLD_SOC_AHB_TOP.v(35)
  // CPLD_SOC_AHB_TOP.v(35)
  // CPLD_SOC_AHB_TOP.v(35)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \reg0_b18|reg0_b16  (
    .c({n2[18],n2[16]}),
    .clk(clk25m),
    .d({_al_u1652_o,_al_u1652_o}),
    .sr(rst_n_pad),
    .q({timer[18],timer[16]}));  // CPLD_SOC_AHB_TOP.v(35)
  // CPLD_SOC_AHB_TOP.v(35)
  // CPLD_SOC_AHB_TOP.v(35)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \reg0_b1|reg0_b19  (
    .c({n2[1],n2[19]}),
    .clk(clk25m),
    .d({_al_u1652_o,_al_u1652_o}),
    .sr(rst_n_pad),
    .q({timer[1],timer[19]}));  // CPLD_SOC_AHB_TOP.v(35)
  // CPLD_SOC_AHB_TOP.v(35)
  // CPLD_SOC_AHB_TOP.v(35)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \reg0_b20|reg0_b8  (
    .c({n2[20],n2[8]}),
    .clk(clk25m),
    .d({_al_u1652_o,_al_u1652_o}),
    .sr(rst_n_pad),
    .q({timer[20],timer[8]}));  // CPLD_SOC_AHB_TOP.v(35)
  // CPLD_SOC_AHB_TOP.v(35)
  // CPLD_SOC_AHB_TOP.v(35)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \reg0_b21|reg0_b7  (
    .c({n2[21],n2[7]}),
    .clk(clk25m),
    .d({_al_u1652_o,_al_u1652_o}),
    .sr(rst_n_pad),
    .q({timer[21],timer[7]}));  // CPLD_SOC_AHB_TOP.v(35)
  // CPLD_SOC_AHB_TOP.v(35)
  // CPLD_SOC_AHB_TOP.v(35)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \reg0_b22|reg0_b6  (
    .c({n2[22],n2[6]}),
    .clk(clk25m),
    .d({_al_u1652_o,_al_u1652_o}),
    .sr(rst_n_pad),
    .q({timer[22],timer[6]}));  // CPLD_SOC_AHB_TOP.v(35)
  // CPLD_SOC_AHB_TOP.v(35)
  // CPLD_SOC_AHB_TOP.v(35)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \reg0_b23|reg0_b5  (
    .c({n2[23],n2[5]}),
    .clk(clk25m),
    .d({_al_u1652_o,_al_u1652_o}),
    .sr(rst_n_pad),
    .q({timer[23],timer[5]}));  // CPLD_SOC_AHB_TOP.v(35)
  // CPLD_SOC_AHB_TOP.v(35)
  // CPLD_SOC_AHB_TOP.v(35)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \reg0_b28|reg0_b4  (
    .c({n2[28],n2[4]}),
    .clk(clk25m),
    .d({_al_u1652_o,_al_u1652_o}),
    .sr(rst_n_pad),
    .q({timer[28],timer[4]}));  // CPLD_SOC_AHB_TOP.v(35)
  // CPLD_SOC_AHB_TOP.v(35)
  // CPLD_SOC_AHB_TOP.v(35)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \reg0_b29|reg0_b9  (
    .c({n2[29],n2[9]}),
    .clk(clk25m),
    .d({_al_u1652_o,_al_u1652_o}),
    .sr(rst_n_pad),
    .q({timer[29],timer[9]}));  // CPLD_SOC_AHB_TOP.v(35)
  // CPLD_SOC_AHB_TOP.v(35)
  // CPLD_SOC_AHB_TOP.v(35)
  EF2_PHY_LSLICE #(
    //.LUTF0("(C*~D)"),
    //.LUTF1("(C*~D)"),
    //.LUTG0("(C*~D)"),
    //.LUTG1("(C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUTF0(16'b0000000011110000),
    .INIT_LUTF1(16'b0000000011110000),
    .INIT_LUTG0(16'b0000000011110000),
    .INIT_LUTG1(16'b0000000011110000),
    .LSFMUX0("FUNC5"),
    .LSFMUX1("FUNC5"),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \reg0_b2|reg0_b31  (
    .c({n2[2],n2[31]}),
    .clk(clk25m),
    .d({_al_u1652_o,_al_u1652_o}),
    .sr(rst_n_pad),
    .q({timer[2],timer[31]}));  // CPLD_SOC_AHB_TOP.v(35)
  // CPLD_SOC_AHB_TOP.v(35)
  // CPLD_SOC_AHB_TOP.v(35)
  EF2_PHY_MSLICE #(
    //.LUT0("(C*~D)"),
    //.LUT1("(C*~D)"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b0000000011110000),
    .INIT_LUT1(16'b0000000011110000),
    .MODE("LOGIC"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \reg0_b3|reg0_b30  (
    .c({n2[3],n2[30]}),
    .clk(clk25m),
    .d({_al_u1652_o,_al_u1652_o}),
    .sr(rst_n_pad),
    .q({timer[3],timer[30]}));  // CPLD_SOC_AHB_TOP.v(35)
  EF2_PHY_SPAD #(
    //.CLKSRC("CLK"),
    //.LOCATION("P105"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DO_DFFMODE("FF"),
    .DO_REGSET("SET"),
    .DRIVE("16"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .OUTCEMUX("CE"),
    .OUTCLKMUX("CLK"),
    .OUTRSTMUX("INV"),
    .SRMODE("ASYNC"),
    .TSMUX("INV"))
    reg1_b0_DO (
    .ce(_al_n1_en),
    .clk(clk25m),
    .do({open_n41459,n4_neg}),
    .rst(rst_n_pad),
    .ts(1'b1),
    .opad(ledout[0]));  // CPLD_SOC_AHB_TOP.v(49)
  // CPLD_SOC_AHB_TOP.v(49)
  // CPLD_SOC_AHB_TOP.v(49)
  EF2_PHY_MSLICE #(
    //.LUT0("~(~C*A*~(D*~B))"),
    //.LUT1("~(A*~(~C*~(~D*~B)))"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1111011111110101),
    .INIT_LUT1(16'b0101111101011101),
    .MODE("LOGIC"),
    .REG0_REGSET("SET"),
    .REG0_SD("F"),
    .REG1_REGSET("SET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \reg1_b2|reg1_b3  (
    .a({_al_u2984_o,_al_u2984_o}),
    .b({_al_u1652_o,_al_u1652_o}),
    .c({_al_u2988_o,_al_u2988_o}),
    .clk(clk25m),
    .d({ledout_pad[2],ledout_pad[3]}),
    .sr(rst_n_pad),
    .q({ledout_pad[2],ledout_pad[3]}));  // CPLD_SOC_AHB_TOP.v(49)

endmodule 

module AL_BUFKEEP
  (
  i,
  o
  );

  input i;
  output o;

  parameter KEEP = "OUT";

  buf u1 (o, i);

endmodule 

