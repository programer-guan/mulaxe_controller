// Verilog netlist created by TD v4.5.12562
// Thu Dec 19 17:42:02 2019

`timescale 1ns / 1ps
module CPLD_SOC_AHB_TOP  // CPLD_SOC_AHB_TOP.v(1)
  (
  clkin,
  limit_l,
  limit_r,
  rst_n,
  dir,
  gpio_out,
  ledout,
  pwm
  );

  input clkin;  // CPLD_SOC_AHB_TOP.v(3)
  input [15:0] limit_l;  // CPLD_SOC_AHB_TOP.v(5)
  input [15:0] limit_r;  // CPLD_SOC_AHB_TOP.v(6)
  input rst_n;  // CPLD_SOC_AHB_TOP.v(4)
  output [15:0] dir;  // CPLD_SOC_AHB_TOP.v(7)
  output [31:0] gpio_out;  // CPLD_SOC_AHB_TOP.v(8)
  output [3:0] ledout;  // CPLD_SOC_AHB_TOP.v(10)
  output [15:0] pwm;  // CPLD_SOC_AHB_TOP.v(7)

  wire [26:0] \PWM0/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWM0/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWM0/n12 ;
  wire [26:0] \PWM0/n13 ;
  wire [31:0] \PWM0/n23 ;
  wire [24:0] \PWM0/n26 ;
  wire [23:0] \PWM0/n31 ;
  wire [31:0] \PWM0/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWM1/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWM1/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWM1/n12 ;
  wire [26:0] \PWM1/n13 ;
  wire [31:0] \PWM1/n23 ;
  wire [24:0] \PWM1/n26 ;
  wire [23:0] \PWM1/n31 ;
  wire [31:0] \PWM1/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWM2/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWM2/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWM2/n12 ;
  wire [26:0] \PWM2/n13 ;
  wire [31:0] \PWM2/n23 ;
  wire [24:0] \PWM2/n26 ;
  wire [23:0] \PWM2/n31 ;
  wire [31:0] \PWM2/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWM3/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWM3/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWM3/n12 ;
  wire [26:0] \PWM3/n13 ;
  wire [31:0] \PWM3/n23 ;
  wire [24:0] \PWM3/n26 ;
  wire [23:0] \PWM3/n31 ;
  wire [31:0] \PWM3/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWM4/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWM4/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWM4/n12 ;
  wire [26:0] \PWM4/n13 ;
  wire [31:0] \PWM4/n23 ;
  wire [24:0] \PWM4/n26 ;
  wire [23:0] \PWM4/n31 ;
  wire [31:0] \PWM4/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWM5/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWM5/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWM5/n12 ;
  wire [26:0] \PWM5/n13 ;
  wire [31:0] \PWM5/n23 ;
  wire [24:0] \PWM5/n26 ;
  wire [23:0] \PWM5/n31 ;
  wire [31:0] \PWM5/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWM6/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWM6/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWM6/n12 ;
  wire [26:0] \PWM6/n13 ;
  wire [31:0] \PWM6/n23 ;
  wire [24:0] \PWM6/n26 ;
  wire [23:0] \PWM6/n31 ;
  wire [31:0] \PWM6/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWM7/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWM7/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWM7/n12 ;
  wire [26:0] \PWM7/n13 ;
  wire [31:0] \PWM7/n23 ;
  wire [24:0] \PWM7/n26 ;
  wire [23:0] \PWM7/n31 ;
  wire [31:0] \PWM7/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWM8/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWM8/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWM8/n12 ;
  wire [26:0] \PWM8/n13 ;
  wire [31:0] \PWM8/n23 ;
  wire [24:0] \PWM8/n26 ;
  wire [23:0] \PWM8/n31 ;
  wire [31:0] \PWM8/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWM9/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWM9/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWM9/n12 ;
  wire [26:0] \PWM9/n13 ;
  wire [31:0] \PWM9/n23 ;
  wire [24:0] \PWM9/n26 ;
  wire [23:0] \PWM9/n31 ;
  wire [31:0] \PWM9/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWMA/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWMA/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWMA/n12 ;
  wire [26:0] \PWMA/n13 ;
  wire [31:0] \PWMA/n23 ;
  wire [24:0] \PWMA/n26 ;
  wire [23:0] \PWMA/n31 ;
  wire [31:0] \PWMA/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWMB/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWMB/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWMB/n12 ;
  wire [26:0] \PWMB/n13 ;
  wire [31:0] \PWMB/n23 ;
  wire [24:0] \PWMB/n26 ;
  wire [23:0] \PWMB/n31 ;
  wire [31:0] \PWMB/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWMC/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWMC/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWMC/n12 ;
  wire [26:0] \PWMC/n13 ;
  wire [31:0] \PWMC/n23 ;
  wire [24:0] \PWMC/n26 ;
  wire [23:0] \PWMC/n31 ;
  wire [31:0] \PWMC/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWMD/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWMD/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWMD/n12 ;
  wire [26:0] \PWMD/n13 ;
  wire [31:0] \PWMD/n23 ;
  wire [24:0] \PWMD/n26 ;
  wire [23:0] \PWMD/n31 ;
  wire [31:0] \PWMD/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWME/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWME/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWME/n12 ;
  wire [26:0] \PWME/n13 ;
  wire [31:0] \PWME/n23 ;
  wire [24:0] \PWME/n26 ;
  wire [23:0] \PWME/n31 ;
  wire [31:0] \PWME/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWMF/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWMF/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWMF/n12 ;
  wire [26:0] \PWMF/n13 ;
  wire [31:0] \PWMF/n23 ;
  wire [24:0] \PWMF/n26 ;
  wire [23:0] \PWMF/n31 ;
  wire [31:0] \PWMF/pnumr ;  // src/OnePWM.v(47)
  wire [31:0] \U_AHB/h2h_haddr ;  // src/AHB.v(23)
  wire [31:0] \U_AHB/h2h_haddrw ;  // src/AHB.v(16)
  wire [31:0] \U_AHB/h2h_hrdata ;  // src/AHB.v(18)
  wire [31:0] \U_AHB/h2h_hwdata ;  // src/AHB.v(17)
  wire [31:0] \U_AHB/n118 ;
  wire [31:0] \U_AHB/n42 ;
  wire [15:0] dir_pad;  // CPLD_SOC_AHB_TOP.v(7)
  wire [31:0] freq0;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freq1;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freq2;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freq3;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freq4;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freq5;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freq6;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freq7;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freq8;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freq9;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freqA;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freqB;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freqC;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freqD;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freqE;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freqF;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] gpio_out_pad;  // CPLD_SOC_AHB_TOP.v(8)
  wire [3:0] ledout_pad;  // CPLD_SOC_AHB_TOP.v(10)
  wire [15:0] limit_l_pad;  // CPLD_SOC_AHB_TOP.v(5)
  wire [15:0] limit_r_pad;  // CPLD_SOC_AHB_TOP.v(6)
  wire [3:0] n10;
  wire [31:0] n2;
  wire [31:0] n3;
  wire [32:0] pnum0;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnum1;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnum2;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnum3;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnum4;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnum5;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnum6;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnum7;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnum8;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnum9;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnumA;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnumB;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnumC;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnumD;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnumE;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnumF;  // CPLD_SOC_AHB_TOP.v(54)
  wire [23:0] pnumcnt0;  // CPLD_SOC_AHB_TOP.v(61)
  wire [23:0] pnumcnt1;  // CPLD_SOC_AHB_TOP.v(62)
  wire [23:0] pnumcnt2;  // CPLD_SOC_AHB_TOP.v(63)
  wire [23:0] pnumcnt3;  // CPLD_SOC_AHB_TOP.v(64)
  wire [23:0] pnumcnt4;  // CPLD_SOC_AHB_TOP.v(65)
  wire [23:0] pnumcnt5;  // CPLD_SOC_AHB_TOP.v(66)
  wire [23:0] pnumcnt6;  // CPLD_SOC_AHB_TOP.v(67)
  wire [23:0] pnumcnt7;  // CPLD_SOC_AHB_TOP.v(68)
  wire [23:0] pnumcnt8;  // CPLD_SOC_AHB_TOP.v(69)
  wire [23:0] pnumcnt9;  // CPLD_SOC_AHB_TOP.v(70)
  wire [23:0] pnumcntA;  // CPLD_SOC_AHB_TOP.v(71)
  wire [23:0] pnumcntB;  // CPLD_SOC_AHB_TOP.v(72)
  wire [23:0] pnumcntC;  // CPLD_SOC_AHB_TOP.v(73)
  wire [23:0] pnumcntD;  // CPLD_SOC_AHB_TOP.v(74)
  wire [23:0] pnumcntE;  // CPLD_SOC_AHB_TOP.v(75)
  wire [23:0] pnumcntF;  // CPLD_SOC_AHB_TOP.v(76)
  wire [15:0] pwm_pad;  // CPLD_SOC_AHB_TOP.v(7)
  wire [31:0] pwm_start_stop;  // CPLD_SOC_AHB_TOP.v(52)
  wire [15:0] pwm_state_read;  // CPLD_SOC_AHB_TOP.v(78)
  wire [31:0] timer;  // CPLD_SOC_AHB_TOP.v(26)
  wire \PWM0/RemaTxNum[0]_keep ;
  wire \PWM0/RemaTxNum[10]_keep ;
  wire \PWM0/RemaTxNum[11]_keep ;
  wire \PWM0/RemaTxNum[12]_keep ;
  wire \PWM0/RemaTxNum[13]_keep ;
  wire \PWM0/RemaTxNum[14]_keep ;
  wire \PWM0/RemaTxNum[15]_keep ;
  wire \PWM0/RemaTxNum[16]_keep ;
  wire \PWM0/RemaTxNum[17]_keep ;
  wire \PWM0/RemaTxNum[18]_keep ;
  wire \PWM0/RemaTxNum[19]_keep ;
  wire \PWM0/RemaTxNum[1]_keep ;
  wire \PWM0/RemaTxNum[20]_keep ;
  wire \PWM0/RemaTxNum[21]_keep ;
  wire \PWM0/RemaTxNum[22]_keep ;
  wire \PWM0/RemaTxNum[23]_keep ;
  wire \PWM0/RemaTxNum[2]_keep ;
  wire \PWM0/RemaTxNum[3]_keep ;
  wire \PWM0/RemaTxNum[4]_keep ;
  wire \PWM0/RemaTxNum[5]_keep ;
  wire \PWM0/RemaTxNum[6]_keep ;
  wire \PWM0/RemaTxNum[7]_keep ;
  wire \PWM0/RemaTxNum[8]_keep ;
  wire \PWM0/RemaTxNum[9]_keep ;
  wire \PWM0/dir_keep ;
  wire \PWM0/mux3_b0_sel_is_3_o ;
  wire \PWM0/n0_lutinv ;
  wire \PWM0/n1 ;
  wire \PWM0/n10 ;
  wire \PWM0/n11 ;
  wire \PWM0/n24 ;
  wire \PWM0/n25_neg_lutinv ;
  wire \PWM0/n32 ;
  wire \PWM0/pnumr[0]_keep ;
  wire \PWM0/pnumr[10]_keep ;
  wire \PWM0/pnumr[11]_keep ;
  wire \PWM0/pnumr[12]_keep ;
  wire \PWM0/pnumr[13]_keep ;
  wire \PWM0/pnumr[14]_keep ;
  wire \PWM0/pnumr[15]_keep ;
  wire \PWM0/pnumr[16]_keep ;
  wire \PWM0/pnumr[17]_keep ;
  wire \PWM0/pnumr[18]_keep ;
  wire \PWM0/pnumr[19]_keep ;
  wire \PWM0/pnumr[1]_keep ;
  wire \PWM0/pnumr[20]_keep ;
  wire \PWM0/pnumr[21]_keep ;
  wire \PWM0/pnumr[22]_keep ;
  wire \PWM0/pnumr[23]_keep ;
  wire \PWM0/pnumr[24]_keep ;
  wire \PWM0/pnumr[25]_keep ;
  wire \PWM0/pnumr[26]_keep ;
  wire \PWM0/pnumr[27]_keep ;
  wire \PWM0/pnumr[28]_keep ;
  wire \PWM0/pnumr[29]_keep ;
  wire \PWM0/pnumr[2]_keep ;
  wire \PWM0/pnumr[30]_keep ;
  wire \PWM0/pnumr[31]_keep ;
  wire \PWM0/pnumr[3]_keep ;
  wire \PWM0/pnumr[4]_keep ;
  wire \PWM0/pnumr[5]_keep ;
  wire \PWM0/pnumr[6]_keep ;
  wire \PWM0/pnumr[7]_keep ;
  wire \PWM0/pnumr[8]_keep ;
  wire \PWM0/pnumr[9]_keep ;
  wire \PWM0/pwm_keep ;
  wire \PWM0/stopreq ;  // src/OnePWM.v(14)
  wire \PWM0/stopreq_keep ;
  wire \PWM0/sub0/c0 ;
  wire \PWM0/sub0/c1 ;
  wire \PWM0/sub0/c10 ;
  wire \PWM0/sub0/c11 ;
  wire \PWM0/sub0/c12 ;
  wire \PWM0/sub0/c13 ;
  wire \PWM0/sub0/c14 ;
  wire \PWM0/sub0/c15 ;
  wire \PWM0/sub0/c16 ;
  wire \PWM0/sub0/c17 ;
  wire \PWM0/sub0/c18 ;
  wire \PWM0/sub0/c19 ;
  wire \PWM0/sub0/c2 ;
  wire \PWM0/sub0/c20 ;
  wire \PWM0/sub0/c21 ;
  wire \PWM0/sub0/c22 ;
  wire \PWM0/sub0/c23 ;
  wire \PWM0/sub0/c24 ;
  wire \PWM0/sub0/c25 ;
  wire \PWM0/sub0/c26 ;
  wire \PWM0/sub0/c3 ;
  wire \PWM0/sub0/c4 ;
  wire \PWM0/sub0/c5 ;
  wire \PWM0/sub0/c6 ;
  wire \PWM0/sub0/c7 ;
  wire \PWM0/sub0/c8 ;
  wire \PWM0/sub0/c9 ;
  wire \PWM0/sub1/c0 ;
  wire \PWM0/sub1/c1 ;
  wire \PWM0/sub1/c10 ;
  wire \PWM0/sub1/c11 ;
  wire \PWM0/sub1/c12 ;
  wire \PWM0/sub1/c13 ;
  wire \PWM0/sub1/c14 ;
  wire \PWM0/sub1/c15 ;
  wire \PWM0/sub1/c16 ;
  wire \PWM0/sub1/c17 ;
  wire \PWM0/sub1/c18 ;
  wire \PWM0/sub1/c19 ;
  wire \PWM0/sub1/c2 ;
  wire \PWM0/sub1/c20 ;
  wire \PWM0/sub1/c21 ;
  wire \PWM0/sub1/c22 ;
  wire \PWM0/sub1/c23 ;
  wire \PWM0/sub1/c3 ;
  wire \PWM0/sub1/c4 ;
  wire \PWM0/sub1/c5 ;
  wire \PWM0/sub1/c6 ;
  wire \PWM0/sub1/c7 ;
  wire \PWM0/sub1/c8 ;
  wire \PWM0/sub1/c9 ;
  wire \PWM0/u14_sel_is_1_o ;
  wire \PWM1/RemaTxNum[0]_keep ;
  wire \PWM1/RemaTxNum[10]_keep ;
  wire \PWM1/RemaTxNum[11]_keep ;
  wire \PWM1/RemaTxNum[12]_keep ;
  wire \PWM1/RemaTxNum[13]_keep ;
  wire \PWM1/RemaTxNum[14]_keep ;
  wire \PWM1/RemaTxNum[15]_keep ;
  wire \PWM1/RemaTxNum[16]_keep ;
  wire \PWM1/RemaTxNum[17]_keep ;
  wire \PWM1/RemaTxNum[18]_keep ;
  wire \PWM1/RemaTxNum[19]_keep ;
  wire \PWM1/RemaTxNum[1]_keep ;
  wire \PWM1/RemaTxNum[20]_keep ;
  wire \PWM1/RemaTxNum[21]_keep ;
  wire \PWM1/RemaTxNum[22]_keep ;
  wire \PWM1/RemaTxNum[23]_keep ;
  wire \PWM1/RemaTxNum[2]_keep ;
  wire \PWM1/RemaTxNum[3]_keep ;
  wire \PWM1/RemaTxNum[4]_keep ;
  wire \PWM1/RemaTxNum[5]_keep ;
  wire \PWM1/RemaTxNum[6]_keep ;
  wire \PWM1/RemaTxNum[7]_keep ;
  wire \PWM1/RemaTxNum[8]_keep ;
  wire \PWM1/RemaTxNum[9]_keep ;
  wire \PWM1/dir_keep ;
  wire \PWM1/mux3_b0_sel_is_3_o ;
  wire \PWM1/n0_lutinv ;
  wire \PWM1/n1 ;
  wire \PWM1/n10 ;
  wire \PWM1/n11 ;
  wire \PWM1/n24 ;
  wire \PWM1/n25_neg_lutinv ;
  wire \PWM1/n32 ;
  wire \PWM1/pnumr[0]_keep ;
  wire \PWM1/pnumr[10]_keep ;
  wire \PWM1/pnumr[11]_keep ;
  wire \PWM1/pnumr[12]_keep ;
  wire \PWM1/pnumr[13]_keep ;
  wire \PWM1/pnumr[14]_keep ;
  wire \PWM1/pnumr[15]_keep ;
  wire \PWM1/pnumr[16]_keep ;
  wire \PWM1/pnumr[17]_keep ;
  wire \PWM1/pnumr[18]_keep ;
  wire \PWM1/pnumr[19]_keep ;
  wire \PWM1/pnumr[1]_keep ;
  wire \PWM1/pnumr[20]_keep ;
  wire \PWM1/pnumr[21]_keep ;
  wire \PWM1/pnumr[22]_keep ;
  wire \PWM1/pnumr[23]_keep ;
  wire \PWM1/pnumr[24]_keep ;
  wire \PWM1/pnumr[25]_keep ;
  wire \PWM1/pnumr[26]_keep ;
  wire \PWM1/pnumr[27]_keep ;
  wire \PWM1/pnumr[28]_keep ;
  wire \PWM1/pnumr[29]_keep ;
  wire \PWM1/pnumr[2]_keep ;
  wire \PWM1/pnumr[30]_keep ;
  wire \PWM1/pnumr[31]_keep ;
  wire \PWM1/pnumr[3]_keep ;
  wire \PWM1/pnumr[4]_keep ;
  wire \PWM1/pnumr[5]_keep ;
  wire \PWM1/pnumr[6]_keep ;
  wire \PWM1/pnumr[7]_keep ;
  wire \PWM1/pnumr[8]_keep ;
  wire \PWM1/pnumr[9]_keep ;
  wire \PWM1/pwm_keep ;
  wire \PWM1/stopreq ;  // src/OnePWM.v(14)
  wire \PWM1/stopreq_keep ;
  wire \PWM1/sub0/c0 ;
  wire \PWM1/sub0/c1 ;
  wire \PWM1/sub0/c10 ;
  wire \PWM1/sub0/c11 ;
  wire \PWM1/sub0/c12 ;
  wire \PWM1/sub0/c13 ;
  wire \PWM1/sub0/c14 ;
  wire \PWM1/sub0/c15 ;
  wire \PWM1/sub0/c16 ;
  wire \PWM1/sub0/c17 ;
  wire \PWM1/sub0/c18 ;
  wire \PWM1/sub0/c19 ;
  wire \PWM1/sub0/c2 ;
  wire \PWM1/sub0/c20 ;
  wire \PWM1/sub0/c21 ;
  wire \PWM1/sub0/c22 ;
  wire \PWM1/sub0/c23 ;
  wire \PWM1/sub0/c24 ;
  wire \PWM1/sub0/c25 ;
  wire \PWM1/sub0/c26 ;
  wire \PWM1/sub0/c3 ;
  wire \PWM1/sub0/c4 ;
  wire \PWM1/sub0/c5 ;
  wire \PWM1/sub0/c6 ;
  wire \PWM1/sub0/c7 ;
  wire \PWM1/sub0/c8 ;
  wire \PWM1/sub0/c9 ;
  wire \PWM1/sub1/c0 ;
  wire \PWM1/sub1/c1 ;
  wire \PWM1/sub1/c10 ;
  wire \PWM1/sub1/c11 ;
  wire \PWM1/sub1/c12 ;
  wire \PWM1/sub1/c13 ;
  wire \PWM1/sub1/c14 ;
  wire \PWM1/sub1/c15 ;
  wire \PWM1/sub1/c16 ;
  wire \PWM1/sub1/c17 ;
  wire \PWM1/sub1/c18 ;
  wire \PWM1/sub1/c19 ;
  wire \PWM1/sub1/c2 ;
  wire \PWM1/sub1/c20 ;
  wire \PWM1/sub1/c21 ;
  wire \PWM1/sub1/c22 ;
  wire \PWM1/sub1/c23 ;
  wire \PWM1/sub1/c3 ;
  wire \PWM1/sub1/c4 ;
  wire \PWM1/sub1/c5 ;
  wire \PWM1/sub1/c6 ;
  wire \PWM1/sub1/c7 ;
  wire \PWM1/sub1/c8 ;
  wire \PWM1/sub1/c9 ;
  wire \PWM1/u14_sel_is_1_o ;
  wire \PWM2/RemaTxNum[0]_keep ;
  wire \PWM2/RemaTxNum[10]_keep ;
  wire \PWM2/RemaTxNum[11]_keep ;
  wire \PWM2/RemaTxNum[12]_keep ;
  wire \PWM2/RemaTxNum[13]_keep ;
  wire \PWM2/RemaTxNum[14]_keep ;
  wire \PWM2/RemaTxNum[15]_keep ;
  wire \PWM2/RemaTxNum[16]_keep ;
  wire \PWM2/RemaTxNum[17]_keep ;
  wire \PWM2/RemaTxNum[18]_keep ;
  wire \PWM2/RemaTxNum[19]_keep ;
  wire \PWM2/RemaTxNum[1]_keep ;
  wire \PWM2/RemaTxNum[20]_keep ;
  wire \PWM2/RemaTxNum[21]_keep ;
  wire \PWM2/RemaTxNum[22]_keep ;
  wire \PWM2/RemaTxNum[23]_keep ;
  wire \PWM2/RemaTxNum[2]_keep ;
  wire \PWM2/RemaTxNum[3]_keep ;
  wire \PWM2/RemaTxNum[4]_keep ;
  wire \PWM2/RemaTxNum[5]_keep ;
  wire \PWM2/RemaTxNum[6]_keep ;
  wire \PWM2/RemaTxNum[7]_keep ;
  wire \PWM2/RemaTxNum[8]_keep ;
  wire \PWM2/RemaTxNum[9]_keep ;
  wire \PWM2/dir_keep ;
  wire \PWM2/mux3_b0_sel_is_3_o ;
  wire \PWM2/n0_lutinv ;
  wire \PWM2/n1 ;
  wire \PWM2/n10 ;
  wire \PWM2/n11 ;
  wire \PWM2/n24 ;
  wire \PWM2/n25_neg_lutinv ;
  wire \PWM2/n32 ;
  wire \PWM2/pnumr[0]_keep ;
  wire \PWM2/pnumr[10]_keep ;
  wire \PWM2/pnumr[11]_keep ;
  wire \PWM2/pnumr[12]_keep ;
  wire \PWM2/pnumr[13]_keep ;
  wire \PWM2/pnumr[14]_keep ;
  wire \PWM2/pnumr[15]_keep ;
  wire \PWM2/pnumr[16]_keep ;
  wire \PWM2/pnumr[17]_keep ;
  wire \PWM2/pnumr[18]_keep ;
  wire \PWM2/pnumr[19]_keep ;
  wire \PWM2/pnumr[1]_keep ;
  wire \PWM2/pnumr[20]_keep ;
  wire \PWM2/pnumr[21]_keep ;
  wire \PWM2/pnumr[22]_keep ;
  wire \PWM2/pnumr[23]_keep ;
  wire \PWM2/pnumr[24]_keep ;
  wire \PWM2/pnumr[25]_keep ;
  wire \PWM2/pnumr[26]_keep ;
  wire \PWM2/pnumr[27]_keep ;
  wire \PWM2/pnumr[28]_keep ;
  wire \PWM2/pnumr[29]_keep ;
  wire \PWM2/pnumr[2]_keep ;
  wire \PWM2/pnumr[30]_keep ;
  wire \PWM2/pnumr[31]_keep ;
  wire \PWM2/pnumr[3]_keep ;
  wire \PWM2/pnumr[4]_keep ;
  wire \PWM2/pnumr[5]_keep ;
  wire \PWM2/pnumr[6]_keep ;
  wire \PWM2/pnumr[7]_keep ;
  wire \PWM2/pnumr[8]_keep ;
  wire \PWM2/pnumr[9]_keep ;
  wire \PWM2/pwm_keep ;
  wire \PWM2/stopreq ;  // src/OnePWM.v(14)
  wire \PWM2/stopreq_keep ;
  wire \PWM2/sub0/c0 ;
  wire \PWM2/sub0/c1 ;
  wire \PWM2/sub0/c10 ;
  wire \PWM2/sub0/c11 ;
  wire \PWM2/sub0/c12 ;
  wire \PWM2/sub0/c13 ;
  wire \PWM2/sub0/c14 ;
  wire \PWM2/sub0/c15 ;
  wire \PWM2/sub0/c16 ;
  wire \PWM2/sub0/c17 ;
  wire \PWM2/sub0/c18 ;
  wire \PWM2/sub0/c19 ;
  wire \PWM2/sub0/c2 ;
  wire \PWM2/sub0/c20 ;
  wire \PWM2/sub0/c21 ;
  wire \PWM2/sub0/c22 ;
  wire \PWM2/sub0/c23 ;
  wire \PWM2/sub0/c24 ;
  wire \PWM2/sub0/c25 ;
  wire \PWM2/sub0/c26 ;
  wire \PWM2/sub0/c3 ;
  wire \PWM2/sub0/c4 ;
  wire \PWM2/sub0/c5 ;
  wire \PWM2/sub0/c6 ;
  wire \PWM2/sub0/c7 ;
  wire \PWM2/sub0/c8 ;
  wire \PWM2/sub0/c9 ;
  wire \PWM2/sub1/c0 ;
  wire \PWM2/sub1/c1 ;
  wire \PWM2/sub1/c10 ;
  wire \PWM2/sub1/c11 ;
  wire \PWM2/sub1/c12 ;
  wire \PWM2/sub1/c13 ;
  wire \PWM2/sub1/c14 ;
  wire \PWM2/sub1/c15 ;
  wire \PWM2/sub1/c16 ;
  wire \PWM2/sub1/c17 ;
  wire \PWM2/sub1/c18 ;
  wire \PWM2/sub1/c19 ;
  wire \PWM2/sub1/c2 ;
  wire \PWM2/sub1/c20 ;
  wire \PWM2/sub1/c21 ;
  wire \PWM2/sub1/c22 ;
  wire \PWM2/sub1/c23 ;
  wire \PWM2/sub1/c3 ;
  wire \PWM2/sub1/c4 ;
  wire \PWM2/sub1/c5 ;
  wire \PWM2/sub1/c6 ;
  wire \PWM2/sub1/c7 ;
  wire \PWM2/sub1/c8 ;
  wire \PWM2/sub1/c9 ;
  wire \PWM2/u14_sel_is_1_o ;
  wire \PWM3/RemaTxNum[0]_keep ;
  wire \PWM3/RemaTxNum[10]_keep ;
  wire \PWM3/RemaTxNum[11]_keep ;
  wire \PWM3/RemaTxNum[12]_keep ;
  wire \PWM3/RemaTxNum[13]_keep ;
  wire \PWM3/RemaTxNum[14]_keep ;
  wire \PWM3/RemaTxNum[15]_keep ;
  wire \PWM3/RemaTxNum[16]_keep ;
  wire \PWM3/RemaTxNum[17]_keep ;
  wire \PWM3/RemaTxNum[18]_keep ;
  wire \PWM3/RemaTxNum[19]_keep ;
  wire \PWM3/RemaTxNum[1]_keep ;
  wire \PWM3/RemaTxNum[20]_keep ;
  wire \PWM3/RemaTxNum[21]_keep ;
  wire \PWM3/RemaTxNum[22]_keep ;
  wire \PWM3/RemaTxNum[23]_keep ;
  wire \PWM3/RemaTxNum[2]_keep ;
  wire \PWM3/RemaTxNum[3]_keep ;
  wire \PWM3/RemaTxNum[4]_keep ;
  wire \PWM3/RemaTxNum[5]_keep ;
  wire \PWM3/RemaTxNum[6]_keep ;
  wire \PWM3/RemaTxNum[7]_keep ;
  wire \PWM3/RemaTxNum[8]_keep ;
  wire \PWM3/RemaTxNum[9]_keep ;
  wire \PWM3/dir_keep ;
  wire \PWM3/mux3_b0_sel_is_3_o ;
  wire \PWM3/n0_lutinv ;
  wire \PWM3/n1 ;
  wire \PWM3/n10 ;
  wire \PWM3/n11 ;
  wire \PWM3/n24 ;
  wire \PWM3/n25_neg_lutinv ;
  wire \PWM3/n32 ;
  wire \PWM3/pnumr[0]_keep ;
  wire \PWM3/pnumr[10]_keep ;
  wire \PWM3/pnumr[11]_keep ;
  wire \PWM3/pnumr[12]_keep ;
  wire \PWM3/pnumr[13]_keep ;
  wire \PWM3/pnumr[14]_keep ;
  wire \PWM3/pnumr[15]_keep ;
  wire \PWM3/pnumr[16]_keep ;
  wire \PWM3/pnumr[17]_keep ;
  wire \PWM3/pnumr[18]_keep ;
  wire \PWM3/pnumr[19]_keep ;
  wire \PWM3/pnumr[1]_keep ;
  wire \PWM3/pnumr[20]_keep ;
  wire \PWM3/pnumr[21]_keep ;
  wire \PWM3/pnumr[22]_keep ;
  wire \PWM3/pnumr[23]_keep ;
  wire \PWM3/pnumr[24]_keep ;
  wire \PWM3/pnumr[25]_keep ;
  wire \PWM3/pnumr[26]_keep ;
  wire \PWM3/pnumr[27]_keep ;
  wire \PWM3/pnumr[28]_keep ;
  wire \PWM3/pnumr[29]_keep ;
  wire \PWM3/pnumr[2]_keep ;
  wire \PWM3/pnumr[30]_keep ;
  wire \PWM3/pnumr[31]_keep ;
  wire \PWM3/pnumr[3]_keep ;
  wire \PWM3/pnumr[4]_keep ;
  wire \PWM3/pnumr[5]_keep ;
  wire \PWM3/pnumr[6]_keep ;
  wire \PWM3/pnumr[7]_keep ;
  wire \PWM3/pnumr[8]_keep ;
  wire \PWM3/pnumr[9]_keep ;
  wire \PWM3/pwm_keep ;
  wire \PWM3/stopreq ;  // src/OnePWM.v(14)
  wire \PWM3/stopreq_keep ;
  wire \PWM3/sub0/c0 ;
  wire \PWM3/sub0/c1 ;
  wire \PWM3/sub0/c10 ;
  wire \PWM3/sub0/c11 ;
  wire \PWM3/sub0/c12 ;
  wire \PWM3/sub0/c13 ;
  wire \PWM3/sub0/c14 ;
  wire \PWM3/sub0/c15 ;
  wire \PWM3/sub0/c16 ;
  wire \PWM3/sub0/c17 ;
  wire \PWM3/sub0/c18 ;
  wire \PWM3/sub0/c19 ;
  wire \PWM3/sub0/c2 ;
  wire \PWM3/sub0/c20 ;
  wire \PWM3/sub0/c21 ;
  wire \PWM3/sub0/c22 ;
  wire \PWM3/sub0/c23 ;
  wire \PWM3/sub0/c24 ;
  wire \PWM3/sub0/c25 ;
  wire \PWM3/sub0/c26 ;
  wire \PWM3/sub0/c3 ;
  wire \PWM3/sub0/c4 ;
  wire \PWM3/sub0/c5 ;
  wire \PWM3/sub0/c6 ;
  wire \PWM3/sub0/c7 ;
  wire \PWM3/sub0/c8 ;
  wire \PWM3/sub0/c9 ;
  wire \PWM3/sub1/c0 ;
  wire \PWM3/sub1/c1 ;
  wire \PWM3/sub1/c10 ;
  wire \PWM3/sub1/c11 ;
  wire \PWM3/sub1/c12 ;
  wire \PWM3/sub1/c13 ;
  wire \PWM3/sub1/c14 ;
  wire \PWM3/sub1/c15 ;
  wire \PWM3/sub1/c16 ;
  wire \PWM3/sub1/c17 ;
  wire \PWM3/sub1/c18 ;
  wire \PWM3/sub1/c19 ;
  wire \PWM3/sub1/c2 ;
  wire \PWM3/sub1/c20 ;
  wire \PWM3/sub1/c21 ;
  wire \PWM3/sub1/c22 ;
  wire \PWM3/sub1/c23 ;
  wire \PWM3/sub1/c3 ;
  wire \PWM3/sub1/c4 ;
  wire \PWM3/sub1/c5 ;
  wire \PWM3/sub1/c6 ;
  wire \PWM3/sub1/c7 ;
  wire \PWM3/sub1/c8 ;
  wire \PWM3/sub1/c9 ;
  wire \PWM3/u14_sel_is_1_o ;
  wire \PWM4/RemaTxNum[0]_keep ;
  wire \PWM4/RemaTxNum[10]_keep ;
  wire \PWM4/RemaTxNum[11]_keep ;
  wire \PWM4/RemaTxNum[12]_keep ;
  wire \PWM4/RemaTxNum[13]_keep ;
  wire \PWM4/RemaTxNum[14]_keep ;
  wire \PWM4/RemaTxNum[15]_keep ;
  wire \PWM4/RemaTxNum[16]_keep ;
  wire \PWM4/RemaTxNum[17]_keep ;
  wire \PWM4/RemaTxNum[18]_keep ;
  wire \PWM4/RemaTxNum[19]_keep ;
  wire \PWM4/RemaTxNum[1]_keep ;
  wire \PWM4/RemaTxNum[20]_keep ;
  wire \PWM4/RemaTxNum[21]_keep ;
  wire \PWM4/RemaTxNum[22]_keep ;
  wire \PWM4/RemaTxNum[23]_keep ;
  wire \PWM4/RemaTxNum[2]_keep ;
  wire \PWM4/RemaTxNum[3]_keep ;
  wire \PWM4/RemaTxNum[4]_keep ;
  wire \PWM4/RemaTxNum[5]_keep ;
  wire \PWM4/RemaTxNum[6]_keep ;
  wire \PWM4/RemaTxNum[7]_keep ;
  wire \PWM4/RemaTxNum[8]_keep ;
  wire \PWM4/RemaTxNum[9]_keep ;
  wire \PWM4/dir_keep ;
  wire \PWM4/mux3_b0_sel_is_3_o ;
  wire \PWM4/n0_lutinv ;
  wire \PWM4/n1 ;
  wire \PWM4/n10 ;
  wire \PWM4/n11 ;
  wire \PWM4/n24 ;
  wire \PWM4/n25_neg_lutinv ;
  wire \PWM4/n32 ;
  wire \PWM4/pnumr[0]_keep ;
  wire \PWM4/pnumr[10]_keep ;
  wire \PWM4/pnumr[11]_keep ;
  wire \PWM4/pnumr[12]_keep ;
  wire \PWM4/pnumr[13]_keep ;
  wire \PWM4/pnumr[14]_keep ;
  wire \PWM4/pnumr[15]_keep ;
  wire \PWM4/pnumr[16]_keep ;
  wire \PWM4/pnumr[17]_keep ;
  wire \PWM4/pnumr[18]_keep ;
  wire \PWM4/pnumr[19]_keep ;
  wire \PWM4/pnumr[1]_keep ;
  wire \PWM4/pnumr[20]_keep ;
  wire \PWM4/pnumr[21]_keep ;
  wire \PWM4/pnumr[22]_keep ;
  wire \PWM4/pnumr[23]_keep ;
  wire \PWM4/pnumr[24]_keep ;
  wire \PWM4/pnumr[25]_keep ;
  wire \PWM4/pnumr[26]_keep ;
  wire \PWM4/pnumr[27]_keep ;
  wire \PWM4/pnumr[28]_keep ;
  wire \PWM4/pnumr[29]_keep ;
  wire \PWM4/pnumr[2]_keep ;
  wire \PWM4/pnumr[30]_keep ;
  wire \PWM4/pnumr[31]_keep ;
  wire \PWM4/pnumr[3]_keep ;
  wire \PWM4/pnumr[4]_keep ;
  wire \PWM4/pnumr[5]_keep ;
  wire \PWM4/pnumr[6]_keep ;
  wire \PWM4/pnumr[7]_keep ;
  wire \PWM4/pnumr[8]_keep ;
  wire \PWM4/pnumr[9]_keep ;
  wire \PWM4/pwm_keep ;
  wire \PWM4/stopreq ;  // src/OnePWM.v(14)
  wire \PWM4/stopreq_keep ;
  wire \PWM4/sub0/c0 ;
  wire \PWM4/sub0/c1 ;
  wire \PWM4/sub0/c10 ;
  wire \PWM4/sub0/c11 ;
  wire \PWM4/sub0/c12 ;
  wire \PWM4/sub0/c13 ;
  wire \PWM4/sub0/c14 ;
  wire \PWM4/sub0/c15 ;
  wire \PWM4/sub0/c16 ;
  wire \PWM4/sub0/c17 ;
  wire \PWM4/sub0/c18 ;
  wire \PWM4/sub0/c19 ;
  wire \PWM4/sub0/c2 ;
  wire \PWM4/sub0/c20 ;
  wire \PWM4/sub0/c21 ;
  wire \PWM4/sub0/c22 ;
  wire \PWM4/sub0/c23 ;
  wire \PWM4/sub0/c24 ;
  wire \PWM4/sub0/c25 ;
  wire \PWM4/sub0/c26 ;
  wire \PWM4/sub0/c3 ;
  wire \PWM4/sub0/c4 ;
  wire \PWM4/sub0/c5 ;
  wire \PWM4/sub0/c6 ;
  wire \PWM4/sub0/c7 ;
  wire \PWM4/sub0/c8 ;
  wire \PWM4/sub0/c9 ;
  wire \PWM4/sub1/c0 ;
  wire \PWM4/sub1/c1 ;
  wire \PWM4/sub1/c10 ;
  wire \PWM4/sub1/c11 ;
  wire \PWM4/sub1/c12 ;
  wire \PWM4/sub1/c13 ;
  wire \PWM4/sub1/c14 ;
  wire \PWM4/sub1/c15 ;
  wire \PWM4/sub1/c16 ;
  wire \PWM4/sub1/c17 ;
  wire \PWM4/sub1/c18 ;
  wire \PWM4/sub1/c19 ;
  wire \PWM4/sub1/c2 ;
  wire \PWM4/sub1/c20 ;
  wire \PWM4/sub1/c21 ;
  wire \PWM4/sub1/c22 ;
  wire \PWM4/sub1/c23 ;
  wire \PWM4/sub1/c3 ;
  wire \PWM4/sub1/c4 ;
  wire \PWM4/sub1/c5 ;
  wire \PWM4/sub1/c6 ;
  wire \PWM4/sub1/c7 ;
  wire \PWM4/sub1/c8 ;
  wire \PWM4/sub1/c9 ;
  wire \PWM4/u14_sel_is_1_o ;
  wire \PWM5/RemaTxNum[0]_keep ;
  wire \PWM5/RemaTxNum[10]_keep ;
  wire \PWM5/RemaTxNum[11]_keep ;
  wire \PWM5/RemaTxNum[12]_keep ;
  wire \PWM5/RemaTxNum[13]_keep ;
  wire \PWM5/RemaTxNum[14]_keep ;
  wire \PWM5/RemaTxNum[15]_keep ;
  wire \PWM5/RemaTxNum[16]_keep ;
  wire \PWM5/RemaTxNum[17]_keep ;
  wire \PWM5/RemaTxNum[18]_keep ;
  wire \PWM5/RemaTxNum[19]_keep ;
  wire \PWM5/RemaTxNum[1]_keep ;
  wire \PWM5/RemaTxNum[20]_keep ;
  wire \PWM5/RemaTxNum[21]_keep ;
  wire \PWM5/RemaTxNum[22]_keep ;
  wire \PWM5/RemaTxNum[23]_keep ;
  wire \PWM5/RemaTxNum[2]_keep ;
  wire \PWM5/RemaTxNum[3]_keep ;
  wire \PWM5/RemaTxNum[4]_keep ;
  wire \PWM5/RemaTxNum[5]_keep ;
  wire \PWM5/RemaTxNum[6]_keep ;
  wire \PWM5/RemaTxNum[7]_keep ;
  wire \PWM5/RemaTxNum[8]_keep ;
  wire \PWM5/RemaTxNum[9]_keep ;
  wire \PWM5/dir_keep ;
  wire \PWM5/mux3_b0_sel_is_3_o ;
  wire \PWM5/n0_lutinv ;
  wire \PWM5/n1 ;
  wire \PWM5/n10 ;
  wire \PWM5/n11 ;
  wire \PWM5/n24 ;
  wire \PWM5/n25_neg_lutinv ;
  wire \PWM5/n32 ;
  wire \PWM5/pnumr[0]_keep ;
  wire \PWM5/pnumr[10]_keep ;
  wire \PWM5/pnumr[11]_keep ;
  wire \PWM5/pnumr[12]_keep ;
  wire \PWM5/pnumr[13]_keep ;
  wire \PWM5/pnumr[14]_keep ;
  wire \PWM5/pnumr[15]_keep ;
  wire \PWM5/pnumr[16]_keep ;
  wire \PWM5/pnumr[17]_keep ;
  wire \PWM5/pnumr[18]_keep ;
  wire \PWM5/pnumr[19]_keep ;
  wire \PWM5/pnumr[1]_keep ;
  wire \PWM5/pnumr[20]_keep ;
  wire \PWM5/pnumr[21]_keep ;
  wire \PWM5/pnumr[22]_keep ;
  wire \PWM5/pnumr[23]_keep ;
  wire \PWM5/pnumr[24]_keep ;
  wire \PWM5/pnumr[25]_keep ;
  wire \PWM5/pnumr[26]_keep ;
  wire \PWM5/pnumr[27]_keep ;
  wire \PWM5/pnumr[28]_keep ;
  wire \PWM5/pnumr[29]_keep ;
  wire \PWM5/pnumr[2]_keep ;
  wire \PWM5/pnumr[30]_keep ;
  wire \PWM5/pnumr[31]_keep ;
  wire \PWM5/pnumr[3]_keep ;
  wire \PWM5/pnumr[4]_keep ;
  wire \PWM5/pnumr[5]_keep ;
  wire \PWM5/pnumr[6]_keep ;
  wire \PWM5/pnumr[7]_keep ;
  wire \PWM5/pnumr[8]_keep ;
  wire \PWM5/pnumr[9]_keep ;
  wire \PWM5/pwm_keep ;
  wire \PWM5/stopreq ;  // src/OnePWM.v(14)
  wire \PWM5/stopreq_keep ;
  wire \PWM5/sub0/c0 ;
  wire \PWM5/sub0/c1 ;
  wire \PWM5/sub0/c10 ;
  wire \PWM5/sub0/c11 ;
  wire \PWM5/sub0/c12 ;
  wire \PWM5/sub0/c13 ;
  wire \PWM5/sub0/c14 ;
  wire \PWM5/sub0/c15 ;
  wire \PWM5/sub0/c16 ;
  wire \PWM5/sub0/c17 ;
  wire \PWM5/sub0/c18 ;
  wire \PWM5/sub0/c19 ;
  wire \PWM5/sub0/c2 ;
  wire \PWM5/sub0/c20 ;
  wire \PWM5/sub0/c21 ;
  wire \PWM5/sub0/c22 ;
  wire \PWM5/sub0/c23 ;
  wire \PWM5/sub0/c24 ;
  wire \PWM5/sub0/c25 ;
  wire \PWM5/sub0/c26 ;
  wire \PWM5/sub0/c3 ;
  wire \PWM5/sub0/c4 ;
  wire \PWM5/sub0/c5 ;
  wire \PWM5/sub0/c6 ;
  wire \PWM5/sub0/c7 ;
  wire \PWM5/sub0/c8 ;
  wire \PWM5/sub0/c9 ;
  wire \PWM5/sub1/c0 ;
  wire \PWM5/sub1/c1 ;
  wire \PWM5/sub1/c10 ;
  wire \PWM5/sub1/c11 ;
  wire \PWM5/sub1/c12 ;
  wire \PWM5/sub1/c13 ;
  wire \PWM5/sub1/c14 ;
  wire \PWM5/sub1/c15 ;
  wire \PWM5/sub1/c16 ;
  wire \PWM5/sub1/c17 ;
  wire \PWM5/sub1/c18 ;
  wire \PWM5/sub1/c19 ;
  wire \PWM5/sub1/c2 ;
  wire \PWM5/sub1/c20 ;
  wire \PWM5/sub1/c21 ;
  wire \PWM5/sub1/c22 ;
  wire \PWM5/sub1/c23 ;
  wire \PWM5/sub1/c3 ;
  wire \PWM5/sub1/c4 ;
  wire \PWM5/sub1/c5 ;
  wire \PWM5/sub1/c6 ;
  wire \PWM5/sub1/c7 ;
  wire \PWM5/sub1/c8 ;
  wire \PWM5/sub1/c9 ;
  wire \PWM5/u14_sel_is_1_o ;
  wire \PWM6/RemaTxNum[0]_keep ;
  wire \PWM6/RemaTxNum[10]_keep ;
  wire \PWM6/RemaTxNum[11]_keep ;
  wire \PWM6/RemaTxNum[12]_keep ;
  wire \PWM6/RemaTxNum[13]_keep ;
  wire \PWM6/RemaTxNum[14]_keep ;
  wire \PWM6/RemaTxNum[15]_keep ;
  wire \PWM6/RemaTxNum[16]_keep ;
  wire \PWM6/RemaTxNum[17]_keep ;
  wire \PWM6/RemaTxNum[18]_keep ;
  wire \PWM6/RemaTxNum[19]_keep ;
  wire \PWM6/RemaTxNum[1]_keep ;
  wire \PWM6/RemaTxNum[20]_keep ;
  wire \PWM6/RemaTxNum[21]_keep ;
  wire \PWM6/RemaTxNum[22]_keep ;
  wire \PWM6/RemaTxNum[23]_keep ;
  wire \PWM6/RemaTxNum[2]_keep ;
  wire \PWM6/RemaTxNum[3]_keep ;
  wire \PWM6/RemaTxNum[4]_keep ;
  wire \PWM6/RemaTxNum[5]_keep ;
  wire \PWM6/RemaTxNum[6]_keep ;
  wire \PWM6/RemaTxNum[7]_keep ;
  wire \PWM6/RemaTxNum[8]_keep ;
  wire \PWM6/RemaTxNum[9]_keep ;
  wire \PWM6/dir_keep ;
  wire \PWM6/mux3_b0_sel_is_3_o ;
  wire \PWM6/n0_lutinv ;
  wire \PWM6/n1 ;
  wire \PWM6/n10 ;
  wire \PWM6/n11 ;
  wire \PWM6/n18_lutinv ;
  wire \PWM6/n24 ;
  wire \PWM6/n25_neg_lutinv ;
  wire \PWM6/n32 ;
  wire \PWM6/pnumr[0]_keep ;
  wire \PWM6/pnumr[10]_keep ;
  wire \PWM6/pnumr[11]_keep ;
  wire \PWM6/pnumr[12]_keep ;
  wire \PWM6/pnumr[13]_keep ;
  wire \PWM6/pnumr[14]_keep ;
  wire \PWM6/pnumr[15]_keep ;
  wire \PWM6/pnumr[16]_keep ;
  wire \PWM6/pnumr[17]_keep ;
  wire \PWM6/pnumr[18]_keep ;
  wire \PWM6/pnumr[19]_keep ;
  wire \PWM6/pnumr[1]_keep ;
  wire \PWM6/pnumr[20]_keep ;
  wire \PWM6/pnumr[21]_keep ;
  wire \PWM6/pnumr[22]_keep ;
  wire \PWM6/pnumr[23]_keep ;
  wire \PWM6/pnumr[24]_keep ;
  wire \PWM6/pnumr[25]_keep ;
  wire \PWM6/pnumr[26]_keep ;
  wire \PWM6/pnumr[27]_keep ;
  wire \PWM6/pnumr[28]_keep ;
  wire \PWM6/pnumr[29]_keep ;
  wire \PWM6/pnumr[2]_keep ;
  wire \PWM6/pnumr[30]_keep ;
  wire \PWM6/pnumr[31]_keep ;
  wire \PWM6/pnumr[3]_keep ;
  wire \PWM6/pnumr[4]_keep ;
  wire \PWM6/pnumr[5]_keep ;
  wire \PWM6/pnumr[6]_keep ;
  wire \PWM6/pnumr[7]_keep ;
  wire \PWM6/pnumr[8]_keep ;
  wire \PWM6/pnumr[9]_keep ;
  wire \PWM6/pwm_keep ;
  wire \PWM6/stopreq ;  // src/OnePWM.v(14)
  wire \PWM6/stopreq_keep ;
  wire \PWM6/sub0/c0 ;
  wire \PWM6/sub0/c1 ;
  wire \PWM6/sub0/c10 ;
  wire \PWM6/sub0/c11 ;
  wire \PWM6/sub0/c12 ;
  wire \PWM6/sub0/c13 ;
  wire \PWM6/sub0/c14 ;
  wire \PWM6/sub0/c15 ;
  wire \PWM6/sub0/c16 ;
  wire \PWM6/sub0/c17 ;
  wire \PWM6/sub0/c18 ;
  wire \PWM6/sub0/c19 ;
  wire \PWM6/sub0/c2 ;
  wire \PWM6/sub0/c20 ;
  wire \PWM6/sub0/c21 ;
  wire \PWM6/sub0/c22 ;
  wire \PWM6/sub0/c23 ;
  wire \PWM6/sub0/c24 ;
  wire \PWM6/sub0/c25 ;
  wire \PWM6/sub0/c26 ;
  wire \PWM6/sub0/c3 ;
  wire \PWM6/sub0/c4 ;
  wire \PWM6/sub0/c5 ;
  wire \PWM6/sub0/c6 ;
  wire \PWM6/sub0/c7 ;
  wire \PWM6/sub0/c8 ;
  wire \PWM6/sub0/c9 ;
  wire \PWM6/sub1/c0 ;
  wire \PWM6/sub1/c1 ;
  wire \PWM6/sub1/c10 ;
  wire \PWM6/sub1/c11 ;
  wire \PWM6/sub1/c12 ;
  wire \PWM6/sub1/c13 ;
  wire \PWM6/sub1/c14 ;
  wire \PWM6/sub1/c15 ;
  wire \PWM6/sub1/c16 ;
  wire \PWM6/sub1/c17 ;
  wire \PWM6/sub1/c18 ;
  wire \PWM6/sub1/c19 ;
  wire \PWM6/sub1/c2 ;
  wire \PWM6/sub1/c20 ;
  wire \PWM6/sub1/c21 ;
  wire \PWM6/sub1/c22 ;
  wire \PWM6/sub1/c23 ;
  wire \PWM6/sub1/c3 ;
  wire \PWM6/sub1/c4 ;
  wire \PWM6/sub1/c5 ;
  wire \PWM6/sub1/c6 ;
  wire \PWM6/sub1/c7 ;
  wire \PWM6/sub1/c8 ;
  wire \PWM6/sub1/c9 ;
  wire \PWM6/u14_sel_is_1_o ;
  wire \PWM7/RemaTxNum[0]_keep ;
  wire \PWM7/RemaTxNum[10]_keep ;
  wire \PWM7/RemaTxNum[11]_keep ;
  wire \PWM7/RemaTxNum[12]_keep ;
  wire \PWM7/RemaTxNum[13]_keep ;
  wire \PWM7/RemaTxNum[14]_keep ;
  wire \PWM7/RemaTxNum[15]_keep ;
  wire \PWM7/RemaTxNum[16]_keep ;
  wire \PWM7/RemaTxNum[17]_keep ;
  wire \PWM7/RemaTxNum[18]_keep ;
  wire \PWM7/RemaTxNum[19]_keep ;
  wire \PWM7/RemaTxNum[1]_keep ;
  wire \PWM7/RemaTxNum[20]_keep ;
  wire \PWM7/RemaTxNum[21]_keep ;
  wire \PWM7/RemaTxNum[22]_keep ;
  wire \PWM7/RemaTxNum[23]_keep ;
  wire \PWM7/RemaTxNum[2]_keep ;
  wire \PWM7/RemaTxNum[3]_keep ;
  wire \PWM7/RemaTxNum[4]_keep ;
  wire \PWM7/RemaTxNum[5]_keep ;
  wire \PWM7/RemaTxNum[6]_keep ;
  wire \PWM7/RemaTxNum[7]_keep ;
  wire \PWM7/RemaTxNum[8]_keep ;
  wire \PWM7/RemaTxNum[9]_keep ;
  wire \PWM7/dir_keep ;
  wire \PWM7/mux3_b0_sel_is_3_o ;
  wire \PWM7/n0_lutinv ;
  wire \PWM7/n1 ;
  wire \PWM7/n10 ;
  wire \PWM7/n11 ;
  wire \PWM7/n24 ;
  wire \PWM7/n25_neg_lutinv ;
  wire \PWM7/n32 ;
  wire \PWM7/pnumr[0]_keep ;
  wire \PWM7/pnumr[10]_keep ;
  wire \PWM7/pnumr[11]_keep ;
  wire \PWM7/pnumr[12]_keep ;
  wire \PWM7/pnumr[13]_keep ;
  wire \PWM7/pnumr[14]_keep ;
  wire \PWM7/pnumr[15]_keep ;
  wire \PWM7/pnumr[16]_keep ;
  wire \PWM7/pnumr[17]_keep ;
  wire \PWM7/pnumr[18]_keep ;
  wire \PWM7/pnumr[19]_keep ;
  wire \PWM7/pnumr[1]_keep ;
  wire \PWM7/pnumr[20]_keep ;
  wire \PWM7/pnumr[21]_keep ;
  wire \PWM7/pnumr[22]_keep ;
  wire \PWM7/pnumr[23]_keep ;
  wire \PWM7/pnumr[24]_keep ;
  wire \PWM7/pnumr[25]_keep ;
  wire \PWM7/pnumr[26]_keep ;
  wire \PWM7/pnumr[27]_keep ;
  wire \PWM7/pnumr[28]_keep ;
  wire \PWM7/pnumr[29]_keep ;
  wire \PWM7/pnumr[2]_keep ;
  wire \PWM7/pnumr[30]_keep ;
  wire \PWM7/pnumr[31]_keep ;
  wire \PWM7/pnumr[3]_keep ;
  wire \PWM7/pnumr[4]_keep ;
  wire \PWM7/pnumr[5]_keep ;
  wire \PWM7/pnumr[6]_keep ;
  wire \PWM7/pnumr[7]_keep ;
  wire \PWM7/pnumr[8]_keep ;
  wire \PWM7/pnumr[9]_keep ;
  wire \PWM7/pwm_keep ;
  wire \PWM7/stopreq ;  // src/OnePWM.v(14)
  wire \PWM7/stopreq_keep ;
  wire \PWM7/sub0/c0 ;
  wire \PWM7/sub0/c1 ;
  wire \PWM7/sub0/c10 ;
  wire \PWM7/sub0/c11 ;
  wire \PWM7/sub0/c12 ;
  wire \PWM7/sub0/c13 ;
  wire \PWM7/sub0/c14 ;
  wire \PWM7/sub0/c15 ;
  wire \PWM7/sub0/c16 ;
  wire \PWM7/sub0/c17 ;
  wire \PWM7/sub0/c18 ;
  wire \PWM7/sub0/c19 ;
  wire \PWM7/sub0/c2 ;
  wire \PWM7/sub0/c20 ;
  wire \PWM7/sub0/c21 ;
  wire \PWM7/sub0/c22 ;
  wire \PWM7/sub0/c23 ;
  wire \PWM7/sub0/c24 ;
  wire \PWM7/sub0/c25 ;
  wire \PWM7/sub0/c26 ;
  wire \PWM7/sub0/c3 ;
  wire \PWM7/sub0/c4 ;
  wire \PWM7/sub0/c5 ;
  wire \PWM7/sub0/c6 ;
  wire \PWM7/sub0/c7 ;
  wire \PWM7/sub0/c8 ;
  wire \PWM7/sub0/c9 ;
  wire \PWM7/sub1/c0 ;
  wire \PWM7/sub1/c1 ;
  wire \PWM7/sub1/c10 ;
  wire \PWM7/sub1/c11 ;
  wire \PWM7/sub1/c12 ;
  wire \PWM7/sub1/c13 ;
  wire \PWM7/sub1/c14 ;
  wire \PWM7/sub1/c15 ;
  wire \PWM7/sub1/c16 ;
  wire \PWM7/sub1/c17 ;
  wire \PWM7/sub1/c18 ;
  wire \PWM7/sub1/c19 ;
  wire \PWM7/sub1/c2 ;
  wire \PWM7/sub1/c20 ;
  wire \PWM7/sub1/c21 ;
  wire \PWM7/sub1/c22 ;
  wire \PWM7/sub1/c23 ;
  wire \PWM7/sub1/c3 ;
  wire \PWM7/sub1/c4 ;
  wire \PWM7/sub1/c5 ;
  wire \PWM7/sub1/c6 ;
  wire \PWM7/sub1/c7 ;
  wire \PWM7/sub1/c8 ;
  wire \PWM7/sub1/c9 ;
  wire \PWM7/u14_sel_is_1_o ;
  wire \PWM8/RemaTxNum[0]_keep ;
  wire \PWM8/RemaTxNum[10]_keep ;
  wire \PWM8/RemaTxNum[11]_keep ;
  wire \PWM8/RemaTxNum[12]_keep ;
  wire \PWM8/RemaTxNum[13]_keep ;
  wire \PWM8/RemaTxNum[14]_keep ;
  wire \PWM8/RemaTxNum[15]_keep ;
  wire \PWM8/RemaTxNum[16]_keep ;
  wire \PWM8/RemaTxNum[17]_keep ;
  wire \PWM8/RemaTxNum[18]_keep ;
  wire \PWM8/RemaTxNum[19]_keep ;
  wire \PWM8/RemaTxNum[1]_keep ;
  wire \PWM8/RemaTxNum[20]_keep ;
  wire \PWM8/RemaTxNum[21]_keep ;
  wire \PWM8/RemaTxNum[22]_keep ;
  wire \PWM8/RemaTxNum[23]_keep ;
  wire \PWM8/RemaTxNum[2]_keep ;
  wire \PWM8/RemaTxNum[3]_keep ;
  wire \PWM8/RemaTxNum[4]_keep ;
  wire \PWM8/RemaTxNum[5]_keep ;
  wire \PWM8/RemaTxNum[6]_keep ;
  wire \PWM8/RemaTxNum[7]_keep ;
  wire \PWM8/RemaTxNum[8]_keep ;
  wire \PWM8/RemaTxNum[9]_keep ;
  wire \PWM8/dir_keep ;
  wire \PWM8/mux3_b0_sel_is_3_o ;
  wire \PWM8/n0_lutinv ;
  wire \PWM8/n1 ;
  wire \PWM8/n10 ;
  wire \PWM8/n11 ;
  wire \PWM8/n24 ;
  wire \PWM8/n25_neg_lutinv ;
  wire \PWM8/n32 ;
  wire \PWM8/pnumr[0]_keep ;
  wire \PWM8/pnumr[10]_keep ;
  wire \PWM8/pnumr[11]_keep ;
  wire \PWM8/pnumr[12]_keep ;
  wire \PWM8/pnumr[13]_keep ;
  wire \PWM8/pnumr[14]_keep ;
  wire \PWM8/pnumr[15]_keep ;
  wire \PWM8/pnumr[16]_keep ;
  wire \PWM8/pnumr[17]_keep ;
  wire \PWM8/pnumr[18]_keep ;
  wire \PWM8/pnumr[19]_keep ;
  wire \PWM8/pnumr[1]_keep ;
  wire \PWM8/pnumr[20]_keep ;
  wire \PWM8/pnumr[21]_keep ;
  wire \PWM8/pnumr[22]_keep ;
  wire \PWM8/pnumr[23]_keep ;
  wire \PWM8/pnumr[24]_keep ;
  wire \PWM8/pnumr[25]_keep ;
  wire \PWM8/pnumr[26]_keep ;
  wire \PWM8/pnumr[27]_keep ;
  wire \PWM8/pnumr[28]_keep ;
  wire \PWM8/pnumr[29]_keep ;
  wire \PWM8/pnumr[2]_keep ;
  wire \PWM8/pnumr[30]_keep ;
  wire \PWM8/pnumr[31]_keep ;
  wire \PWM8/pnumr[3]_keep ;
  wire \PWM8/pnumr[4]_keep ;
  wire \PWM8/pnumr[5]_keep ;
  wire \PWM8/pnumr[6]_keep ;
  wire \PWM8/pnumr[7]_keep ;
  wire \PWM8/pnumr[8]_keep ;
  wire \PWM8/pnumr[9]_keep ;
  wire \PWM8/pwm_keep ;
  wire \PWM8/stopreq ;  // src/OnePWM.v(14)
  wire \PWM8/stopreq_keep ;
  wire \PWM8/sub0/c0 ;
  wire \PWM8/sub0/c1 ;
  wire \PWM8/sub0/c10 ;
  wire \PWM8/sub0/c11 ;
  wire \PWM8/sub0/c12 ;
  wire \PWM8/sub0/c13 ;
  wire \PWM8/sub0/c14 ;
  wire \PWM8/sub0/c15 ;
  wire \PWM8/sub0/c16 ;
  wire \PWM8/sub0/c17 ;
  wire \PWM8/sub0/c18 ;
  wire \PWM8/sub0/c19 ;
  wire \PWM8/sub0/c2 ;
  wire \PWM8/sub0/c20 ;
  wire \PWM8/sub0/c21 ;
  wire \PWM8/sub0/c22 ;
  wire \PWM8/sub0/c23 ;
  wire \PWM8/sub0/c24 ;
  wire \PWM8/sub0/c25 ;
  wire \PWM8/sub0/c26 ;
  wire \PWM8/sub0/c3 ;
  wire \PWM8/sub0/c4 ;
  wire \PWM8/sub0/c5 ;
  wire \PWM8/sub0/c6 ;
  wire \PWM8/sub0/c7 ;
  wire \PWM8/sub0/c8 ;
  wire \PWM8/sub0/c9 ;
  wire \PWM8/sub1/c0 ;
  wire \PWM8/sub1/c1 ;
  wire \PWM8/sub1/c10 ;
  wire \PWM8/sub1/c11 ;
  wire \PWM8/sub1/c12 ;
  wire \PWM8/sub1/c13 ;
  wire \PWM8/sub1/c14 ;
  wire \PWM8/sub1/c15 ;
  wire \PWM8/sub1/c16 ;
  wire \PWM8/sub1/c17 ;
  wire \PWM8/sub1/c18 ;
  wire \PWM8/sub1/c19 ;
  wire \PWM8/sub1/c2 ;
  wire \PWM8/sub1/c20 ;
  wire \PWM8/sub1/c21 ;
  wire \PWM8/sub1/c22 ;
  wire \PWM8/sub1/c23 ;
  wire \PWM8/sub1/c3 ;
  wire \PWM8/sub1/c4 ;
  wire \PWM8/sub1/c5 ;
  wire \PWM8/sub1/c6 ;
  wire \PWM8/sub1/c7 ;
  wire \PWM8/sub1/c8 ;
  wire \PWM8/sub1/c9 ;
  wire \PWM8/u14_sel_is_1_o ;
  wire \PWM9/RemaTxNum[0]_keep ;
  wire \PWM9/RemaTxNum[10]_keep ;
  wire \PWM9/RemaTxNum[11]_keep ;
  wire \PWM9/RemaTxNum[12]_keep ;
  wire \PWM9/RemaTxNum[13]_keep ;
  wire \PWM9/RemaTxNum[14]_keep ;
  wire \PWM9/RemaTxNum[15]_keep ;
  wire \PWM9/RemaTxNum[16]_keep ;
  wire \PWM9/RemaTxNum[17]_keep ;
  wire \PWM9/RemaTxNum[18]_keep ;
  wire \PWM9/RemaTxNum[19]_keep ;
  wire \PWM9/RemaTxNum[1]_keep ;
  wire \PWM9/RemaTxNum[20]_keep ;
  wire \PWM9/RemaTxNum[21]_keep ;
  wire \PWM9/RemaTxNum[22]_keep ;
  wire \PWM9/RemaTxNum[23]_keep ;
  wire \PWM9/RemaTxNum[2]_keep ;
  wire \PWM9/RemaTxNum[3]_keep ;
  wire \PWM9/RemaTxNum[4]_keep ;
  wire \PWM9/RemaTxNum[5]_keep ;
  wire \PWM9/RemaTxNum[6]_keep ;
  wire \PWM9/RemaTxNum[7]_keep ;
  wire \PWM9/RemaTxNum[8]_keep ;
  wire \PWM9/RemaTxNum[9]_keep ;
  wire \PWM9/dir_keep ;
  wire \PWM9/mux3_b0_sel_is_3_o ;
  wire \PWM9/n0_lutinv ;
  wire \PWM9/n1 ;
  wire \PWM9/n10 ;
  wire \PWM9/n11 ;
  wire \PWM9/n24 ;
  wire \PWM9/n25_neg_lutinv ;
  wire \PWM9/n32 ;
  wire \PWM9/pnumr[0]_keep ;
  wire \PWM9/pnumr[10]_keep ;
  wire \PWM9/pnumr[11]_keep ;
  wire \PWM9/pnumr[12]_keep ;
  wire \PWM9/pnumr[13]_keep ;
  wire \PWM9/pnumr[14]_keep ;
  wire \PWM9/pnumr[15]_keep ;
  wire \PWM9/pnumr[16]_keep ;
  wire \PWM9/pnumr[17]_keep ;
  wire \PWM9/pnumr[18]_keep ;
  wire \PWM9/pnumr[19]_keep ;
  wire \PWM9/pnumr[1]_keep ;
  wire \PWM9/pnumr[20]_keep ;
  wire \PWM9/pnumr[21]_keep ;
  wire \PWM9/pnumr[22]_keep ;
  wire \PWM9/pnumr[23]_keep ;
  wire \PWM9/pnumr[24]_keep ;
  wire \PWM9/pnumr[25]_keep ;
  wire \PWM9/pnumr[26]_keep ;
  wire \PWM9/pnumr[27]_keep ;
  wire \PWM9/pnumr[28]_keep ;
  wire \PWM9/pnumr[29]_keep ;
  wire \PWM9/pnumr[2]_keep ;
  wire \PWM9/pnumr[30]_keep ;
  wire \PWM9/pnumr[31]_keep ;
  wire \PWM9/pnumr[3]_keep ;
  wire \PWM9/pnumr[4]_keep ;
  wire \PWM9/pnumr[5]_keep ;
  wire \PWM9/pnumr[6]_keep ;
  wire \PWM9/pnumr[7]_keep ;
  wire \PWM9/pnumr[8]_keep ;
  wire \PWM9/pnumr[9]_keep ;
  wire \PWM9/pwm_keep ;
  wire \PWM9/stopreq ;  // src/OnePWM.v(14)
  wire \PWM9/stopreq_keep ;
  wire \PWM9/sub0/c0 ;
  wire \PWM9/sub0/c1 ;
  wire \PWM9/sub0/c10 ;
  wire \PWM9/sub0/c11 ;
  wire \PWM9/sub0/c12 ;
  wire \PWM9/sub0/c13 ;
  wire \PWM9/sub0/c14 ;
  wire \PWM9/sub0/c15 ;
  wire \PWM9/sub0/c16 ;
  wire \PWM9/sub0/c17 ;
  wire \PWM9/sub0/c18 ;
  wire \PWM9/sub0/c19 ;
  wire \PWM9/sub0/c2 ;
  wire \PWM9/sub0/c20 ;
  wire \PWM9/sub0/c21 ;
  wire \PWM9/sub0/c22 ;
  wire \PWM9/sub0/c23 ;
  wire \PWM9/sub0/c24 ;
  wire \PWM9/sub0/c25 ;
  wire \PWM9/sub0/c26 ;
  wire \PWM9/sub0/c3 ;
  wire \PWM9/sub0/c4 ;
  wire \PWM9/sub0/c5 ;
  wire \PWM9/sub0/c6 ;
  wire \PWM9/sub0/c7 ;
  wire \PWM9/sub0/c8 ;
  wire \PWM9/sub0/c9 ;
  wire \PWM9/sub1/c0 ;
  wire \PWM9/sub1/c1 ;
  wire \PWM9/sub1/c10 ;
  wire \PWM9/sub1/c11 ;
  wire \PWM9/sub1/c12 ;
  wire \PWM9/sub1/c13 ;
  wire \PWM9/sub1/c14 ;
  wire \PWM9/sub1/c15 ;
  wire \PWM9/sub1/c16 ;
  wire \PWM9/sub1/c17 ;
  wire \PWM9/sub1/c18 ;
  wire \PWM9/sub1/c19 ;
  wire \PWM9/sub1/c2 ;
  wire \PWM9/sub1/c20 ;
  wire \PWM9/sub1/c21 ;
  wire \PWM9/sub1/c22 ;
  wire \PWM9/sub1/c23 ;
  wire \PWM9/sub1/c3 ;
  wire \PWM9/sub1/c4 ;
  wire \PWM9/sub1/c5 ;
  wire \PWM9/sub1/c6 ;
  wire \PWM9/sub1/c7 ;
  wire \PWM9/sub1/c8 ;
  wire \PWM9/sub1/c9 ;
  wire \PWM9/u14_sel_is_1_o ;
  wire \PWMA/RemaTxNum[0]_keep ;
  wire \PWMA/RemaTxNum[10]_keep ;
  wire \PWMA/RemaTxNum[11]_keep ;
  wire \PWMA/RemaTxNum[12]_keep ;
  wire \PWMA/RemaTxNum[13]_keep ;
  wire \PWMA/RemaTxNum[14]_keep ;
  wire \PWMA/RemaTxNum[15]_keep ;
  wire \PWMA/RemaTxNum[16]_keep ;
  wire \PWMA/RemaTxNum[17]_keep ;
  wire \PWMA/RemaTxNum[18]_keep ;
  wire \PWMA/RemaTxNum[19]_keep ;
  wire \PWMA/RemaTxNum[1]_keep ;
  wire \PWMA/RemaTxNum[20]_keep ;
  wire \PWMA/RemaTxNum[21]_keep ;
  wire \PWMA/RemaTxNum[22]_keep ;
  wire \PWMA/RemaTxNum[23]_keep ;
  wire \PWMA/RemaTxNum[2]_keep ;
  wire \PWMA/RemaTxNum[3]_keep ;
  wire \PWMA/RemaTxNum[4]_keep ;
  wire \PWMA/RemaTxNum[5]_keep ;
  wire \PWMA/RemaTxNum[6]_keep ;
  wire \PWMA/RemaTxNum[7]_keep ;
  wire \PWMA/RemaTxNum[8]_keep ;
  wire \PWMA/RemaTxNum[9]_keep ;
  wire \PWMA/dir_keep ;
  wire \PWMA/mux3_b0_sel_is_3_o ;
  wire \PWMA/n0_lutinv ;
  wire \PWMA/n1 ;
  wire \PWMA/n10 ;
  wire \PWMA/n11 ;
  wire \PWMA/n24 ;
  wire \PWMA/n25_neg_lutinv ;
  wire \PWMA/n32 ;
  wire \PWMA/pnumr[0]_keep ;
  wire \PWMA/pnumr[10]_keep ;
  wire \PWMA/pnumr[11]_keep ;
  wire \PWMA/pnumr[12]_keep ;
  wire \PWMA/pnumr[13]_keep ;
  wire \PWMA/pnumr[14]_keep ;
  wire \PWMA/pnumr[15]_keep ;
  wire \PWMA/pnumr[16]_keep ;
  wire \PWMA/pnumr[17]_keep ;
  wire \PWMA/pnumr[18]_keep ;
  wire \PWMA/pnumr[19]_keep ;
  wire \PWMA/pnumr[1]_keep ;
  wire \PWMA/pnumr[20]_keep ;
  wire \PWMA/pnumr[21]_keep ;
  wire \PWMA/pnumr[22]_keep ;
  wire \PWMA/pnumr[23]_keep ;
  wire \PWMA/pnumr[24]_keep ;
  wire \PWMA/pnumr[25]_keep ;
  wire \PWMA/pnumr[26]_keep ;
  wire \PWMA/pnumr[27]_keep ;
  wire \PWMA/pnumr[28]_keep ;
  wire \PWMA/pnumr[29]_keep ;
  wire \PWMA/pnumr[2]_keep ;
  wire \PWMA/pnumr[30]_keep ;
  wire \PWMA/pnumr[31]_keep ;
  wire \PWMA/pnumr[3]_keep ;
  wire \PWMA/pnumr[4]_keep ;
  wire \PWMA/pnumr[5]_keep ;
  wire \PWMA/pnumr[6]_keep ;
  wire \PWMA/pnumr[7]_keep ;
  wire \PWMA/pnumr[8]_keep ;
  wire \PWMA/pnumr[9]_keep ;
  wire \PWMA/pwm_keep ;
  wire \PWMA/stopreq ;  // src/OnePWM.v(14)
  wire \PWMA/stopreq_keep ;
  wire \PWMA/sub0/c0 ;
  wire \PWMA/sub0/c1 ;
  wire \PWMA/sub0/c10 ;
  wire \PWMA/sub0/c11 ;
  wire \PWMA/sub0/c12 ;
  wire \PWMA/sub0/c13 ;
  wire \PWMA/sub0/c14 ;
  wire \PWMA/sub0/c15 ;
  wire \PWMA/sub0/c16 ;
  wire \PWMA/sub0/c17 ;
  wire \PWMA/sub0/c18 ;
  wire \PWMA/sub0/c19 ;
  wire \PWMA/sub0/c2 ;
  wire \PWMA/sub0/c20 ;
  wire \PWMA/sub0/c21 ;
  wire \PWMA/sub0/c22 ;
  wire \PWMA/sub0/c23 ;
  wire \PWMA/sub0/c24 ;
  wire \PWMA/sub0/c25 ;
  wire \PWMA/sub0/c26 ;
  wire \PWMA/sub0/c3 ;
  wire \PWMA/sub0/c4 ;
  wire \PWMA/sub0/c5 ;
  wire \PWMA/sub0/c6 ;
  wire \PWMA/sub0/c7 ;
  wire \PWMA/sub0/c8 ;
  wire \PWMA/sub0/c9 ;
  wire \PWMA/sub1/c0 ;
  wire \PWMA/sub1/c1 ;
  wire \PWMA/sub1/c10 ;
  wire \PWMA/sub1/c11 ;
  wire \PWMA/sub1/c12 ;
  wire \PWMA/sub1/c13 ;
  wire \PWMA/sub1/c14 ;
  wire \PWMA/sub1/c15 ;
  wire \PWMA/sub1/c16 ;
  wire \PWMA/sub1/c17 ;
  wire \PWMA/sub1/c18 ;
  wire \PWMA/sub1/c19 ;
  wire \PWMA/sub1/c2 ;
  wire \PWMA/sub1/c20 ;
  wire \PWMA/sub1/c21 ;
  wire \PWMA/sub1/c22 ;
  wire \PWMA/sub1/c23 ;
  wire \PWMA/sub1/c3 ;
  wire \PWMA/sub1/c4 ;
  wire \PWMA/sub1/c5 ;
  wire \PWMA/sub1/c6 ;
  wire \PWMA/sub1/c7 ;
  wire \PWMA/sub1/c8 ;
  wire \PWMA/sub1/c9 ;
  wire \PWMA/u14_sel_is_1_o ;
  wire \PWMB/RemaTxNum[0]_keep ;
  wire \PWMB/RemaTxNum[10]_keep ;
  wire \PWMB/RemaTxNum[11]_keep ;
  wire \PWMB/RemaTxNum[12]_keep ;
  wire \PWMB/RemaTxNum[13]_keep ;
  wire \PWMB/RemaTxNum[14]_keep ;
  wire \PWMB/RemaTxNum[15]_keep ;
  wire \PWMB/RemaTxNum[16]_keep ;
  wire \PWMB/RemaTxNum[17]_keep ;
  wire \PWMB/RemaTxNum[18]_keep ;
  wire \PWMB/RemaTxNum[19]_keep ;
  wire \PWMB/RemaTxNum[1]_keep ;
  wire \PWMB/RemaTxNum[20]_keep ;
  wire \PWMB/RemaTxNum[21]_keep ;
  wire \PWMB/RemaTxNum[22]_keep ;
  wire \PWMB/RemaTxNum[23]_keep ;
  wire \PWMB/RemaTxNum[2]_keep ;
  wire \PWMB/RemaTxNum[3]_keep ;
  wire \PWMB/RemaTxNum[4]_keep ;
  wire \PWMB/RemaTxNum[5]_keep ;
  wire \PWMB/RemaTxNum[6]_keep ;
  wire \PWMB/RemaTxNum[7]_keep ;
  wire \PWMB/RemaTxNum[8]_keep ;
  wire \PWMB/RemaTxNum[9]_keep ;
  wire \PWMB/dir_keep ;
  wire \PWMB/mux3_b0_sel_is_3_o ;
  wire \PWMB/n0_lutinv ;
  wire \PWMB/n1 ;
  wire \PWMB/n10 ;
  wire \PWMB/n11 ;
  wire \PWMB/n24 ;
  wire \PWMB/n25_neg_lutinv ;
  wire \PWMB/n32 ;
  wire \PWMB/pnumr[0]_keep ;
  wire \PWMB/pnumr[10]_keep ;
  wire \PWMB/pnumr[11]_keep ;
  wire \PWMB/pnumr[12]_keep ;
  wire \PWMB/pnumr[13]_keep ;
  wire \PWMB/pnumr[14]_keep ;
  wire \PWMB/pnumr[15]_keep ;
  wire \PWMB/pnumr[16]_keep ;
  wire \PWMB/pnumr[17]_keep ;
  wire \PWMB/pnumr[18]_keep ;
  wire \PWMB/pnumr[19]_keep ;
  wire \PWMB/pnumr[1]_keep ;
  wire \PWMB/pnumr[20]_keep ;
  wire \PWMB/pnumr[21]_keep ;
  wire \PWMB/pnumr[22]_keep ;
  wire \PWMB/pnumr[23]_keep ;
  wire \PWMB/pnumr[24]_keep ;
  wire \PWMB/pnumr[25]_keep ;
  wire \PWMB/pnumr[26]_keep ;
  wire \PWMB/pnumr[27]_keep ;
  wire \PWMB/pnumr[28]_keep ;
  wire \PWMB/pnumr[29]_keep ;
  wire \PWMB/pnumr[2]_keep ;
  wire \PWMB/pnumr[30]_keep ;
  wire \PWMB/pnumr[31]_keep ;
  wire \PWMB/pnumr[3]_keep ;
  wire \PWMB/pnumr[4]_keep ;
  wire \PWMB/pnumr[5]_keep ;
  wire \PWMB/pnumr[6]_keep ;
  wire \PWMB/pnumr[7]_keep ;
  wire \PWMB/pnumr[8]_keep ;
  wire \PWMB/pnumr[9]_keep ;
  wire \PWMB/pwm_keep ;
  wire \PWMB/stopreq ;  // src/OnePWM.v(14)
  wire \PWMB/stopreq_keep ;
  wire \PWMB/sub0/c0 ;
  wire \PWMB/sub0/c1 ;
  wire \PWMB/sub0/c10 ;
  wire \PWMB/sub0/c11 ;
  wire \PWMB/sub0/c12 ;
  wire \PWMB/sub0/c13 ;
  wire \PWMB/sub0/c14 ;
  wire \PWMB/sub0/c15 ;
  wire \PWMB/sub0/c16 ;
  wire \PWMB/sub0/c17 ;
  wire \PWMB/sub0/c18 ;
  wire \PWMB/sub0/c19 ;
  wire \PWMB/sub0/c2 ;
  wire \PWMB/sub0/c20 ;
  wire \PWMB/sub0/c21 ;
  wire \PWMB/sub0/c22 ;
  wire \PWMB/sub0/c23 ;
  wire \PWMB/sub0/c24 ;
  wire \PWMB/sub0/c25 ;
  wire \PWMB/sub0/c26 ;
  wire \PWMB/sub0/c3 ;
  wire \PWMB/sub0/c4 ;
  wire \PWMB/sub0/c5 ;
  wire \PWMB/sub0/c6 ;
  wire \PWMB/sub0/c7 ;
  wire \PWMB/sub0/c8 ;
  wire \PWMB/sub0/c9 ;
  wire \PWMB/sub1/c0 ;
  wire \PWMB/sub1/c1 ;
  wire \PWMB/sub1/c10 ;
  wire \PWMB/sub1/c11 ;
  wire \PWMB/sub1/c12 ;
  wire \PWMB/sub1/c13 ;
  wire \PWMB/sub1/c14 ;
  wire \PWMB/sub1/c15 ;
  wire \PWMB/sub1/c16 ;
  wire \PWMB/sub1/c17 ;
  wire \PWMB/sub1/c18 ;
  wire \PWMB/sub1/c19 ;
  wire \PWMB/sub1/c2 ;
  wire \PWMB/sub1/c20 ;
  wire \PWMB/sub1/c21 ;
  wire \PWMB/sub1/c22 ;
  wire \PWMB/sub1/c23 ;
  wire \PWMB/sub1/c3 ;
  wire \PWMB/sub1/c4 ;
  wire \PWMB/sub1/c5 ;
  wire \PWMB/sub1/c6 ;
  wire \PWMB/sub1/c7 ;
  wire \PWMB/sub1/c8 ;
  wire \PWMB/sub1/c9 ;
  wire \PWMB/u14_sel_is_1_o ;
  wire \PWMC/RemaTxNum[0]_keep ;
  wire \PWMC/RemaTxNum[10]_keep ;
  wire \PWMC/RemaTxNum[11]_keep ;
  wire \PWMC/RemaTxNum[12]_keep ;
  wire \PWMC/RemaTxNum[13]_keep ;
  wire \PWMC/RemaTxNum[14]_keep ;
  wire \PWMC/RemaTxNum[15]_keep ;
  wire \PWMC/RemaTxNum[16]_keep ;
  wire \PWMC/RemaTxNum[17]_keep ;
  wire \PWMC/RemaTxNum[18]_keep ;
  wire \PWMC/RemaTxNum[19]_keep ;
  wire \PWMC/RemaTxNum[1]_keep ;
  wire \PWMC/RemaTxNum[20]_keep ;
  wire \PWMC/RemaTxNum[21]_keep ;
  wire \PWMC/RemaTxNum[22]_keep ;
  wire \PWMC/RemaTxNum[23]_keep ;
  wire \PWMC/RemaTxNum[2]_keep ;
  wire \PWMC/RemaTxNum[3]_keep ;
  wire \PWMC/RemaTxNum[4]_keep ;
  wire \PWMC/RemaTxNum[5]_keep ;
  wire \PWMC/RemaTxNum[6]_keep ;
  wire \PWMC/RemaTxNum[7]_keep ;
  wire \PWMC/RemaTxNum[8]_keep ;
  wire \PWMC/RemaTxNum[9]_keep ;
  wire \PWMC/dir_keep ;
  wire \PWMC/mux3_b0_sel_is_3_o ;
  wire \PWMC/n0_lutinv ;
  wire \PWMC/n1 ;
  wire \PWMC/n10 ;
  wire \PWMC/n11 ;
  wire \PWMC/n24 ;
  wire \PWMC/n25_neg_lutinv ;
  wire \PWMC/n32 ;
  wire \PWMC/pnumr[0]_keep ;
  wire \PWMC/pnumr[10]_keep ;
  wire \PWMC/pnumr[11]_keep ;
  wire \PWMC/pnumr[12]_keep ;
  wire \PWMC/pnumr[13]_keep ;
  wire \PWMC/pnumr[14]_keep ;
  wire \PWMC/pnumr[15]_keep ;
  wire \PWMC/pnumr[16]_keep ;
  wire \PWMC/pnumr[17]_keep ;
  wire \PWMC/pnumr[18]_keep ;
  wire \PWMC/pnumr[19]_keep ;
  wire \PWMC/pnumr[1]_keep ;
  wire \PWMC/pnumr[20]_keep ;
  wire \PWMC/pnumr[21]_keep ;
  wire \PWMC/pnumr[22]_keep ;
  wire \PWMC/pnumr[23]_keep ;
  wire \PWMC/pnumr[24]_keep ;
  wire \PWMC/pnumr[25]_keep ;
  wire \PWMC/pnumr[26]_keep ;
  wire \PWMC/pnumr[27]_keep ;
  wire \PWMC/pnumr[28]_keep ;
  wire \PWMC/pnumr[29]_keep ;
  wire \PWMC/pnumr[2]_keep ;
  wire \PWMC/pnumr[30]_keep ;
  wire \PWMC/pnumr[31]_keep ;
  wire \PWMC/pnumr[3]_keep ;
  wire \PWMC/pnumr[4]_keep ;
  wire \PWMC/pnumr[5]_keep ;
  wire \PWMC/pnumr[6]_keep ;
  wire \PWMC/pnumr[7]_keep ;
  wire \PWMC/pnumr[8]_keep ;
  wire \PWMC/pnumr[9]_keep ;
  wire \PWMC/pwm_keep ;
  wire \PWMC/stopreq ;  // src/OnePWM.v(14)
  wire \PWMC/stopreq_keep ;
  wire \PWMC/sub0/c0 ;
  wire \PWMC/sub0/c1 ;
  wire \PWMC/sub0/c10 ;
  wire \PWMC/sub0/c11 ;
  wire \PWMC/sub0/c12 ;
  wire \PWMC/sub0/c13 ;
  wire \PWMC/sub0/c14 ;
  wire \PWMC/sub0/c15 ;
  wire \PWMC/sub0/c16 ;
  wire \PWMC/sub0/c17 ;
  wire \PWMC/sub0/c18 ;
  wire \PWMC/sub0/c19 ;
  wire \PWMC/sub0/c2 ;
  wire \PWMC/sub0/c20 ;
  wire \PWMC/sub0/c21 ;
  wire \PWMC/sub0/c22 ;
  wire \PWMC/sub0/c23 ;
  wire \PWMC/sub0/c24 ;
  wire \PWMC/sub0/c25 ;
  wire \PWMC/sub0/c26 ;
  wire \PWMC/sub0/c3 ;
  wire \PWMC/sub0/c4 ;
  wire \PWMC/sub0/c5 ;
  wire \PWMC/sub0/c6 ;
  wire \PWMC/sub0/c7 ;
  wire \PWMC/sub0/c8 ;
  wire \PWMC/sub0/c9 ;
  wire \PWMC/sub1/c0 ;
  wire \PWMC/sub1/c1 ;
  wire \PWMC/sub1/c10 ;
  wire \PWMC/sub1/c11 ;
  wire \PWMC/sub1/c12 ;
  wire \PWMC/sub1/c13 ;
  wire \PWMC/sub1/c14 ;
  wire \PWMC/sub1/c15 ;
  wire \PWMC/sub1/c16 ;
  wire \PWMC/sub1/c17 ;
  wire \PWMC/sub1/c18 ;
  wire \PWMC/sub1/c19 ;
  wire \PWMC/sub1/c2 ;
  wire \PWMC/sub1/c20 ;
  wire \PWMC/sub1/c21 ;
  wire \PWMC/sub1/c22 ;
  wire \PWMC/sub1/c23 ;
  wire \PWMC/sub1/c3 ;
  wire \PWMC/sub1/c4 ;
  wire \PWMC/sub1/c5 ;
  wire \PWMC/sub1/c6 ;
  wire \PWMC/sub1/c7 ;
  wire \PWMC/sub1/c8 ;
  wire \PWMC/sub1/c9 ;
  wire \PWMC/u14_sel_is_1_o ;
  wire \PWMD/RemaTxNum[0]_keep ;
  wire \PWMD/RemaTxNum[10]_keep ;
  wire \PWMD/RemaTxNum[11]_keep ;
  wire \PWMD/RemaTxNum[12]_keep ;
  wire \PWMD/RemaTxNum[13]_keep ;
  wire \PWMD/RemaTxNum[14]_keep ;
  wire \PWMD/RemaTxNum[15]_keep ;
  wire \PWMD/RemaTxNum[16]_keep ;
  wire \PWMD/RemaTxNum[17]_keep ;
  wire \PWMD/RemaTxNum[18]_keep ;
  wire \PWMD/RemaTxNum[19]_keep ;
  wire \PWMD/RemaTxNum[1]_keep ;
  wire \PWMD/RemaTxNum[20]_keep ;
  wire \PWMD/RemaTxNum[21]_keep ;
  wire \PWMD/RemaTxNum[22]_keep ;
  wire \PWMD/RemaTxNum[23]_keep ;
  wire \PWMD/RemaTxNum[2]_keep ;
  wire \PWMD/RemaTxNum[3]_keep ;
  wire \PWMD/RemaTxNum[4]_keep ;
  wire \PWMD/RemaTxNum[5]_keep ;
  wire \PWMD/RemaTxNum[6]_keep ;
  wire \PWMD/RemaTxNum[7]_keep ;
  wire \PWMD/RemaTxNum[8]_keep ;
  wire \PWMD/RemaTxNum[9]_keep ;
  wire \PWMD/dir_keep ;
  wire \PWMD/mux3_b0_sel_is_3_o ;
  wire \PWMD/n0_lutinv ;
  wire \PWMD/n1 ;
  wire \PWMD/n10 ;
  wire \PWMD/n11 ;
  wire \PWMD/n24 ;
  wire \PWMD/n25_neg_lutinv ;
  wire \PWMD/n32 ;
  wire \PWMD/pnumr[0]_keep ;
  wire \PWMD/pnumr[10]_keep ;
  wire \PWMD/pnumr[11]_keep ;
  wire \PWMD/pnumr[12]_keep ;
  wire \PWMD/pnumr[13]_keep ;
  wire \PWMD/pnumr[14]_keep ;
  wire \PWMD/pnumr[15]_keep ;
  wire \PWMD/pnumr[16]_keep ;
  wire \PWMD/pnumr[17]_keep ;
  wire \PWMD/pnumr[18]_keep ;
  wire \PWMD/pnumr[19]_keep ;
  wire \PWMD/pnumr[1]_keep ;
  wire \PWMD/pnumr[20]_keep ;
  wire \PWMD/pnumr[21]_keep ;
  wire \PWMD/pnumr[22]_keep ;
  wire \PWMD/pnumr[23]_keep ;
  wire \PWMD/pnumr[24]_keep ;
  wire \PWMD/pnumr[25]_keep ;
  wire \PWMD/pnumr[26]_keep ;
  wire \PWMD/pnumr[27]_keep ;
  wire \PWMD/pnumr[28]_keep ;
  wire \PWMD/pnumr[29]_keep ;
  wire \PWMD/pnumr[2]_keep ;
  wire \PWMD/pnumr[30]_keep ;
  wire \PWMD/pnumr[31]_keep ;
  wire \PWMD/pnumr[3]_keep ;
  wire \PWMD/pnumr[4]_keep ;
  wire \PWMD/pnumr[5]_keep ;
  wire \PWMD/pnumr[6]_keep ;
  wire \PWMD/pnumr[7]_keep ;
  wire \PWMD/pnumr[8]_keep ;
  wire \PWMD/pnumr[9]_keep ;
  wire \PWMD/pwm_keep ;
  wire \PWMD/stopreq ;  // src/OnePWM.v(14)
  wire \PWMD/stopreq_keep ;
  wire \PWMD/sub0/c0 ;
  wire \PWMD/sub0/c1 ;
  wire \PWMD/sub0/c10 ;
  wire \PWMD/sub0/c11 ;
  wire \PWMD/sub0/c12 ;
  wire \PWMD/sub0/c13 ;
  wire \PWMD/sub0/c14 ;
  wire \PWMD/sub0/c15 ;
  wire \PWMD/sub0/c16 ;
  wire \PWMD/sub0/c17 ;
  wire \PWMD/sub0/c18 ;
  wire \PWMD/sub0/c19 ;
  wire \PWMD/sub0/c2 ;
  wire \PWMD/sub0/c20 ;
  wire \PWMD/sub0/c21 ;
  wire \PWMD/sub0/c22 ;
  wire \PWMD/sub0/c23 ;
  wire \PWMD/sub0/c24 ;
  wire \PWMD/sub0/c25 ;
  wire \PWMD/sub0/c26 ;
  wire \PWMD/sub0/c3 ;
  wire \PWMD/sub0/c4 ;
  wire \PWMD/sub0/c5 ;
  wire \PWMD/sub0/c6 ;
  wire \PWMD/sub0/c7 ;
  wire \PWMD/sub0/c8 ;
  wire \PWMD/sub0/c9 ;
  wire \PWMD/sub1/c0 ;
  wire \PWMD/sub1/c1 ;
  wire \PWMD/sub1/c10 ;
  wire \PWMD/sub1/c11 ;
  wire \PWMD/sub1/c12 ;
  wire \PWMD/sub1/c13 ;
  wire \PWMD/sub1/c14 ;
  wire \PWMD/sub1/c15 ;
  wire \PWMD/sub1/c16 ;
  wire \PWMD/sub1/c17 ;
  wire \PWMD/sub1/c18 ;
  wire \PWMD/sub1/c19 ;
  wire \PWMD/sub1/c2 ;
  wire \PWMD/sub1/c20 ;
  wire \PWMD/sub1/c21 ;
  wire \PWMD/sub1/c22 ;
  wire \PWMD/sub1/c23 ;
  wire \PWMD/sub1/c3 ;
  wire \PWMD/sub1/c4 ;
  wire \PWMD/sub1/c5 ;
  wire \PWMD/sub1/c6 ;
  wire \PWMD/sub1/c7 ;
  wire \PWMD/sub1/c8 ;
  wire \PWMD/sub1/c9 ;
  wire \PWMD/u14_sel_is_1_o ;
  wire \PWME/RemaTxNum[0]_keep ;
  wire \PWME/RemaTxNum[10]_keep ;
  wire \PWME/RemaTxNum[11]_keep ;
  wire \PWME/RemaTxNum[12]_keep ;
  wire \PWME/RemaTxNum[13]_keep ;
  wire \PWME/RemaTxNum[14]_keep ;
  wire \PWME/RemaTxNum[15]_keep ;
  wire \PWME/RemaTxNum[16]_keep ;
  wire \PWME/RemaTxNum[17]_keep ;
  wire \PWME/RemaTxNum[18]_keep ;
  wire \PWME/RemaTxNum[19]_keep ;
  wire \PWME/RemaTxNum[1]_keep ;
  wire \PWME/RemaTxNum[20]_keep ;
  wire \PWME/RemaTxNum[21]_keep ;
  wire \PWME/RemaTxNum[22]_keep ;
  wire \PWME/RemaTxNum[23]_keep ;
  wire \PWME/RemaTxNum[2]_keep ;
  wire \PWME/RemaTxNum[3]_keep ;
  wire \PWME/RemaTxNum[4]_keep ;
  wire \PWME/RemaTxNum[5]_keep ;
  wire \PWME/RemaTxNum[6]_keep ;
  wire \PWME/RemaTxNum[7]_keep ;
  wire \PWME/RemaTxNum[8]_keep ;
  wire \PWME/RemaTxNum[9]_keep ;
  wire \PWME/dir_keep ;
  wire \PWME/mux3_b0_sel_is_3_o ;
  wire \PWME/n0_lutinv ;
  wire \PWME/n1 ;
  wire \PWME/n10 ;
  wire \PWME/n11 ;
  wire \PWME/n24 ;
  wire \PWME/n25_neg_lutinv ;
  wire \PWME/n32 ;
  wire \PWME/pnumr[0]_keep ;
  wire \PWME/pnumr[10]_keep ;
  wire \PWME/pnumr[11]_keep ;
  wire \PWME/pnumr[12]_keep ;
  wire \PWME/pnumr[13]_keep ;
  wire \PWME/pnumr[14]_keep ;
  wire \PWME/pnumr[15]_keep ;
  wire \PWME/pnumr[16]_keep ;
  wire \PWME/pnumr[17]_keep ;
  wire \PWME/pnumr[18]_keep ;
  wire \PWME/pnumr[19]_keep ;
  wire \PWME/pnumr[1]_keep ;
  wire \PWME/pnumr[20]_keep ;
  wire \PWME/pnumr[21]_keep ;
  wire \PWME/pnumr[22]_keep ;
  wire \PWME/pnumr[23]_keep ;
  wire \PWME/pnumr[24]_keep ;
  wire \PWME/pnumr[25]_keep ;
  wire \PWME/pnumr[26]_keep ;
  wire \PWME/pnumr[27]_keep ;
  wire \PWME/pnumr[28]_keep ;
  wire \PWME/pnumr[29]_keep ;
  wire \PWME/pnumr[2]_keep ;
  wire \PWME/pnumr[30]_keep ;
  wire \PWME/pnumr[31]_keep ;
  wire \PWME/pnumr[3]_keep ;
  wire \PWME/pnumr[4]_keep ;
  wire \PWME/pnumr[5]_keep ;
  wire \PWME/pnumr[6]_keep ;
  wire \PWME/pnumr[7]_keep ;
  wire \PWME/pnumr[8]_keep ;
  wire \PWME/pnumr[9]_keep ;
  wire \PWME/pwm_keep ;
  wire \PWME/stopreq ;  // src/OnePWM.v(14)
  wire \PWME/stopreq_keep ;
  wire \PWME/sub0/c0 ;
  wire \PWME/sub0/c1 ;
  wire \PWME/sub0/c10 ;
  wire \PWME/sub0/c11 ;
  wire \PWME/sub0/c12 ;
  wire \PWME/sub0/c13 ;
  wire \PWME/sub0/c14 ;
  wire \PWME/sub0/c15 ;
  wire \PWME/sub0/c16 ;
  wire \PWME/sub0/c17 ;
  wire \PWME/sub0/c18 ;
  wire \PWME/sub0/c19 ;
  wire \PWME/sub0/c2 ;
  wire \PWME/sub0/c20 ;
  wire \PWME/sub0/c21 ;
  wire \PWME/sub0/c22 ;
  wire \PWME/sub0/c23 ;
  wire \PWME/sub0/c24 ;
  wire \PWME/sub0/c25 ;
  wire \PWME/sub0/c26 ;
  wire \PWME/sub0/c3 ;
  wire \PWME/sub0/c4 ;
  wire \PWME/sub0/c5 ;
  wire \PWME/sub0/c6 ;
  wire \PWME/sub0/c7 ;
  wire \PWME/sub0/c8 ;
  wire \PWME/sub0/c9 ;
  wire \PWME/sub1/c0 ;
  wire \PWME/sub1/c1 ;
  wire \PWME/sub1/c10 ;
  wire \PWME/sub1/c11 ;
  wire \PWME/sub1/c12 ;
  wire \PWME/sub1/c13 ;
  wire \PWME/sub1/c14 ;
  wire \PWME/sub1/c15 ;
  wire \PWME/sub1/c16 ;
  wire \PWME/sub1/c17 ;
  wire \PWME/sub1/c18 ;
  wire \PWME/sub1/c19 ;
  wire \PWME/sub1/c2 ;
  wire \PWME/sub1/c20 ;
  wire \PWME/sub1/c21 ;
  wire \PWME/sub1/c22 ;
  wire \PWME/sub1/c23 ;
  wire \PWME/sub1/c3 ;
  wire \PWME/sub1/c4 ;
  wire \PWME/sub1/c5 ;
  wire \PWME/sub1/c6 ;
  wire \PWME/sub1/c7 ;
  wire \PWME/sub1/c8 ;
  wire \PWME/sub1/c9 ;
  wire \PWME/u14_sel_is_1_o ;
  wire \PWMF/RemaTxNum[0]_keep ;
  wire \PWMF/RemaTxNum[10]_keep ;
  wire \PWMF/RemaTxNum[11]_keep ;
  wire \PWMF/RemaTxNum[12]_keep ;
  wire \PWMF/RemaTxNum[13]_keep ;
  wire \PWMF/RemaTxNum[14]_keep ;
  wire \PWMF/RemaTxNum[15]_keep ;
  wire \PWMF/RemaTxNum[16]_keep ;
  wire \PWMF/RemaTxNum[17]_keep ;
  wire \PWMF/RemaTxNum[18]_keep ;
  wire \PWMF/RemaTxNum[19]_keep ;
  wire \PWMF/RemaTxNum[1]_keep ;
  wire \PWMF/RemaTxNum[20]_keep ;
  wire \PWMF/RemaTxNum[21]_keep ;
  wire \PWMF/RemaTxNum[22]_keep ;
  wire \PWMF/RemaTxNum[23]_keep ;
  wire \PWMF/RemaTxNum[2]_keep ;
  wire \PWMF/RemaTxNum[3]_keep ;
  wire \PWMF/RemaTxNum[4]_keep ;
  wire \PWMF/RemaTxNum[5]_keep ;
  wire \PWMF/RemaTxNum[6]_keep ;
  wire \PWMF/RemaTxNum[7]_keep ;
  wire \PWMF/RemaTxNum[8]_keep ;
  wire \PWMF/RemaTxNum[9]_keep ;
  wire \PWMF/dir_keep ;
  wire \PWMF/mux3_b0_sel_is_3_o ;
  wire \PWMF/n0_lutinv ;
  wire \PWMF/n1 ;
  wire \PWMF/n10 ;
  wire \PWMF/n11 ;
  wire \PWMF/n24 ;
  wire \PWMF/n25_neg_lutinv ;
  wire \PWMF/n32 ;
  wire \PWMF/pnumr[0]_keep ;
  wire \PWMF/pnumr[10]_keep ;
  wire \PWMF/pnumr[11]_keep ;
  wire \PWMF/pnumr[12]_keep ;
  wire \PWMF/pnumr[13]_keep ;
  wire \PWMF/pnumr[14]_keep ;
  wire \PWMF/pnumr[15]_keep ;
  wire \PWMF/pnumr[16]_keep ;
  wire \PWMF/pnumr[17]_keep ;
  wire \PWMF/pnumr[18]_keep ;
  wire \PWMF/pnumr[19]_keep ;
  wire \PWMF/pnumr[1]_keep ;
  wire \PWMF/pnumr[20]_keep ;
  wire \PWMF/pnumr[21]_keep ;
  wire \PWMF/pnumr[22]_keep ;
  wire \PWMF/pnumr[23]_keep ;
  wire \PWMF/pnumr[24]_keep ;
  wire \PWMF/pnumr[25]_keep ;
  wire \PWMF/pnumr[26]_keep ;
  wire \PWMF/pnumr[27]_keep ;
  wire \PWMF/pnumr[28]_keep ;
  wire \PWMF/pnumr[29]_keep ;
  wire \PWMF/pnumr[2]_keep ;
  wire \PWMF/pnumr[30]_keep ;
  wire \PWMF/pnumr[31]_keep ;
  wire \PWMF/pnumr[3]_keep ;
  wire \PWMF/pnumr[4]_keep ;
  wire \PWMF/pnumr[5]_keep ;
  wire \PWMF/pnumr[6]_keep ;
  wire \PWMF/pnumr[7]_keep ;
  wire \PWMF/pnumr[8]_keep ;
  wire \PWMF/pnumr[9]_keep ;
  wire \PWMF/pwm_keep ;
  wire \PWMF/stopreq ;  // src/OnePWM.v(14)
  wire \PWMF/stopreq_keep ;
  wire \PWMF/sub0/c0 ;
  wire \PWMF/sub0/c1 ;
  wire \PWMF/sub0/c10 ;
  wire \PWMF/sub0/c11 ;
  wire \PWMF/sub0/c12 ;
  wire \PWMF/sub0/c13 ;
  wire \PWMF/sub0/c14 ;
  wire \PWMF/sub0/c15 ;
  wire \PWMF/sub0/c16 ;
  wire \PWMF/sub0/c17 ;
  wire \PWMF/sub0/c18 ;
  wire \PWMF/sub0/c19 ;
  wire \PWMF/sub0/c2 ;
  wire \PWMF/sub0/c20 ;
  wire \PWMF/sub0/c21 ;
  wire \PWMF/sub0/c22 ;
  wire \PWMF/sub0/c23 ;
  wire \PWMF/sub0/c24 ;
  wire \PWMF/sub0/c25 ;
  wire \PWMF/sub0/c26 ;
  wire \PWMF/sub0/c3 ;
  wire \PWMF/sub0/c4 ;
  wire \PWMF/sub0/c5 ;
  wire \PWMF/sub0/c6 ;
  wire \PWMF/sub0/c7 ;
  wire \PWMF/sub0/c8 ;
  wire \PWMF/sub0/c9 ;
  wire \PWMF/sub1/c0 ;
  wire \PWMF/sub1/c1 ;
  wire \PWMF/sub1/c10 ;
  wire \PWMF/sub1/c11 ;
  wire \PWMF/sub1/c12 ;
  wire \PWMF/sub1/c13 ;
  wire \PWMF/sub1/c14 ;
  wire \PWMF/sub1/c15 ;
  wire \PWMF/sub1/c16 ;
  wire \PWMF/sub1/c17 ;
  wire \PWMF/sub1/c18 ;
  wire \PWMF/sub1/c19 ;
  wire \PWMF/sub1/c2 ;
  wire \PWMF/sub1/c20 ;
  wire \PWMF/sub1/c21 ;
  wire \PWMF/sub1/c22 ;
  wire \PWMF/sub1/c23 ;
  wire \PWMF/sub1/c3 ;
  wire \PWMF/sub1/c4 ;
  wire \PWMF/sub1/c5 ;
  wire \PWMF/sub1/c6 ;
  wire \PWMF/sub1/c7 ;
  wire \PWMF/sub1/c8 ;
  wire \PWMF/sub1/c9 ;
  wire \PWMF/u14_sel_is_1_o ;
  wire \U_AHB/h2h_hwrite ;  // src/AHB.v(22)
  wire \U_AHB/h2h_hwritew ;  // src/AHB.v(19)
  wire \U_AHB/n10 ;
  wire \U_AHB/n102 ;
  wire \U_AHB/n104_lutinv ;
  wire \U_AHB/n105 ;
  wire \U_AHB/n108 ;
  wire \U_AHB/n111 ;
  wire \U_AHB/n113_lutinv ;
  wire \U_AHB/n12 ;
  wire \U_AHB/n14 ;
  wire \U_AHB/n16 ;
  wire \U_AHB/n18 ;
  wire \U_AHB/n2 ;
  wire \U_AHB/n20 ;
  wire \U_AHB/n22 ;
  wire \U_AHB/n24 ;
  wire \U_AHB/n26 ;
  wire \U_AHB/n28 ;
  wire \U_AHB/n30 ;
  wire \U_AHB/n32 ;
  wire \U_AHB/n34 ;
  wire \U_AHB/n36 ;
  wire \U_AHB/n38 ;
  wire \U_AHB/n4 ;
  wire \U_AHB/n45 ;
  wire \U_AHB/n47 ;
  wire \U_AHB/n51 ;
  wire \U_AHB/n53 ;
  wire \U_AHB/n55 ;
  wire \U_AHB/n57 ;
  wire \U_AHB/n59 ;
  wire \U_AHB/n61 ;
  wire \U_AHB/n63 ;
  wire \U_AHB/n65 ;
  wire \U_AHB/n67 ;
  wire \U_AHB/n69 ;
  wire \U_AHB/n71 ;
  wire \U_AHB/n73 ;
  wire \U_AHB/n75 ;
  wire \U_AHB/n77 ;
  wire \U_AHB/n79 ;
  wire \U_AHB/n8 ;
  wire \U_AHB/n82 ;
  wire \U_AHB/n87 ;
  wire \U_AHB/n90 ;
  wire \U_AHB/n93 ;
  wire \U_AHB/n95_lutinv ;
  wire \U_AHB/n96 ;
  wire \U_AHB/n99 ;
  wire _al_n1_en;
  wire _al_u1030_o;
  wire _al_u1031_o;
  wire _al_u1032_o;
  wire _al_u1033_o;
  wire _al_u1034_o;
  wire _al_u1035_o;
  wire _al_u1036_o;
  wire _al_u1067_o;
  wire _al_u1068_o;
  wire _al_u1069_o;
  wire _al_u1070_o;
  wire _al_u1071_o;
  wire _al_u1072_o;
  wire _al_u1073_o;
  wire _al_u1104_o;
  wire _al_u1105_o;
  wire _al_u1106_o;
  wire _al_u1107_o;
  wire _al_u1108_o;
  wire _al_u1109_o;
  wire _al_u1110_o;
  wire _al_u1141_o;
  wire _al_u1142_o;
  wire _al_u1143_o;
  wire _al_u1144_o;
  wire _al_u1145_o;
  wire _al_u1146_o;
  wire _al_u1147_o;
  wire _al_u1178_o;
  wire _al_u1179_o;
  wire _al_u1180_o;
  wire _al_u1181_o;
  wire _al_u1182_o;
  wire _al_u1183_o;
  wire _al_u1184_o;
  wire _al_u1215_o;
  wire _al_u1216_o;
  wire _al_u1217_o;
  wire _al_u1218_o;
  wire _al_u1219_o;
  wire _al_u1220_o;
  wire _al_u1221_o;
  wire _al_u1252_o;
  wire _al_u1253_o;
  wire _al_u1254_o;
  wire _al_u1255_o;
  wire _al_u1256_o;
  wire _al_u1257_o;
  wire _al_u1258_o;
  wire _al_u1289_o;
  wire _al_u1290_o;
  wire _al_u1291_o;
  wire _al_u1292_o;
  wire _al_u1293_o;
  wire _al_u1294_o;
  wire _al_u1295_o;
  wire _al_u1360_o;
  wire _al_u1361_o;
  wire _al_u1362_o;
  wire _al_u1363_o;
  wire _al_u1364_o;
  wire _al_u1365_o;
  wire _al_u1366_o;
  wire _al_u1367_o;
  wire _al_u1368_o;
  wire _al_u1369_o;
  wire _al_u1370_o;
  wire _al_u1371_o;
  wire _al_u1372_o;
  wire _al_u1373_o;
  wire _al_u1374_o;
  wire _al_u1375_o;
  wire _al_u1376_o;
  wire _al_u1378_o;
  wire _al_u1379_o;
  wire _al_u1380_o;
  wire _al_u1381_o;
  wire _al_u1382_o;
  wire _al_u1383_o;
  wire _al_u1384_o;
  wire _al_u1385_o;
  wire _al_u1386_o;
  wire _al_u1387_o;
  wire _al_u1388_o;
  wire _al_u1389_o;
  wire _al_u1390_o;
  wire _al_u1391_o;
  wire _al_u1392_o;
  wire _al_u1393_o;
  wire _al_u1395_o;
  wire _al_u1396_o;
  wire _al_u1397_o;
  wire _al_u1398_o;
  wire _al_u1399_o;
  wire _al_u1400_o;
  wire _al_u1401_o;
  wire _al_u1402_o;
  wire _al_u1403_o;
  wire _al_u1404_o;
  wire _al_u1405_o;
  wire _al_u1406_o;
  wire _al_u1407_o;
  wire _al_u1408_o;
  wire _al_u1409_o;
  wire _al_u1410_o;
  wire _al_u1411_o;
  wire _al_u1413_o;
  wire _al_u1414_o;
  wire _al_u1415_o;
  wire _al_u1416_o;
  wire _al_u1417_o;
  wire _al_u1418_o;
  wire _al_u1419_o;
  wire _al_u1420_o;
  wire _al_u1421_o;
  wire _al_u1422_o;
  wire _al_u1423_o;
  wire _al_u1424_o;
  wire _al_u1425_o;
  wire _al_u1426_o;
  wire _al_u1427_o;
  wire _al_u1428_o;
  wire _al_u1430_o;
  wire _al_u1431_o;
  wire _al_u1432_o;
  wire _al_u1433_o;
  wire _al_u1434_o;
  wire _al_u1435_o;
  wire _al_u1436_o;
  wire _al_u1437_o;
  wire _al_u1438_o;
  wire _al_u1439_o;
  wire _al_u1440_o;
  wire _al_u1441_o;
  wire _al_u1442_o;
  wire _al_u1443_o;
  wire _al_u1444_o;
  wire _al_u1445_o;
  wire _al_u1447_o;
  wire _al_u1448_o;
  wire _al_u1449_o;
  wire _al_u1450_o;
  wire _al_u1451_o;
  wire _al_u1452_o;
  wire _al_u1453_o;
  wire _al_u1454_o;
  wire _al_u1455_o;
  wire _al_u1456_o;
  wire _al_u1457_o;
  wire _al_u1458_o;
  wire _al_u1459_o;
  wire _al_u1460_o;
  wire _al_u1461_o;
  wire _al_u1462_o;
  wire _al_u1464_o;
  wire _al_u1465_o;
  wire _al_u1466_o;
  wire _al_u1467_o;
  wire _al_u1468_o;
  wire _al_u1469_o;
  wire _al_u1470_o;
  wire _al_u1471_o;
  wire _al_u1472_o;
  wire _al_u1473_o;
  wire _al_u1474_o;
  wire _al_u1475_o;
  wire _al_u1476_o;
  wire _al_u1477_o;
  wire _al_u1480_o;
  wire _al_u1481_o;
  wire _al_u1482_o;
  wire _al_u1483_o;
  wire _al_u1484_o;
  wire _al_u1485_o;
  wire _al_u1486_o;
  wire _al_u1487_o;
  wire _al_u1488_o;
  wire _al_u1489_o;
  wire _al_u1490_o;
  wire _al_u1491_o;
  wire _al_u1492_o;
  wire _al_u1493_o;
  wire _al_u1494_o;
  wire _al_u1495_o;
  wire _al_u1496_o;
  wire _al_u1498_o;
  wire _al_u1499_o;
  wire _al_u1500_o;
  wire _al_u1501_o;
  wire _al_u1502_o;
  wire _al_u1503_o;
  wire _al_u1504_o;
  wire _al_u1505_o;
  wire _al_u1506_o;
  wire _al_u1507_o;
  wire _al_u1508_o;
  wire _al_u1509_o;
  wire _al_u1510_o;
  wire _al_u1511_o;
  wire _al_u1512_o;
  wire _al_u1513_o;
  wire _al_u1514_o;
  wire _al_u1516_o;
  wire _al_u1517_o;
  wire _al_u1518_o;
  wire _al_u1519_o;
  wire _al_u1520_o;
  wire _al_u1521_o;
  wire _al_u1522_o;
  wire _al_u1523_o;
  wire _al_u1524_o;
  wire _al_u1525_o;
  wire _al_u1526_o;
  wire _al_u1527_o;
  wire _al_u1528_o;
  wire _al_u1529_o;
  wire _al_u1530_o;
  wire _al_u1531_o;
  wire _al_u1533_o;
  wire _al_u1534_o;
  wire _al_u1535_o;
  wire _al_u1536_o;
  wire _al_u1537_o;
  wire _al_u1538_o;
  wire _al_u1539_o;
  wire _al_u1540_o;
  wire _al_u1541_o;
  wire _al_u1542_o;
  wire _al_u1543_o;
  wire _al_u1544_o;
  wire _al_u1545_o;
  wire _al_u1546_o;
  wire _al_u1547_o;
  wire _al_u1548_o;
  wire _al_u1549_o;
  wire _al_u1551_o;
  wire _al_u1552_o;
  wire _al_u1553_o;
  wire _al_u1554_o;
  wire _al_u1555_o;
  wire _al_u1556_o;
  wire _al_u1557_o;
  wire _al_u1558_o;
  wire _al_u1559_o;
  wire _al_u1560_o;
  wire _al_u1561_o;
  wire _al_u1562_o;
  wire _al_u1563_o;
  wire _al_u1564_o;
  wire _al_u1565_o;
  wire _al_u1566_o;
  wire _al_u1568_o;
  wire _al_u1569_o;
  wire _al_u1570_o;
  wire _al_u1571_o;
  wire _al_u1572_o;
  wire _al_u1573_o;
  wire _al_u1574_o;
  wire _al_u1575_o;
  wire _al_u1576_o;
  wire _al_u1577_o;
  wire _al_u1578_o;
  wire _al_u1579_o;
  wire _al_u1580_o;
  wire _al_u1581_o;
  wire _al_u1582_o;
  wire _al_u1583_o;
  wire _al_u1585_o;
  wire _al_u1586_o;
  wire _al_u1587_o;
  wire _al_u1588_o;
  wire _al_u1589_o;
  wire _al_u1590_o;
  wire _al_u1591_o;
  wire _al_u1592_o;
  wire _al_u1593_o;
  wire _al_u1594_o;
  wire _al_u1595_o;
  wire _al_u1596_o;
  wire _al_u1597_o;
  wire _al_u1598_o;
  wire _al_u1599_o;
  wire _al_u1600_o;
  wire _al_u1602_o;
  wire _al_u1603_o;
  wire _al_u1604_o;
  wire _al_u1605_o;
  wire _al_u1606_o;
  wire _al_u1607_o;
  wire _al_u1608_o;
  wire _al_u1609_o;
  wire _al_u1610_o;
  wire _al_u1611_o;
  wire _al_u1612_o;
  wire _al_u1613_o;
  wire _al_u1614_o;
  wire _al_u1615_o;
  wire _al_u1616_o;
  wire _al_u1617_o;
  wire _al_u1618_o;
  wire _al_u1620_o;
  wire _al_u1621_o;
  wire _al_u1622_o;
  wire _al_u1623_o;
  wire _al_u1624_o;
  wire _al_u1625_o;
  wire _al_u1626_o;
  wire _al_u1627_o;
  wire _al_u1628_o;
  wire _al_u1629_o;
  wire _al_u1630_o;
  wire _al_u1631_o;
  wire _al_u1632_o;
  wire _al_u1633_o;
  wire _al_u1634_o;
  wire _al_u1635_o;
  wire _al_u1636_o;
  wire _al_u1638_o;
  wire _al_u1639_o;
  wire _al_u1640_o;
  wire _al_u1641_o;
  wire _al_u1642_o;
  wire _al_u1643_o;
  wire _al_u1644_o;
  wire _al_u1645_o;
  wire _al_u1647_o;
  wire _al_u1648_o;
  wire _al_u1649_o;
  wire _al_u1650_o;
  wire _al_u1651_o;
  wire _al_u1652_o;
  wire _al_u1686_o;
  wire _al_u1687_o;
  wire _al_u1688_o;
  wire _al_u1689_o;
  wire _al_u1690_o;
  wire _al_u1691_o;
  wire _al_u1693_o;
  wire _al_u1695_o;
  wire _al_u1697_o;
  wire _al_u1699_o;
  wire _al_u1701_o;
  wire _al_u1703_o;
  wire _al_u1705_o;
  wire _al_u1707_o;
  wire _al_u1709_o;
  wire _al_u1711_o;
  wire _al_u1713_o;
  wire _al_u1715_o;
  wire _al_u1717_o;
  wire _al_u1719_o;
  wire _al_u1721_o;
  wire _al_u1723_o;
  wire _al_u1725_o;
  wire _al_u1727_o;
  wire _al_u1729_o;
  wire _al_u1731_o;
  wire _al_u1733_o;
  wire _al_u1735_o;
  wire _al_u1737_o;
  wire _al_u1739_o;
  wire _al_u1741_o;
  wire _al_u1742_o;
  wire _al_u1743_o;
  wire _al_u1744_o;
  wire _al_u1745_o;
  wire _al_u1746_o;
  wire _al_u1747_o;
  wire _al_u1748_o;
  wire _al_u1749_o;
  wire _al_u1750_o;
  wire _al_u1751_o;
  wire _al_u1752_o;
  wire _al_u1753_o;
  wire _al_u1754_o;
  wire _al_u1755_o;
  wire _al_u1756_o;
  wire _al_u1757_o;
  wire _al_u1758_o;
  wire _al_u1759_o;
  wire _al_u1760_o;
  wire _al_u1761_o;
  wire _al_u1762_o;
  wire _al_u1763_o;
  wire _al_u1764_o;
  wire _al_u1765_o;
  wire _al_u1768_o;
  wire _al_u1769_o;
  wire _al_u1770_o;
  wire _al_u1771_o;
  wire _al_u1772_o;
  wire _al_u1773_o;
  wire _al_u1775_o;
  wire _al_u1777_o;
  wire _al_u1779_o;
  wire _al_u1781_o;
  wire _al_u1783_o;
  wire _al_u1785_o;
  wire _al_u1787_o;
  wire _al_u1789_o;
  wire _al_u1791_o;
  wire _al_u1793_o;
  wire _al_u1795_o;
  wire _al_u1797_o;
  wire _al_u1799_o;
  wire _al_u1801_o;
  wire _al_u1803_o;
  wire _al_u1805_o;
  wire _al_u1807_o;
  wire _al_u1809_o;
  wire _al_u1811_o;
  wire _al_u1813_o;
  wire _al_u1815_o;
  wire _al_u1817_o;
  wire _al_u1819_o;
  wire _al_u1821_o;
  wire _al_u1823_o;
  wire _al_u1824_o;
  wire _al_u1825_o;
  wire _al_u1826_o;
  wire _al_u1827_o;
  wire _al_u1828_o;
  wire _al_u1829_o;
  wire _al_u1830_o;
  wire _al_u1831_o;
  wire _al_u1832_o;
  wire _al_u1833_o;
  wire _al_u1834_o;
  wire _al_u1835_o;
  wire _al_u1836_o;
  wire _al_u1837_o;
  wire _al_u1838_o;
  wire _al_u1839_o;
  wire _al_u1840_o;
  wire _al_u1841_o;
  wire _al_u1842_o;
  wire _al_u1843_o;
  wire _al_u1844_o;
  wire _al_u1845_o;
  wire _al_u1846_o;
  wire _al_u1847_o;
  wire _al_u1850_o;
  wire _al_u1851_o;
  wire _al_u1852_o;
  wire _al_u1853_o;
  wire _al_u1854_o;
  wire _al_u1855_o;
  wire _al_u1857_o;
  wire _al_u1859_o;
  wire _al_u1861_o;
  wire _al_u1863_o;
  wire _al_u1865_o;
  wire _al_u1867_o;
  wire _al_u1869_o;
  wire _al_u1871_o;
  wire _al_u1873_o;
  wire _al_u1875_o;
  wire _al_u1877_o;
  wire _al_u1879_o;
  wire _al_u1881_o;
  wire _al_u1883_o;
  wire _al_u1885_o;
  wire _al_u1887_o;
  wire _al_u1889_o;
  wire _al_u1891_o;
  wire _al_u1893_o;
  wire _al_u1895_o;
  wire _al_u1897_o;
  wire _al_u1899_o;
  wire _al_u1901_o;
  wire _al_u1903_o;
  wire _al_u1905_o;
  wire _al_u1906_o;
  wire _al_u1907_o;
  wire _al_u1908_o;
  wire _al_u1909_o;
  wire _al_u1910_o;
  wire _al_u1911_o;
  wire _al_u1912_o;
  wire _al_u1913_o;
  wire _al_u1914_o;
  wire _al_u1915_o;
  wire _al_u1916_o;
  wire _al_u1917_o;
  wire _al_u1918_o;
  wire _al_u1919_o;
  wire _al_u1920_o;
  wire _al_u1921_o;
  wire _al_u1922_o;
  wire _al_u1923_o;
  wire _al_u1924_o;
  wire _al_u1925_o;
  wire _al_u1926_o;
  wire _al_u1927_o;
  wire _al_u1930_o;
  wire _al_u1931_o;
  wire _al_u1932_o;
  wire _al_u1933_o;
  wire _al_u1934_o;
  wire _al_u1935_o;
  wire _al_u1937_o;
  wire _al_u1939_o;
  wire _al_u1941_o;
  wire _al_u1943_o;
  wire _al_u1945_o;
  wire _al_u1947_o;
  wire _al_u1949_o;
  wire _al_u1951_o;
  wire _al_u1953_o;
  wire _al_u1955_o;
  wire _al_u1957_o;
  wire _al_u1959_o;
  wire _al_u1961_o;
  wire _al_u1963_o;
  wire _al_u1965_o;
  wire _al_u1967_o;
  wire _al_u1969_o;
  wire _al_u1971_o;
  wire _al_u1973_o;
  wire _al_u1975_o;
  wire _al_u1977_o;
  wire _al_u1979_o;
  wire _al_u1981_o;
  wire _al_u1983_o;
  wire _al_u1985_o;
  wire _al_u1986_o;
  wire _al_u1987_o;
  wire _al_u1988_o;
  wire _al_u1989_o;
  wire _al_u1990_o;
  wire _al_u1991_o;
  wire _al_u1992_o;
  wire _al_u1993_o;
  wire _al_u1994_o;
  wire _al_u1995_o;
  wire _al_u1996_o;
  wire _al_u1997_o;
  wire _al_u1998_o;
  wire _al_u1999_o;
  wire _al_u2000_o;
  wire _al_u2001_o;
  wire _al_u2002_o;
  wire _al_u2003_o;
  wire _al_u2004_o;
  wire _al_u2005_o;
  wire _al_u2006_o;
  wire _al_u2007_o;
  wire _al_u2008_o;
  wire _al_u2009_o;
  wire _al_u2012_o;
  wire _al_u2013_o;
  wire _al_u2014_o;
  wire _al_u2015_o;
  wire _al_u2016_o;
  wire _al_u2017_o;
  wire _al_u2019_o;
  wire _al_u2021_o;
  wire _al_u2023_o;
  wire _al_u2025_o;
  wire _al_u2027_o;
  wire _al_u2029_o;
  wire _al_u2031_o;
  wire _al_u2033_o;
  wire _al_u2035_o;
  wire _al_u2037_o;
  wire _al_u2039_o;
  wire _al_u2041_o;
  wire _al_u2043_o;
  wire _al_u2045_o;
  wire _al_u2047_o;
  wire _al_u2049_o;
  wire _al_u2051_o;
  wire _al_u2053_o;
  wire _al_u2055_o;
  wire _al_u2057_o;
  wire _al_u2059_o;
  wire _al_u2061_o;
  wire _al_u2063_o;
  wire _al_u2065_o;
  wire _al_u2067_o;
  wire _al_u2068_o;
  wire _al_u2069_o;
  wire _al_u2070_o;
  wire _al_u2071_o;
  wire _al_u2072_o;
  wire _al_u2073_o;
  wire _al_u2074_o;
  wire _al_u2075_o;
  wire _al_u2076_o;
  wire _al_u2077_o;
  wire _al_u2078_o;
  wire _al_u2079_o;
  wire _al_u2080_o;
  wire _al_u2081_o;
  wire _al_u2082_o;
  wire _al_u2083_o;
  wire _al_u2084_o;
  wire _al_u2085_o;
  wire _al_u2086_o;
  wire _al_u2087_o;
  wire _al_u2088_o;
  wire _al_u2089_o;
  wire _al_u2090_o;
  wire _al_u2091_o;
  wire _al_u2094_o;
  wire _al_u2095_o;
  wire _al_u2096_o;
  wire _al_u2097_o;
  wire _al_u2098_o;
  wire _al_u2099_o;
  wire _al_u2101_o;
  wire _al_u2103_o;
  wire _al_u2105_o;
  wire _al_u2107_o;
  wire _al_u2109_o;
  wire _al_u2111_o;
  wire _al_u2113_o;
  wire _al_u2115_o;
  wire _al_u2117_o;
  wire _al_u2119_o;
  wire _al_u2121_o;
  wire _al_u2123_o;
  wire _al_u2125_o;
  wire _al_u2127_o;
  wire _al_u2129_o;
  wire _al_u2131_o;
  wire _al_u2133_o;
  wire _al_u2135_o;
  wire _al_u2137_o;
  wire _al_u2139_o;
  wire _al_u2141_o;
  wire _al_u2143_o;
  wire _al_u2145_o;
  wire _al_u2147_o;
  wire _al_u2149_o;
  wire _al_u2150_o;
  wire _al_u2151_o;
  wire _al_u2152_o;
  wire _al_u2153_o;
  wire _al_u2154_o;
  wire _al_u2155_o;
  wire _al_u2156_o;
  wire _al_u2157_o;
  wire _al_u2158_o;
  wire _al_u2159_o;
  wire _al_u2160_o;
  wire _al_u2161_o;
  wire _al_u2162_o;
  wire _al_u2163_o;
  wire _al_u2164_o;
  wire _al_u2165_o;
  wire _al_u2166_o;
  wire _al_u2167_o;
  wire _al_u2168_o;
  wire _al_u2169_o;
  wire _al_u2170_o;
  wire _al_u2171_o;
  wire _al_u2172_o;
  wire _al_u2173_o;
  wire _al_u2176_o;
  wire _al_u2177_o;
  wire _al_u2178_o;
  wire _al_u2179_o;
  wire _al_u2180_o;
  wire _al_u2181_o;
  wire _al_u2183_o;
  wire _al_u2185_o;
  wire _al_u2187_o;
  wire _al_u2189_o;
  wire _al_u2191_o;
  wire _al_u2193_o;
  wire _al_u2195_o;
  wire _al_u2197_o;
  wire _al_u2199_o;
  wire _al_u2201_o;
  wire _al_u2203_o;
  wire _al_u2205_o;
  wire _al_u2207_o;
  wire _al_u2209_o;
  wire _al_u2211_o;
  wire _al_u2213_o;
  wire _al_u2215_o;
  wire _al_u2217_o;
  wire _al_u2219_o;
  wire _al_u2221_o;
  wire _al_u2223_o;
  wire _al_u2225_o;
  wire _al_u2227_o;
  wire _al_u2229_o;
  wire _al_u2231_o;
  wire _al_u2232_o;
  wire _al_u2233_o;
  wire _al_u2234_o;
  wire _al_u2235_o;
  wire _al_u2236_o;
  wire _al_u2237_o;
  wire _al_u2238_o;
  wire _al_u2239_o;
  wire _al_u2240_o;
  wire _al_u2241_o;
  wire _al_u2242_o;
  wire _al_u2243_o;
  wire _al_u2244_o;
  wire _al_u2245_o;
  wire _al_u2246_o;
  wire _al_u2247_o;
  wire _al_u2248_o;
  wire _al_u2249_o;
  wire _al_u2250_o;
  wire _al_u2251_o;
  wire _al_u2252_o;
  wire _al_u2253_o;
  wire _al_u2256_o;
  wire _al_u2257_o;
  wire _al_u2258_o;
  wire _al_u2259_o;
  wire _al_u2260_o;
  wire _al_u2261_o;
  wire _al_u2263_o;
  wire _al_u2265_o;
  wire _al_u2267_o;
  wire _al_u2269_o;
  wire _al_u2271_o;
  wire _al_u2273_o;
  wire _al_u2275_o;
  wire _al_u2277_o;
  wire _al_u2279_o;
  wire _al_u2281_o;
  wire _al_u2283_o;
  wire _al_u2285_o;
  wire _al_u2287_o;
  wire _al_u2289_o;
  wire _al_u2291_o;
  wire _al_u2293_o;
  wire _al_u2295_o;
  wire _al_u2297_o;
  wire _al_u2299_o;
  wire _al_u2301_o;
  wire _al_u2303_o;
  wire _al_u2305_o;
  wire _al_u2307_o;
  wire _al_u2309_o;
  wire _al_u2311_o;
  wire _al_u2312_o;
  wire _al_u2313_o;
  wire _al_u2314_o;
  wire _al_u2315_o;
  wire _al_u2316_o;
  wire _al_u2317_o;
  wire _al_u2318_o;
  wire _al_u2319_o;
  wire _al_u2320_o;
  wire _al_u2321_o;
  wire _al_u2322_o;
  wire _al_u2323_o;
  wire _al_u2324_o;
  wire _al_u2325_o;
  wire _al_u2326_o;
  wire _al_u2327_o;
  wire _al_u2328_o;
  wire _al_u2329_o;
  wire _al_u2330_o;
  wire _al_u2331_o;
  wire _al_u2332_o;
  wire _al_u2333_o;
  wire _al_u2334_o;
  wire _al_u2335_o;
  wire _al_u2338_o;
  wire _al_u2339_o;
  wire _al_u2340_o;
  wire _al_u2341_o;
  wire _al_u2342_o;
  wire _al_u2343_o;
  wire _al_u2345_o;
  wire _al_u2347_o;
  wire _al_u2349_o;
  wire _al_u2351_o;
  wire _al_u2353_o;
  wire _al_u2355_o;
  wire _al_u2357_o;
  wire _al_u2359_o;
  wire _al_u2361_o;
  wire _al_u2363_o;
  wire _al_u2365_o;
  wire _al_u2367_o;
  wire _al_u2369_o;
  wire _al_u2371_o;
  wire _al_u2373_o;
  wire _al_u2375_o;
  wire _al_u2377_o;
  wire _al_u2379_o;
  wire _al_u2381_o;
  wire _al_u2383_o;
  wire _al_u2385_o;
  wire _al_u2387_o;
  wire _al_u2389_o;
  wire _al_u2391_o;
  wire _al_u2393_o;
  wire _al_u2394_o;
  wire _al_u2395_o;
  wire _al_u2396_o;
  wire _al_u2397_o;
  wire _al_u2398_o;
  wire _al_u2399_o;
  wire _al_u2400_o;
  wire _al_u2401_o;
  wire _al_u2402_o;
  wire _al_u2403_o;
  wire _al_u2404_o;
  wire _al_u2405_o;
  wire _al_u2406_o;
  wire _al_u2407_o;
  wire _al_u2408_o;
  wire _al_u2409_o;
  wire _al_u2410_o;
  wire _al_u2411_o;
  wire _al_u2412_o;
  wire _al_u2413_o;
  wire _al_u2414_o;
  wire _al_u2415_o;
  wire _al_u2418_o;
  wire _al_u2419_o;
  wire _al_u2420_o;
  wire _al_u2421_o;
  wire _al_u2422_o;
  wire _al_u2423_o;
  wire _al_u2425_o;
  wire _al_u2427_o;
  wire _al_u2429_o;
  wire _al_u2431_o;
  wire _al_u2433_o;
  wire _al_u2435_o;
  wire _al_u2437_o;
  wire _al_u2439_o;
  wire _al_u2441_o;
  wire _al_u2443_o;
  wire _al_u2445_o;
  wire _al_u2447_o;
  wire _al_u2449_o;
  wire _al_u2451_o;
  wire _al_u2453_o;
  wire _al_u2455_o;
  wire _al_u2457_o;
  wire _al_u2459_o;
  wire _al_u2461_o;
  wire _al_u2463_o;
  wire _al_u2465_o;
  wire _al_u2467_o;
  wire _al_u2469_o;
  wire _al_u2471_o;
  wire _al_u2473_o;
  wire _al_u2474_o;
  wire _al_u2475_o;
  wire _al_u2476_o;
  wire _al_u2477_o;
  wire _al_u2478_o;
  wire _al_u2479_o;
  wire _al_u2480_o;
  wire _al_u2481_o;
  wire _al_u2482_o;
  wire _al_u2483_o;
  wire _al_u2484_o;
  wire _al_u2485_o;
  wire _al_u2486_o;
  wire _al_u2487_o;
  wire _al_u2488_o;
  wire _al_u2489_o;
  wire _al_u2490_o;
  wire _al_u2491_o;
  wire _al_u2492_o;
  wire _al_u2493_o;
  wire _al_u2494_o;
  wire _al_u2495_o;
  wire _al_u2496_o;
  wire _al_u2497_o;
  wire _al_u2500_o;
  wire _al_u2501_o;
  wire _al_u2502_o;
  wire _al_u2503_o;
  wire _al_u2504_o;
  wire _al_u2505_o;
  wire _al_u2507_o;
  wire _al_u2509_o;
  wire _al_u2511_o;
  wire _al_u2513_o;
  wire _al_u2515_o;
  wire _al_u2517_o;
  wire _al_u2519_o;
  wire _al_u2521_o;
  wire _al_u2523_o;
  wire _al_u2525_o;
  wire _al_u2527_o;
  wire _al_u2529_o;
  wire _al_u2531_o;
  wire _al_u2533_o;
  wire _al_u2535_o;
  wire _al_u2537_o;
  wire _al_u2539_o;
  wire _al_u2541_o;
  wire _al_u2543_o;
  wire _al_u2545_o;
  wire _al_u2547_o;
  wire _al_u2549_o;
  wire _al_u2551_o;
  wire _al_u2553_o;
  wire _al_u2555_o;
  wire _al_u2556_o;
  wire _al_u2557_o;
  wire _al_u2558_o;
  wire _al_u2559_o;
  wire _al_u2560_o;
  wire _al_u2561_o;
  wire _al_u2562_o;
  wire _al_u2563_o;
  wire _al_u2564_o;
  wire _al_u2565_o;
  wire _al_u2566_o;
  wire _al_u2567_o;
  wire _al_u2568_o;
  wire _al_u2569_o;
  wire _al_u2570_o;
  wire _al_u2571_o;
  wire _al_u2572_o;
  wire _al_u2573_o;
  wire _al_u2574_o;
  wire _al_u2575_o;
  wire _al_u2576_o;
  wire _al_u2579_o;
  wire _al_u2580_o;
  wire _al_u2581_o;
  wire _al_u2582_o;
  wire _al_u2583_o;
  wire _al_u2584_o;
  wire _al_u2586_o;
  wire _al_u2588_o;
  wire _al_u2590_o;
  wire _al_u2592_o;
  wire _al_u2594_o;
  wire _al_u2596_o;
  wire _al_u2598_o;
  wire _al_u2600_o;
  wire _al_u2602_o;
  wire _al_u2604_o;
  wire _al_u2606_o;
  wire _al_u2608_o;
  wire _al_u2610_o;
  wire _al_u2612_o;
  wire _al_u2614_o;
  wire _al_u2616_o;
  wire _al_u2618_o;
  wire _al_u2620_o;
  wire _al_u2622_o;
  wire _al_u2624_o;
  wire _al_u2626_o;
  wire _al_u2628_o;
  wire _al_u2630_o;
  wire _al_u2632_o;
  wire _al_u2634_o;
  wire _al_u2635_o;
  wire _al_u2636_o;
  wire _al_u2637_o;
  wire _al_u2638_o;
  wire _al_u2639_o;
  wire _al_u2640_o;
  wire _al_u2641_o;
  wire _al_u2642_o;
  wire _al_u2643_o;
  wire _al_u2644_o;
  wire _al_u2645_o;
  wire _al_u2646_o;
  wire _al_u2647_o;
  wire _al_u2648_o;
  wire _al_u2649_o;
  wire _al_u2650_o;
  wire _al_u2651_o;
  wire _al_u2652_o;
  wire _al_u2653_o;
  wire _al_u2654_o;
  wire _al_u2655_o;
  wire _al_u2656_o;
  wire _al_u2657_o;
  wire _al_u2658_o;
  wire _al_u2661_o;
  wire _al_u2662_o;
  wire _al_u2663_o;
  wire _al_u2664_o;
  wire _al_u2665_o;
  wire _al_u2666_o;
  wire _al_u2668_o;
  wire _al_u2670_o;
  wire _al_u2672_o;
  wire _al_u2674_o;
  wire _al_u2676_o;
  wire _al_u2678_o;
  wire _al_u2680_o;
  wire _al_u2682_o;
  wire _al_u2684_o;
  wire _al_u2686_o;
  wire _al_u2688_o;
  wire _al_u2690_o;
  wire _al_u2692_o;
  wire _al_u2694_o;
  wire _al_u2696_o;
  wire _al_u2698_o;
  wire _al_u2700_o;
  wire _al_u2702_o;
  wire _al_u2704_o;
  wire _al_u2706_o;
  wire _al_u2708_o;
  wire _al_u2710_o;
  wire _al_u2712_o;
  wire _al_u2714_o;
  wire _al_u2716_o;
  wire _al_u2717_o;
  wire _al_u2718_o;
  wire _al_u2719_o;
  wire _al_u2720_o;
  wire _al_u2721_o;
  wire _al_u2722_o;
  wire _al_u2723_o;
  wire _al_u2724_o;
  wire _al_u2725_o;
  wire _al_u2726_o;
  wire _al_u2727_o;
  wire _al_u2728_o;
  wire _al_u2729_o;
  wire _al_u2730_o;
  wire _al_u2731_o;
  wire _al_u2732_o;
  wire _al_u2733_o;
  wire _al_u2734_o;
  wire _al_u2735_o;
  wire _al_u2736_o;
  wire _al_u2737_o;
  wire _al_u2740_o;
  wire _al_u2741_o;
  wire _al_u2742_o;
  wire _al_u2743_o;
  wire _al_u2744_o;
  wire _al_u2745_o;
  wire _al_u2747_o;
  wire _al_u2749_o;
  wire _al_u2751_o;
  wire _al_u2753_o;
  wire _al_u2755_o;
  wire _al_u2757_o;
  wire _al_u2759_o;
  wire _al_u2761_o;
  wire _al_u2763_o;
  wire _al_u2765_o;
  wire _al_u2767_o;
  wire _al_u2769_o;
  wire _al_u2771_o;
  wire _al_u2773_o;
  wire _al_u2775_o;
  wire _al_u2777_o;
  wire _al_u2779_o;
  wire _al_u2781_o;
  wire _al_u2783_o;
  wire _al_u2785_o;
  wire _al_u2787_o;
  wire _al_u2789_o;
  wire _al_u2791_o;
  wire _al_u2793_o;
  wire _al_u2795_o;
  wire _al_u2796_o;
  wire _al_u2797_o;
  wire _al_u2798_o;
  wire _al_u2799_o;
  wire _al_u2800_o;
  wire _al_u2801_o;
  wire _al_u2802_o;
  wire _al_u2803_o;
  wire _al_u2804_o;
  wire _al_u2805_o;
  wire _al_u2806_o;
  wire _al_u2807_o;
  wire _al_u2808_o;
  wire _al_u2809_o;
  wire _al_u2810_o;
  wire _al_u2811_o;
  wire _al_u2812_o;
  wire _al_u2813_o;
  wire _al_u2814_o;
  wire _al_u2815_o;
  wire _al_u2816_o;
  wire _al_u2817_o;
  wire _al_u2820_o;
  wire _al_u2821_o;
  wire _al_u2822_o;
  wire _al_u2823_o;
  wire _al_u2824_o;
  wire _al_u2825_o;
  wire _al_u2827_o;
  wire _al_u2829_o;
  wire _al_u2831_o;
  wire _al_u2833_o;
  wire _al_u2835_o;
  wire _al_u2837_o;
  wire _al_u2839_o;
  wire _al_u2841_o;
  wire _al_u2843_o;
  wire _al_u2845_o;
  wire _al_u2847_o;
  wire _al_u2849_o;
  wire _al_u2851_o;
  wire _al_u2853_o;
  wire _al_u2855_o;
  wire _al_u2857_o;
  wire _al_u2859_o;
  wire _al_u2861_o;
  wire _al_u2863_o;
  wire _al_u2865_o;
  wire _al_u2867_o;
  wire _al_u2869_o;
  wire _al_u2871_o;
  wire _al_u2873_o;
  wire _al_u2875_o;
  wire _al_u2876_o;
  wire _al_u2877_o;
  wire _al_u2878_o;
  wire _al_u2879_o;
  wire _al_u2880_o;
  wire _al_u2881_o;
  wire _al_u2882_o;
  wire _al_u2883_o;
  wire _al_u2884_o;
  wire _al_u2885_o;
  wire _al_u2886_o;
  wire _al_u2887_o;
  wire _al_u2888_o;
  wire _al_u2889_o;
  wire _al_u2890_o;
  wire _al_u2891_o;
  wire _al_u2892_o;
  wire _al_u2893_o;
  wire _al_u2894_o;
  wire _al_u2895_o;
  wire _al_u2896_o;
  wire _al_u2899_o;
  wire _al_u2900_o;
  wire _al_u2901_o;
  wire _al_u2902_o;
  wire _al_u2903_o;
  wire _al_u2904_o;
  wire _al_u2906_o;
  wire _al_u2908_o;
  wire _al_u2910_o;
  wire _al_u2912_o;
  wire _al_u2914_o;
  wire _al_u2916_o;
  wire _al_u2918_o;
  wire _al_u2920_o;
  wire _al_u2922_o;
  wire _al_u2924_o;
  wire _al_u2926_o;
  wire _al_u2928_o;
  wire _al_u2930_o;
  wire _al_u2932_o;
  wire _al_u2934_o;
  wire _al_u2936_o;
  wire _al_u2938_o;
  wire _al_u2940_o;
  wire _al_u2942_o;
  wire _al_u2944_o;
  wire _al_u2946_o;
  wire _al_u2948_o;
  wire _al_u2950_o;
  wire _al_u2952_o;
  wire _al_u2954_o;
  wire _al_u2955_o;
  wire _al_u2956_o;
  wire _al_u2957_o;
  wire _al_u2958_o;
  wire _al_u2959_o;
  wire _al_u2960_o;
  wire _al_u2961_o;
  wire _al_u2962_o;
  wire _al_u2963_o;
  wire _al_u2964_o;
  wire _al_u2965_o;
  wire _al_u2966_o;
  wire _al_u2967_o;
  wire _al_u2968_o;
  wire _al_u2969_o;
  wire _al_u2970_o;
  wire _al_u2971_o;
  wire _al_u2972_o;
  wire _al_u2973_o;
  wire _al_u2974_o;
  wire _al_u2975_o;
  wire _al_u2976_o;
  wire _al_u2977_o;
  wire _al_u2978_o;
  wire _al_u2980_o;
  wire _al_u2981_o;
  wire _al_u2982_o;
  wire _al_u2983_o;
  wire _al_u2984_o;
  wire _al_u2985_o;
  wire _al_u2986_o;
  wire _al_u2987_o;
  wire _al_u2988_o;
  wire _al_u3007_o;
  wire _al_u3008_o;
  wire _al_u3010_o;
  wire _al_u3011_o;
  wire _al_u3013_o;
  wire _al_u3014_o;
  wire _al_u3016_o;
  wire _al_u3017_o;
  wire _al_u3019_o;
  wire _al_u3020_o;
  wire _al_u3022_o;
  wire _al_u3023_o;
  wire _al_u3025_o;
  wire _al_u3026_o;
  wire _al_u3028_o;
  wire _al_u3029_o;
  wire _al_u3031_o;
  wire _al_u3032_o;
  wire _al_u3034_o;
  wire _al_u3035_o;
  wire _al_u3037_o;
  wire _al_u3038_o;
  wire _al_u3040_o;
  wire _al_u3041_o;
  wire _al_u3043_o;
  wire _al_u3044_o;
  wire _al_u3046_o;
  wire _al_u3047_o;
  wire _al_u3049_o;
  wire _al_u3050_o;
  wire _al_u3052_o;
  wire _al_u3053_o;
  wire _al_u3055_o;
  wire _al_u3061_o;
  wire _al_u3062_o;
  wire _al_u3065_o;
  wire _al_u3068_o;
  wire _al_u3070_o;
  wire _al_u3072_o;
  wire _al_u3074_o;
  wire _al_u3076_o;
  wire _al_u3078_o;
  wire _al_u3080_o;
  wire _al_u3082_o;
  wire _al_u3085_o;
  wire _al_u3087_o;
  wire _al_u3089_o;
  wire _al_u3092_o;
  wire _al_u3094_o;
  wire _al_u3095_o;
  wire _al_u3096_o;
  wire _al_u3097_o;
  wire _al_u3098_o;
  wire _al_u3100_o;
  wire _al_u3101_o;
  wire _al_u3102_o;
  wire _al_u3103_o;
  wire _al_u3104_o;
  wire _al_u3105_o;
  wire _al_u3106_o;
  wire _al_u3107_o;
  wire _al_u3108_o;
  wire _al_u3109_o;
  wire _al_u3111_o;
  wire _al_u3112_o;
  wire _al_u3113_o;
  wire _al_u3114_o;
  wire _al_u3115_o;
  wire _al_u3116_o;
  wire _al_u3117_o;
  wire _al_u3118_o;
  wire _al_u3119_o;
  wire _al_u3120_o;
  wire _al_u3122_o;
  wire _al_u3123_o;
  wire _al_u3124_o;
  wire _al_u3125_o;
  wire _al_u3126_o;
  wire _al_u3127_o;
  wire _al_u3128_o;
  wire _al_u3129_o;
  wire _al_u3130_o;
  wire _al_u3131_o;
  wire _al_u3133_o;
  wire _al_u3134_o;
  wire _al_u3135_o;
  wire _al_u3136_o;
  wire _al_u3137_o;
  wire _al_u3138_o;
  wire _al_u3139_o;
  wire _al_u3140_o;
  wire _al_u3141_o;
  wire _al_u3142_o;
  wire _al_u3143_o;
  wire _al_u3145_o;
  wire _al_u3146_o;
  wire _al_u3147_o;
  wire _al_u3148_o;
  wire _al_u3149_o;
  wire _al_u3150_o;
  wire _al_u3151_o;
  wire _al_u3152_o;
  wire _al_u3153_o;
  wire _al_u3154_o;
  wire _al_u3156_o;
  wire _al_u3157_o;
  wire _al_u3158_o;
  wire _al_u3159_o;
  wire _al_u3160_o;
  wire _al_u3161_o;
  wire _al_u3162_o;
  wire _al_u3163_o;
  wire _al_u3164_o;
  wire _al_u3165_o;
  wire _al_u3167_o;
  wire _al_u3168_o;
  wire _al_u3169_o;
  wire _al_u3170_o;
  wire _al_u3171_o;
  wire _al_u3172_o;
  wire _al_u3173_o;
  wire _al_u3174_o;
  wire _al_u3175_o;
  wire _al_u3176_o;
  wire _al_u3178_o;
  wire _al_u3179_o;
  wire _al_u3180_o;
  wire _al_u3181_o;
  wire _al_u3182_o;
  wire _al_u3183_o;
  wire _al_u3184_o;
  wire _al_u3185_o;
  wire _al_u3186_o;
  wire _al_u3187_o;
  wire _al_u3189_o;
  wire _al_u3190_o;
  wire _al_u3191_o;
  wire _al_u3192_o;
  wire _al_u3193_o;
  wire _al_u3194_o;
  wire _al_u3195_o;
  wire _al_u3196_o;
  wire _al_u3197_o;
  wire _al_u3198_o;
  wire _al_u3200_o;
  wire _al_u3201_o;
  wire _al_u3202_o;
  wire _al_u3203_o;
  wire _al_u3204_o;
  wire _al_u3205_o;
  wire _al_u3206_o;
  wire _al_u3207_o;
  wire _al_u3208_o;
  wire _al_u3209_o;
  wire _al_u3211_o;
  wire _al_u3212_o;
  wire _al_u3213_o;
  wire _al_u3214_o;
  wire _al_u3215_o;
  wire _al_u3216_o;
  wire _al_u3217_o;
  wire _al_u3218_o;
  wire _al_u3219_o;
  wire _al_u3220_o;
  wire _al_u3222_o;
  wire _al_u3223_o;
  wire _al_u3224_o;
  wire _al_u3225_o;
  wire _al_u3226_o;
  wire _al_u3227_o;
  wire _al_u3228_o;
  wire _al_u3229_o;
  wire _al_u3230_o;
  wire _al_u3231_o;
  wire _al_u3233_o;
  wire _al_u3234_o;
  wire _al_u3235_o;
  wire _al_u3236_o;
  wire _al_u3237_o;
  wire _al_u3238_o;
  wire _al_u3239_o;
  wire _al_u3240_o;
  wire _al_u3241_o;
  wire _al_u3242_o;
  wire _al_u3244_o;
  wire _al_u3245_o;
  wire _al_u3246_o;
  wire _al_u3247_o;
  wire _al_u3248_o;
  wire _al_u3249_o;
  wire _al_u3250_o;
  wire _al_u3251_o;
  wire _al_u3252_o;
  wire _al_u3253_o;
  wire _al_u3255_o;
  wire _al_u3256_o;
  wire _al_u3257_o;
  wire _al_u3258_o;
  wire _al_u3259_o;
  wire _al_u3260_o;
  wire _al_u3261_o;
  wire _al_u3262_o;
  wire _al_u3263_o;
  wire _al_u3264_o;
  wire _al_u3266_o;
  wire _al_u3267_o;
  wire _al_u3268_o;
  wire _al_u3269_o;
  wire _al_u3270_o;
  wire _al_u3271_o;
  wire _al_u3272_o;
  wire _al_u3273_o;
  wire _al_u3274_o;
  wire _al_u3275_o;
  wire _al_u3277_o;
  wire _al_u3278_o;
  wire _al_u3279_o;
  wire _al_u3280_o;
  wire _al_u3281_o;
  wire _al_u3282_o;
  wire _al_u3283_o;
  wire _al_u3284_o;
  wire _al_u3285_o;
  wire _al_u3286_o;
  wire _al_u3288_o;
  wire _al_u3289_o;
  wire _al_u3290_o;
  wire _al_u3291_o;
  wire _al_u3292_o;
  wire _al_u3293_o;
  wire _al_u3294_o;
  wire _al_u3295_o;
  wire _al_u3296_o;
  wire _al_u3297_o;
  wire _al_u3299_o;
  wire _al_u3300_o;
  wire _al_u3301_o;
  wire _al_u3302_o;
  wire _al_u3303_o;
  wire _al_u3304_o;
  wire _al_u3305_o;
  wire _al_u3306_o;
  wire _al_u3307_o;
  wire _al_u3308_o;
  wire _al_u3310_o;
  wire _al_u3311_o;
  wire _al_u3312_o;
  wire _al_u3313_o;
  wire _al_u3314_o;
  wire _al_u3315_o;
  wire _al_u3316_o;
  wire _al_u3317_o;
  wire _al_u3318_o;
  wire _al_u3319_o;
  wire _al_u3321_o;
  wire _al_u3322_o;
  wire _al_u3323_o;
  wire _al_u3324_o;
  wire _al_u3325_o;
  wire _al_u3326_o;
  wire _al_u3327_o;
  wire _al_u3328_o;
  wire _al_u3329_o;
  wire _al_u3330_o;
  wire _al_u3332_o;
  wire _al_u3333_o;
  wire _al_u3334_o;
  wire _al_u3335_o;
  wire _al_u3336_o;
  wire _al_u3337_o;
  wire _al_u3338_o;
  wire _al_u3339_o;
  wire _al_u3340_o;
  wire _al_u3341_o;
  wire _al_u3343_o;
  wire _al_u3344_o;
  wire _al_u3345_o;
  wire _al_u3346_o;
  wire _al_u3347_o;
  wire _al_u3348_o;
  wire _al_u3349_o;
  wire _al_u3350_o;
  wire _al_u3351_o;
  wire _al_u3352_o;
  wire _al_u734_o;
  wire _al_u735_o;
  wire _al_u736_o;
  wire _al_u737_o;
  wire _al_u738_o;
  wire _al_u739_o;
  wire _al_u740_o;
  wire _al_u771_o;
  wire _al_u772_o;
  wire _al_u773_o;
  wire _al_u774_o;
  wire _al_u775_o;
  wire _al_u776_o;
  wire _al_u777_o;
  wire _al_u808_o;
  wire _al_u809_o;
  wire _al_u810_o;
  wire _al_u811_o;
  wire _al_u812_o;
  wire _al_u813_o;
  wire _al_u814_o;
  wire _al_u845_o;
  wire _al_u846_o;
  wire _al_u847_o;
  wire _al_u848_o;
  wire _al_u849_o;
  wire _al_u850_o;
  wire _al_u851_o;
  wire _al_u882_o;
  wire _al_u883_o;
  wire _al_u884_o;
  wire _al_u885_o;
  wire _al_u886_o;
  wire _al_u887_o;
  wire _al_u888_o;
  wire _al_u919_o;
  wire _al_u920_o;
  wire _al_u921_o;
  wire _al_u922_o;
  wire _al_u923_o;
  wire _al_u924_o;
  wire _al_u925_o;
  wire _al_u956_o;
  wire _al_u957_o;
  wire _al_u958_o;
  wire _al_u959_o;
  wire _al_u960_o;
  wire _al_u961_o;
  wire _al_u962_o;
  wire _al_u993_o;
  wire _al_u994_o;
  wire _al_u995_o;
  wire _al_u996_o;
  wire _al_u997_o;
  wire _al_u998_o;
  wire _al_u999_o;
  wire \add0/c0 ;
  wire \add0/c1 ;
  wire \add0/c10 ;
  wire \add0/c11 ;
  wire \add0/c12 ;
  wire \add0/c13 ;
  wire \add0/c14 ;
  wire \add0/c15 ;
  wire \add0/c16 ;
  wire \add0/c17 ;
  wire \add0/c18 ;
  wire \add0/c19 ;
  wire \add0/c2 ;
  wire \add0/c20 ;
  wire \add0/c21 ;
  wire \add0/c22 ;
  wire \add0/c23 ;
  wire \add0/c24 ;
  wire \add0/c25 ;
  wire \add0/c26 ;
  wire \add0/c27 ;
  wire \add0/c28 ;
  wire \add0/c29 ;
  wire \add0/c3 ;
  wire \add0/c30 ;
  wire \add0/c31 ;
  wire \add0/c4 ;
  wire \add0/c5 ;
  wire \add0/c6 ;
  wire \add0/c7 ;
  wire \add0/c8 ;
  wire \add0/c9 ;
  wire clk100m;  // CPLD_SOC_AHB_TOP.v(13)
  wire clk100m_keep;
  wire clk25m;  // CPLD_SOC_AHB_TOP.v(13)
  wire clkin_pad;  // CPLD_SOC_AHB_TOP.v(3)
  wire n4_neg;
  wire \pwm[0]_d ;
  wire \pwm[10]_d ;
  wire \pwm[11]_d ;
  wire \pwm[12]_d ;
  wire \pwm[13]_d ;
  wire \pwm[14]_d ;
  wire \pwm[15]_d ;
  wire \pwm[1]_d ;
  wire \pwm[2]_d ;
  wire \pwm[3]_d ;
  wire \pwm[4]_d ;
  wire \pwm[5]_d ;
  wire \pwm[6]_d ;
  wire \pwm[7]_d ;
  wire \pwm[8]_d ;
  wire \pwm[9]_d ;
  wire rst_n_pad;  // CPLD_SOC_AHB_TOP.v(4)
  wire rstn;  // CPLD_SOC_AHB_TOP.v(13)

  reg_ar_as_w1 \PWM0/State_reg  (
    .clk(clk100m),
    .d(\PWM0/n10 ),
    .en(1'b1),
    .reset(~rstn),
    .set(1'b0),
    .q(pwm_state_read[0]));  // src/OnePWM.v(26)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[0]  (
    .i(\PWM0/RemaTxNum[0]_keep ),
    .o(pnumcnt0[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[10]  (
    .i(\PWM0/RemaTxNum[10]_keep ),
    .o(pnumcnt0[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[11]  (
    .i(\PWM0/RemaTxNum[11]_keep ),
    .o(pnumcnt0[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[12]  (
    .i(\PWM0/RemaTxNum[12]_keep ),
    .o(pnumcnt0[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[13]  (
    .i(\PWM0/RemaTxNum[13]_keep ),
    .o(pnumcnt0[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[14]  (
    .i(\PWM0/RemaTxNum[14]_keep ),
    .o(pnumcnt0[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[15]  (
    .i(\PWM0/RemaTxNum[15]_keep ),
    .o(pnumcnt0[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[16]  (
    .i(\PWM0/RemaTxNum[16]_keep ),
    .o(pnumcnt0[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[17]  (
    .i(\PWM0/RemaTxNum[17]_keep ),
    .o(pnumcnt0[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[18]  (
    .i(\PWM0/RemaTxNum[18]_keep ),
    .o(pnumcnt0[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[19]  (
    .i(\PWM0/RemaTxNum[19]_keep ),
    .o(pnumcnt0[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[1]  (
    .i(\PWM0/RemaTxNum[1]_keep ),
    .o(pnumcnt0[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[20]  (
    .i(\PWM0/RemaTxNum[20]_keep ),
    .o(pnumcnt0[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[21]  (
    .i(\PWM0/RemaTxNum[21]_keep ),
    .o(pnumcnt0[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[22]  (
    .i(\PWM0/RemaTxNum[22]_keep ),
    .o(pnumcnt0[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[23]  (
    .i(\PWM0/RemaTxNum[23]_keep ),
    .o(pnumcnt0[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[2]  (
    .i(\PWM0/RemaTxNum[2]_keep ),
    .o(pnumcnt0[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[3]  (
    .i(\PWM0/RemaTxNum[3]_keep ),
    .o(pnumcnt0[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[4]  (
    .i(\PWM0/RemaTxNum[4]_keep ),
    .o(pnumcnt0[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[5]  (
    .i(\PWM0/RemaTxNum[5]_keep ),
    .o(pnumcnt0[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[6]  (
    .i(\PWM0/RemaTxNum[6]_keep ),
    .o(pnumcnt0[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[7]  (
    .i(\PWM0/RemaTxNum[7]_keep ),
    .o(pnumcnt0[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[8]  (
    .i(\PWM0/RemaTxNum[8]_keep ),
    .o(pnumcnt0[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[9]  (
    .i(\PWM0/RemaTxNum[9]_keep ),
    .o(pnumcnt0[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_dir  (
    .i(\PWM0/dir_keep ),
    .o(dir_pad[0]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[0]  (
    .i(\PWM0/pnumr[0]_keep ),
    .o(\PWM0/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[10]  (
    .i(\PWM0/pnumr[10]_keep ),
    .o(\PWM0/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[11]  (
    .i(\PWM0/pnumr[11]_keep ),
    .o(\PWM0/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[12]  (
    .i(\PWM0/pnumr[12]_keep ),
    .o(\PWM0/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[13]  (
    .i(\PWM0/pnumr[13]_keep ),
    .o(\PWM0/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[14]  (
    .i(\PWM0/pnumr[14]_keep ),
    .o(\PWM0/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[15]  (
    .i(\PWM0/pnumr[15]_keep ),
    .o(\PWM0/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[16]  (
    .i(\PWM0/pnumr[16]_keep ),
    .o(\PWM0/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[17]  (
    .i(\PWM0/pnumr[17]_keep ),
    .o(\PWM0/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[18]  (
    .i(\PWM0/pnumr[18]_keep ),
    .o(\PWM0/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[19]  (
    .i(\PWM0/pnumr[19]_keep ),
    .o(\PWM0/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[1]  (
    .i(\PWM0/pnumr[1]_keep ),
    .o(\PWM0/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[20]  (
    .i(\PWM0/pnumr[20]_keep ),
    .o(\PWM0/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[21]  (
    .i(\PWM0/pnumr[21]_keep ),
    .o(\PWM0/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[22]  (
    .i(\PWM0/pnumr[22]_keep ),
    .o(\PWM0/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[23]  (
    .i(\PWM0/pnumr[23]_keep ),
    .o(\PWM0/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[24]  (
    .i(\PWM0/pnumr[24]_keep ),
    .o(\PWM0/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[25]  (
    .i(\PWM0/pnumr[25]_keep ),
    .o(\PWM0/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[26]  (
    .i(\PWM0/pnumr[26]_keep ),
    .o(\PWM0/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[27]  (
    .i(\PWM0/pnumr[27]_keep ),
    .o(\PWM0/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[28]  (
    .i(\PWM0/pnumr[28]_keep ),
    .o(\PWM0/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[29]  (
    .i(\PWM0/pnumr[29]_keep ),
    .o(\PWM0/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[2]  (
    .i(\PWM0/pnumr[2]_keep ),
    .o(\PWM0/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[30]  (
    .i(\PWM0/pnumr[30]_keep ),
    .o(\PWM0/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[31]  (
    .i(\PWM0/pnumr[31]_keep ),
    .o(\PWM0/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[3]  (
    .i(\PWM0/pnumr[3]_keep ),
    .o(\PWM0/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[4]  (
    .i(\PWM0/pnumr[4]_keep ),
    .o(\PWM0/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[5]  (
    .i(\PWM0/pnumr[5]_keep ),
    .o(\PWM0/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[6]  (
    .i(\PWM0/pnumr[6]_keep ),
    .o(\PWM0/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[7]  (
    .i(\PWM0/pnumr[7]_keep ),
    .o(\PWM0/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[8]  (
    .i(\PWM0/pnumr[8]_keep ),
    .o(\PWM0/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[9]  (
    .i(\PWM0/pnumr[9]_keep ),
    .o(\PWM0/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pwm  (
    .i(\PWM0/pwm_keep ),
    .o(pwm_pad[0]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_stopreq  (
    .i(\PWM0/stopreq_keep ),
    .o(\PWM0/stopreq ));  // src/OnePWM.v(14)
  reg_ar_as_w1 \PWM0/dir_reg  (
    .clk(clk100m),
    .d(\PWM0/n32 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/dir_keep ));  // src/OnePWM.v(58)
  reg_sr_as_w1 \PWM0/pwm_reg  (
    .clk(clk100m),
    .d(\pwm[0]_d ),
    .en(1'b1),
    .reset(~\PWM0/u14_sel_is_1_o ),
    .set(1'b0),
    .q(\PWM0/pwm_keep ));  // src/OnePWM.v(45)
  reg_sr_as_w1 \PWM0/reg0_b0  (
    .clk(clk100m),
    .d(\PWM0/n13 [0]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [0]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b1  (
    .clk(clk100m),
    .d(\PWM0/n13 [1]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [1]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b10  (
    .clk(clk100m),
    .d(\PWM0/n13 [10]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [10]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b11  (
    .clk(clk100m),
    .d(\PWM0/n13 [11]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [11]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b12  (
    .clk(clk100m),
    .d(\PWM0/n13 [12]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [12]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b13  (
    .clk(clk100m),
    .d(\PWM0/n13 [13]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [13]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b14  (
    .clk(clk100m),
    .d(\PWM0/n13 [14]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [14]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b15  (
    .clk(clk100m),
    .d(\PWM0/n13 [15]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [15]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b16  (
    .clk(clk100m),
    .d(\PWM0/n13 [16]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [16]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b17  (
    .clk(clk100m),
    .d(\PWM0/n13 [17]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [17]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b18  (
    .clk(clk100m),
    .d(\PWM0/n13 [18]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [18]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b19  (
    .clk(clk100m),
    .d(\PWM0/n13 [19]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [19]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b2  (
    .clk(clk100m),
    .d(\PWM0/n13 [2]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [2]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b20  (
    .clk(clk100m),
    .d(\PWM0/n13 [20]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [20]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b21  (
    .clk(clk100m),
    .d(\PWM0/n13 [21]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [21]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b22  (
    .clk(clk100m),
    .d(\PWM0/n13 [22]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [22]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b23  (
    .clk(clk100m),
    .d(\PWM0/n13 [23]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [23]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b24  (
    .clk(clk100m),
    .d(\PWM0/n13 [24]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [24]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b25  (
    .clk(clk100m),
    .d(\PWM0/n13 [25]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [25]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b26  (
    .clk(clk100m),
    .d(\PWM0/n13 [26]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [26]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b3  (
    .clk(clk100m),
    .d(\PWM0/n13 [3]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [3]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b4  (
    .clk(clk100m),
    .d(\PWM0/n13 [4]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [4]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b5  (
    .clk(clk100m),
    .d(\PWM0/n13 [5]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [5]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b6  (
    .clk(clk100m),
    .d(\PWM0/n13 [6]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [6]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b7  (
    .clk(clk100m),
    .d(\PWM0/n13 [7]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [7]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b8  (
    .clk(clk100m),
    .d(\PWM0/n13 [8]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [8]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b9  (
    .clk(clk100m),
    .d(\PWM0/n13 [9]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b0  (
    .clk(clk100m),
    .d(freq0[0]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [0]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b1  (
    .clk(clk100m),
    .d(freq0[1]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [1]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b10  (
    .clk(clk100m),
    .d(freq0[10]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [10]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b11  (
    .clk(clk100m),
    .d(freq0[11]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [11]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b12  (
    .clk(clk100m),
    .d(freq0[12]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [12]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b13  (
    .clk(clk100m),
    .d(freq0[13]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [13]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b14  (
    .clk(clk100m),
    .d(freq0[14]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [14]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b15  (
    .clk(clk100m),
    .d(freq0[15]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [15]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b16  (
    .clk(clk100m),
    .d(freq0[16]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [16]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b17  (
    .clk(clk100m),
    .d(freq0[17]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [17]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b18  (
    .clk(clk100m),
    .d(freq0[18]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [18]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b19  (
    .clk(clk100m),
    .d(freq0[19]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [19]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b2  (
    .clk(clk100m),
    .d(freq0[2]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [2]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b20  (
    .clk(clk100m),
    .d(freq0[20]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [20]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b21  (
    .clk(clk100m),
    .d(freq0[21]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [21]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b22  (
    .clk(clk100m),
    .d(freq0[22]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [22]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b23  (
    .clk(clk100m),
    .d(freq0[23]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [23]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b24  (
    .clk(clk100m),
    .d(freq0[24]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [24]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b25  (
    .clk(clk100m),
    .d(freq0[25]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [25]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b26  (
    .clk(clk100m),
    .d(freq0[26]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [26]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b3  (
    .clk(clk100m),
    .d(freq0[3]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [3]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b4  (
    .clk(clk100m),
    .d(freq0[4]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [4]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b5  (
    .clk(clk100m),
    .d(freq0[5]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [5]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b6  (
    .clk(clk100m),
    .d(freq0[6]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [6]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b7  (
    .clk(clk100m),
    .d(freq0[7]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [7]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b8  (
    .clk(clk100m),
    .d(freq0[8]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [8]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b9  (
    .clk(clk100m),
    .d(freq0[9]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg2_b0  (
    .clk(clk100m),
    .d(\PWM0/n23 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[0]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b1  (
    .clk(clk100m),
    .d(\PWM0/n23 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[1]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b10  (
    .clk(clk100m),
    .d(\PWM0/n23 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[10]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b11  (
    .clk(clk100m),
    .d(\PWM0/n23 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[11]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b12  (
    .clk(clk100m),
    .d(\PWM0/n23 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[12]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b13  (
    .clk(clk100m),
    .d(\PWM0/n23 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[13]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b14  (
    .clk(clk100m),
    .d(\PWM0/n23 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[14]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b15  (
    .clk(clk100m),
    .d(\PWM0/n23 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[15]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b16  (
    .clk(clk100m),
    .d(\PWM0/n23 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[16]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b17  (
    .clk(clk100m),
    .d(\PWM0/n23 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[17]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b18  (
    .clk(clk100m),
    .d(\PWM0/n23 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[18]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b19  (
    .clk(clk100m),
    .d(\PWM0/n23 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[19]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b2  (
    .clk(clk100m),
    .d(\PWM0/n23 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[2]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b20  (
    .clk(clk100m),
    .d(\PWM0/n23 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[20]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b21  (
    .clk(clk100m),
    .d(\PWM0/n23 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[21]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b22  (
    .clk(clk100m),
    .d(\PWM0/n23 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[22]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b23  (
    .clk(clk100m),
    .d(\PWM0/n23 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[23]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b24  (
    .clk(clk100m),
    .d(\PWM0/n23 [24]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[24]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b25  (
    .clk(clk100m),
    .d(\PWM0/n23 [25]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[25]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b26  (
    .clk(clk100m),
    .d(\PWM0/n23 [26]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[26]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b27  (
    .clk(clk100m),
    .d(\PWM0/n23 [27]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[27]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b28  (
    .clk(clk100m),
    .d(\PWM0/n23 [28]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[28]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b29  (
    .clk(clk100m),
    .d(\PWM0/n23 [29]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[29]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b3  (
    .clk(clk100m),
    .d(\PWM0/n23 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[3]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b30  (
    .clk(clk100m),
    .d(\PWM0/n23 [30]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[30]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b31  (
    .clk(clk100m),
    .d(\PWM0/n23 [31]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[31]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b4  (
    .clk(clk100m),
    .d(\PWM0/n23 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[4]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b5  (
    .clk(clk100m),
    .d(\PWM0/n23 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[5]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b6  (
    .clk(clk100m),
    .d(\PWM0/n23 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[6]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b7  (
    .clk(clk100m),
    .d(\PWM0/n23 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[7]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b8  (
    .clk(clk100m),
    .d(\PWM0/n23 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[8]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b9  (
    .clk(clk100m),
    .d(\PWM0/n23 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[9]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg3_b0  (
    .clk(clk100m),
    .d(\PWM0/n31 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[0]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b1  (
    .clk(clk100m),
    .d(\PWM0/n31 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[1]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b10  (
    .clk(clk100m),
    .d(\PWM0/n31 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[10]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b11  (
    .clk(clk100m),
    .d(\PWM0/n31 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[11]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b12  (
    .clk(clk100m),
    .d(\PWM0/n31 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[12]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b13  (
    .clk(clk100m),
    .d(\PWM0/n31 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[13]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b14  (
    .clk(clk100m),
    .d(\PWM0/n31 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[14]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b15  (
    .clk(clk100m),
    .d(\PWM0/n31 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[15]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b16  (
    .clk(clk100m),
    .d(\PWM0/n31 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[16]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b17  (
    .clk(clk100m),
    .d(\PWM0/n31 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[17]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b18  (
    .clk(clk100m),
    .d(\PWM0/n31 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[18]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b19  (
    .clk(clk100m),
    .d(\PWM0/n31 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[19]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b2  (
    .clk(clk100m),
    .d(\PWM0/n31 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[2]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b20  (
    .clk(clk100m),
    .d(\PWM0/n31 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[20]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b21  (
    .clk(clk100m),
    .d(\PWM0/n31 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[21]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b22  (
    .clk(clk100m),
    .d(\PWM0/n31 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[22]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b23  (
    .clk(clk100m),
    .d(\PWM0/n31 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[23]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b3  (
    .clk(clk100m),
    .d(\PWM0/n31 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[3]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b4  (
    .clk(clk100m),
    .d(\PWM0/n31 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[4]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b5  (
    .clk(clk100m),
    .d(\PWM0/n31 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[5]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b6  (
    .clk(clk100m),
    .d(\PWM0/n31 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[6]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b7  (
    .clk(clk100m),
    .d(\PWM0/n31 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[7]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b8  (
    .clk(clk100m),
    .d(\PWM0/n31 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[8]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b9  (
    .clk(clk100m),
    .d(\PWM0/n31 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[9]_keep ));  // src/OnePWM.v(58)
  reg_ar_ss_w1 \PWM0/stopreq_reg  (
    .clk(clk100m),
    .d(\PWM0/n1 ),
    .en(1'b1),
    .reset(1'b0),
    .set(pwm_start_stop[0]),
    .q(\PWM0/stopreq_keep ));  // src/OnePWM.v(15)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub0/u0  (
    .a(\PWM0/FreCnt [0]),
    .b(1'b1),
    .c(\PWM0/sub0/c0 ),
    .o({\PWM0/sub0/c1 ,\PWM0/n12 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub0/u1  (
    .a(\PWM0/FreCnt [1]),
    .b(1'b0),
    .c(\PWM0/sub0/c1 ),
    .o({\PWM0/sub0/c2 ,\PWM0/n12 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub0/u10  (
    .a(\PWM0/FreCnt [10]),
    .b(1'b0),
    .c(\PWM0/sub0/c10 ),
    .o({\PWM0/sub0/c11 ,\PWM0/n12 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub0/u11  (
    .a(\PWM0/FreCnt [11]),
    .b(1'b0),
    .c(\PWM0/sub0/c11 ),
    .o({\PWM0/sub0/c12 ,\PWM0/n12 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub0/u12  (
    .a(\PWM0/FreCnt [12]),
    .b(1'b0),
    .c(\PWM0/sub0/c12 ),
    .o({\PWM0/sub0/c13 ,\PWM0/n12 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub0/u13  (
    .a(\PWM0/FreCnt [13]),
    .b(1'b0),
    .c(\PWM0/sub0/c13 ),
    .o({\PWM0/sub0/c14 ,\PWM0/n12 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub0/u14  (
    .a(\PWM0/FreCnt [14]),
    .b(1'b0),
    .c(\PWM0/sub0/c14 ),
    .o({\PWM0/sub0/c15 ,\PWM0/n12 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub0/u15  (
    .a(\PWM0/FreCnt [15]),
    .b(1'b0),
    .c(\PWM0/sub0/c15 ),
    .o({\PWM0/sub0/c16 ,\PWM0/n12 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub0/u16  (
    .a(\PWM0/FreCnt [16]),
    .b(1'b0),
    .c(\PWM0/sub0/c16 ),
    .o({\PWM0/sub0/c17 ,\PWM0/n12 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub0/u17  (
    .a(\PWM0/FreCnt [17]),
    .b(1'b0),
    .c(\PWM0/sub0/c17 ),
    .o({\PWM0/sub0/c18 ,\PWM0/n12 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub0/u18  (
    .a(\PWM0/FreCnt [18]),
    .b(1'b0),
    .c(\PWM0/sub0/c18 ),
    .o({\PWM0/sub0/c19 ,\PWM0/n12 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub0/u19  (
    .a(\PWM0/FreCnt [19]),
    .b(1'b0),
    .c(\PWM0/sub0/c19 ),
    .o({\PWM0/sub0/c20 ,\PWM0/n12 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub0/u2  (
    .a(\PWM0/FreCnt [2]),
    .b(1'b0),
    .c(\PWM0/sub0/c2 ),
    .o({\PWM0/sub0/c3 ,\PWM0/n12 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub0/u20  (
    .a(\PWM0/FreCnt [20]),
    .b(1'b0),
    .c(\PWM0/sub0/c20 ),
    .o({\PWM0/sub0/c21 ,\PWM0/n12 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub0/u21  (
    .a(\PWM0/FreCnt [21]),
    .b(1'b0),
    .c(\PWM0/sub0/c21 ),
    .o({\PWM0/sub0/c22 ,\PWM0/n12 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub0/u22  (
    .a(\PWM0/FreCnt [22]),
    .b(1'b0),
    .c(\PWM0/sub0/c22 ),
    .o({\PWM0/sub0/c23 ,\PWM0/n12 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub0/u23  (
    .a(\PWM0/FreCnt [23]),
    .b(1'b0),
    .c(\PWM0/sub0/c23 ),
    .o({\PWM0/sub0/c24 ,\PWM0/n12 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub0/u24  (
    .a(\PWM0/FreCnt [24]),
    .b(1'b0),
    .c(\PWM0/sub0/c24 ),
    .o({\PWM0/sub0/c25 ,\PWM0/n12 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub0/u25  (
    .a(\PWM0/FreCnt [25]),
    .b(1'b0),
    .c(\PWM0/sub0/c25 ),
    .o({\PWM0/sub0/c26 ,\PWM0/n12 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub0/u26  (
    .a(\PWM0/FreCnt [26]),
    .b(1'b0),
    .c(\PWM0/sub0/c26 ),
    .o({open_n0,\PWM0/n12 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub0/u3  (
    .a(\PWM0/FreCnt [3]),
    .b(1'b0),
    .c(\PWM0/sub0/c3 ),
    .o({\PWM0/sub0/c4 ,\PWM0/n12 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub0/u4  (
    .a(\PWM0/FreCnt [4]),
    .b(1'b0),
    .c(\PWM0/sub0/c4 ),
    .o({\PWM0/sub0/c5 ,\PWM0/n12 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub0/u5  (
    .a(\PWM0/FreCnt [5]),
    .b(1'b0),
    .c(\PWM0/sub0/c5 ),
    .o({\PWM0/sub0/c6 ,\PWM0/n12 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub0/u6  (
    .a(\PWM0/FreCnt [6]),
    .b(1'b0),
    .c(\PWM0/sub0/c6 ),
    .o({\PWM0/sub0/c7 ,\PWM0/n12 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub0/u7  (
    .a(\PWM0/FreCnt [7]),
    .b(1'b0),
    .c(\PWM0/sub0/c7 ),
    .o({\PWM0/sub0/c8 ,\PWM0/n12 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub0/u8  (
    .a(\PWM0/FreCnt [8]),
    .b(1'b0),
    .c(\PWM0/sub0/c8 ),
    .o({\PWM0/sub0/c9 ,\PWM0/n12 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub0/u9  (
    .a(\PWM0/FreCnt [9]),
    .b(1'b0),
    .c(\PWM0/sub0/c9 ),
    .o({\PWM0/sub0/c10 ,\PWM0/n12 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \PWM0/sub0/ucin  (
    .a(1'b0),
    .o({\PWM0/sub0/c0 ,open_n3}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub1/u0  (
    .a(pnumcnt0[0]),
    .b(1'b1),
    .c(\PWM0/sub1/c0 ),
    .o({\PWM0/sub1/c1 ,\PWM0/n26 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub1/u1  (
    .a(pnumcnt0[1]),
    .b(1'b0),
    .c(\PWM0/sub1/c1 ),
    .o({\PWM0/sub1/c2 ,\PWM0/n26 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub1/u10  (
    .a(pnumcnt0[10]),
    .b(1'b0),
    .c(\PWM0/sub1/c10 ),
    .o({\PWM0/sub1/c11 ,\PWM0/n26 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub1/u11  (
    .a(pnumcnt0[11]),
    .b(1'b0),
    .c(\PWM0/sub1/c11 ),
    .o({\PWM0/sub1/c12 ,\PWM0/n26 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub1/u12  (
    .a(pnumcnt0[12]),
    .b(1'b0),
    .c(\PWM0/sub1/c12 ),
    .o({\PWM0/sub1/c13 ,\PWM0/n26 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub1/u13  (
    .a(pnumcnt0[13]),
    .b(1'b0),
    .c(\PWM0/sub1/c13 ),
    .o({\PWM0/sub1/c14 ,\PWM0/n26 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub1/u14  (
    .a(pnumcnt0[14]),
    .b(1'b0),
    .c(\PWM0/sub1/c14 ),
    .o({\PWM0/sub1/c15 ,\PWM0/n26 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub1/u15  (
    .a(pnumcnt0[15]),
    .b(1'b0),
    .c(\PWM0/sub1/c15 ),
    .o({\PWM0/sub1/c16 ,\PWM0/n26 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub1/u16  (
    .a(pnumcnt0[16]),
    .b(1'b0),
    .c(\PWM0/sub1/c16 ),
    .o({\PWM0/sub1/c17 ,\PWM0/n26 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub1/u17  (
    .a(pnumcnt0[17]),
    .b(1'b0),
    .c(\PWM0/sub1/c17 ),
    .o({\PWM0/sub1/c18 ,\PWM0/n26 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub1/u18  (
    .a(pnumcnt0[18]),
    .b(1'b0),
    .c(\PWM0/sub1/c18 ),
    .o({\PWM0/sub1/c19 ,\PWM0/n26 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub1/u19  (
    .a(pnumcnt0[19]),
    .b(1'b0),
    .c(\PWM0/sub1/c19 ),
    .o({\PWM0/sub1/c20 ,\PWM0/n26 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub1/u2  (
    .a(pnumcnt0[2]),
    .b(1'b0),
    .c(\PWM0/sub1/c2 ),
    .o({\PWM0/sub1/c3 ,\PWM0/n26 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub1/u20  (
    .a(pnumcnt0[20]),
    .b(1'b0),
    .c(\PWM0/sub1/c20 ),
    .o({\PWM0/sub1/c21 ,\PWM0/n26 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub1/u21  (
    .a(pnumcnt0[21]),
    .b(1'b0),
    .c(\PWM0/sub1/c21 ),
    .o({\PWM0/sub1/c22 ,\PWM0/n26 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub1/u22  (
    .a(pnumcnt0[22]),
    .b(1'b0),
    .c(\PWM0/sub1/c22 ),
    .o({\PWM0/sub1/c23 ,\PWM0/n26 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub1/u23  (
    .a(pnumcnt0[23]),
    .b(1'b0),
    .c(\PWM0/sub1/c23 ),
    .o({open_n4,\PWM0/n26 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub1/u3  (
    .a(pnumcnt0[3]),
    .b(1'b0),
    .c(\PWM0/sub1/c3 ),
    .o({\PWM0/sub1/c4 ,\PWM0/n26 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub1/u4  (
    .a(pnumcnt0[4]),
    .b(1'b0),
    .c(\PWM0/sub1/c4 ),
    .o({\PWM0/sub1/c5 ,\PWM0/n26 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub1/u5  (
    .a(pnumcnt0[5]),
    .b(1'b0),
    .c(\PWM0/sub1/c5 ),
    .o({\PWM0/sub1/c6 ,\PWM0/n26 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub1/u6  (
    .a(pnumcnt0[6]),
    .b(1'b0),
    .c(\PWM0/sub1/c6 ),
    .o({\PWM0/sub1/c7 ,\PWM0/n26 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub1/u7  (
    .a(pnumcnt0[7]),
    .b(1'b0),
    .c(\PWM0/sub1/c7 ),
    .o({\PWM0/sub1/c8 ,\PWM0/n26 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub1/u8  (
    .a(pnumcnt0[8]),
    .b(1'b0),
    .c(\PWM0/sub1/c8 ),
    .o({\PWM0/sub1/c9 ,\PWM0/n26 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM0/sub1/u9  (
    .a(pnumcnt0[9]),
    .b(1'b0),
    .c(\PWM0/sub1/c9 ),
    .o({\PWM0/sub1/c10 ,\PWM0/n26 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \PWM0/sub1/ucin  (
    .a(1'b0),
    .o({\PWM0/sub1/c0 ,open_n7}));
  reg_ar_as_w1 \PWM1/State_reg  (
    .clk(clk100m),
    .d(\PWM1/n10 ),
    .en(1'b1),
    .reset(~rstn),
    .set(1'b0),
    .q(pwm_state_read[1]));  // src/OnePWM.v(26)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[0]  (
    .i(\PWM1/RemaTxNum[0]_keep ),
    .o(pnumcnt1[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[10]  (
    .i(\PWM1/RemaTxNum[10]_keep ),
    .o(pnumcnt1[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[11]  (
    .i(\PWM1/RemaTxNum[11]_keep ),
    .o(pnumcnt1[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[12]  (
    .i(\PWM1/RemaTxNum[12]_keep ),
    .o(pnumcnt1[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[13]  (
    .i(\PWM1/RemaTxNum[13]_keep ),
    .o(pnumcnt1[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[14]  (
    .i(\PWM1/RemaTxNum[14]_keep ),
    .o(pnumcnt1[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[15]  (
    .i(\PWM1/RemaTxNum[15]_keep ),
    .o(pnumcnt1[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[16]  (
    .i(\PWM1/RemaTxNum[16]_keep ),
    .o(pnumcnt1[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[17]  (
    .i(\PWM1/RemaTxNum[17]_keep ),
    .o(pnumcnt1[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[18]  (
    .i(\PWM1/RemaTxNum[18]_keep ),
    .o(pnumcnt1[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[19]  (
    .i(\PWM1/RemaTxNum[19]_keep ),
    .o(pnumcnt1[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[1]  (
    .i(\PWM1/RemaTxNum[1]_keep ),
    .o(pnumcnt1[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[20]  (
    .i(\PWM1/RemaTxNum[20]_keep ),
    .o(pnumcnt1[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[21]  (
    .i(\PWM1/RemaTxNum[21]_keep ),
    .o(pnumcnt1[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[22]  (
    .i(\PWM1/RemaTxNum[22]_keep ),
    .o(pnumcnt1[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[23]  (
    .i(\PWM1/RemaTxNum[23]_keep ),
    .o(pnumcnt1[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[2]  (
    .i(\PWM1/RemaTxNum[2]_keep ),
    .o(pnumcnt1[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[3]  (
    .i(\PWM1/RemaTxNum[3]_keep ),
    .o(pnumcnt1[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[4]  (
    .i(\PWM1/RemaTxNum[4]_keep ),
    .o(pnumcnt1[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[5]  (
    .i(\PWM1/RemaTxNum[5]_keep ),
    .o(pnumcnt1[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[6]  (
    .i(\PWM1/RemaTxNum[6]_keep ),
    .o(pnumcnt1[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[7]  (
    .i(\PWM1/RemaTxNum[7]_keep ),
    .o(pnumcnt1[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[8]  (
    .i(\PWM1/RemaTxNum[8]_keep ),
    .o(pnumcnt1[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[9]  (
    .i(\PWM1/RemaTxNum[9]_keep ),
    .o(pnumcnt1[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_dir  (
    .i(\PWM1/dir_keep ),
    .o(dir_pad[1]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[0]  (
    .i(\PWM1/pnumr[0]_keep ),
    .o(\PWM1/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[10]  (
    .i(\PWM1/pnumr[10]_keep ),
    .o(\PWM1/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[11]  (
    .i(\PWM1/pnumr[11]_keep ),
    .o(\PWM1/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[12]  (
    .i(\PWM1/pnumr[12]_keep ),
    .o(\PWM1/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[13]  (
    .i(\PWM1/pnumr[13]_keep ),
    .o(\PWM1/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[14]  (
    .i(\PWM1/pnumr[14]_keep ),
    .o(\PWM1/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[15]  (
    .i(\PWM1/pnumr[15]_keep ),
    .o(\PWM1/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[16]  (
    .i(\PWM1/pnumr[16]_keep ),
    .o(\PWM1/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[17]  (
    .i(\PWM1/pnumr[17]_keep ),
    .o(\PWM1/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[18]  (
    .i(\PWM1/pnumr[18]_keep ),
    .o(\PWM1/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[19]  (
    .i(\PWM1/pnumr[19]_keep ),
    .o(\PWM1/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[1]  (
    .i(\PWM1/pnumr[1]_keep ),
    .o(\PWM1/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[20]  (
    .i(\PWM1/pnumr[20]_keep ),
    .o(\PWM1/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[21]  (
    .i(\PWM1/pnumr[21]_keep ),
    .o(\PWM1/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[22]  (
    .i(\PWM1/pnumr[22]_keep ),
    .o(\PWM1/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[23]  (
    .i(\PWM1/pnumr[23]_keep ),
    .o(\PWM1/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[24]  (
    .i(\PWM1/pnumr[24]_keep ),
    .o(\PWM1/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[25]  (
    .i(\PWM1/pnumr[25]_keep ),
    .o(\PWM1/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[26]  (
    .i(\PWM1/pnumr[26]_keep ),
    .o(\PWM1/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[27]  (
    .i(\PWM1/pnumr[27]_keep ),
    .o(\PWM1/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[28]  (
    .i(\PWM1/pnumr[28]_keep ),
    .o(\PWM1/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[29]  (
    .i(\PWM1/pnumr[29]_keep ),
    .o(\PWM1/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[2]  (
    .i(\PWM1/pnumr[2]_keep ),
    .o(\PWM1/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[30]  (
    .i(\PWM1/pnumr[30]_keep ),
    .o(\PWM1/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[31]  (
    .i(\PWM1/pnumr[31]_keep ),
    .o(\PWM1/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[3]  (
    .i(\PWM1/pnumr[3]_keep ),
    .o(\PWM1/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[4]  (
    .i(\PWM1/pnumr[4]_keep ),
    .o(\PWM1/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[5]  (
    .i(\PWM1/pnumr[5]_keep ),
    .o(\PWM1/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[6]  (
    .i(\PWM1/pnumr[6]_keep ),
    .o(\PWM1/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[7]  (
    .i(\PWM1/pnumr[7]_keep ),
    .o(\PWM1/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[8]  (
    .i(\PWM1/pnumr[8]_keep ),
    .o(\PWM1/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[9]  (
    .i(\PWM1/pnumr[9]_keep ),
    .o(\PWM1/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pwm  (
    .i(\PWM1/pwm_keep ),
    .o(pwm_pad[1]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_stopreq  (
    .i(\PWM1/stopreq_keep ),
    .o(\PWM1/stopreq ));  // src/OnePWM.v(14)
  reg_ar_as_w1 \PWM1/dir_reg  (
    .clk(clk100m),
    .d(\PWM1/n32 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/dir_keep ));  // src/OnePWM.v(58)
  reg_sr_as_w1 \PWM1/pwm_reg  (
    .clk(clk100m),
    .d(\pwm[1]_d ),
    .en(1'b1),
    .reset(~\PWM1/u14_sel_is_1_o ),
    .set(1'b0),
    .q(\PWM1/pwm_keep ));  // src/OnePWM.v(45)
  reg_sr_as_w1 \PWM1/reg0_b0  (
    .clk(clk100m),
    .d(\PWM1/n13 [0]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [0]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b1  (
    .clk(clk100m),
    .d(\PWM1/n13 [1]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [1]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b10  (
    .clk(clk100m),
    .d(\PWM1/n13 [10]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [10]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b11  (
    .clk(clk100m),
    .d(\PWM1/n13 [11]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [11]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b12  (
    .clk(clk100m),
    .d(\PWM1/n13 [12]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [12]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b13  (
    .clk(clk100m),
    .d(\PWM1/n13 [13]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [13]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b14  (
    .clk(clk100m),
    .d(\PWM1/n13 [14]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [14]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b15  (
    .clk(clk100m),
    .d(\PWM1/n13 [15]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [15]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b16  (
    .clk(clk100m),
    .d(\PWM1/n13 [16]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [16]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b17  (
    .clk(clk100m),
    .d(\PWM1/n13 [17]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [17]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b18  (
    .clk(clk100m),
    .d(\PWM1/n13 [18]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [18]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b19  (
    .clk(clk100m),
    .d(\PWM1/n13 [19]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [19]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b2  (
    .clk(clk100m),
    .d(\PWM1/n13 [2]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [2]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b20  (
    .clk(clk100m),
    .d(\PWM1/n13 [20]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [20]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b21  (
    .clk(clk100m),
    .d(\PWM1/n13 [21]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [21]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b22  (
    .clk(clk100m),
    .d(\PWM1/n13 [22]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [22]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b23  (
    .clk(clk100m),
    .d(\PWM1/n13 [23]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [23]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b24  (
    .clk(clk100m),
    .d(\PWM1/n13 [24]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [24]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b25  (
    .clk(clk100m),
    .d(\PWM1/n13 [25]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [25]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b26  (
    .clk(clk100m),
    .d(\PWM1/n13 [26]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [26]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b3  (
    .clk(clk100m),
    .d(\PWM1/n13 [3]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [3]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b4  (
    .clk(clk100m),
    .d(\PWM1/n13 [4]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [4]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b5  (
    .clk(clk100m),
    .d(\PWM1/n13 [5]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [5]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b6  (
    .clk(clk100m),
    .d(\PWM1/n13 [6]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [6]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b7  (
    .clk(clk100m),
    .d(\PWM1/n13 [7]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [7]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b8  (
    .clk(clk100m),
    .d(\PWM1/n13 [8]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [8]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b9  (
    .clk(clk100m),
    .d(\PWM1/n13 [9]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b0  (
    .clk(clk100m),
    .d(freq1[0]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [0]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b1  (
    .clk(clk100m),
    .d(freq1[1]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [1]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b10  (
    .clk(clk100m),
    .d(freq1[10]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [10]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b11  (
    .clk(clk100m),
    .d(freq1[11]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [11]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b12  (
    .clk(clk100m),
    .d(freq1[12]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [12]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b13  (
    .clk(clk100m),
    .d(freq1[13]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [13]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b14  (
    .clk(clk100m),
    .d(freq1[14]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [14]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b15  (
    .clk(clk100m),
    .d(freq1[15]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [15]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b16  (
    .clk(clk100m),
    .d(freq1[16]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [16]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b17  (
    .clk(clk100m),
    .d(freq1[17]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [17]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b18  (
    .clk(clk100m),
    .d(freq1[18]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [18]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b19  (
    .clk(clk100m),
    .d(freq1[19]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [19]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b2  (
    .clk(clk100m),
    .d(freq1[2]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [2]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b20  (
    .clk(clk100m),
    .d(freq1[20]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [20]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b21  (
    .clk(clk100m),
    .d(freq1[21]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [21]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b22  (
    .clk(clk100m),
    .d(freq1[22]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [22]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b23  (
    .clk(clk100m),
    .d(freq1[23]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [23]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b24  (
    .clk(clk100m),
    .d(freq1[24]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [24]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b25  (
    .clk(clk100m),
    .d(freq1[25]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [25]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b26  (
    .clk(clk100m),
    .d(freq1[26]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [26]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b3  (
    .clk(clk100m),
    .d(freq1[3]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [3]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b4  (
    .clk(clk100m),
    .d(freq1[4]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [4]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b5  (
    .clk(clk100m),
    .d(freq1[5]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [5]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b6  (
    .clk(clk100m),
    .d(freq1[6]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [6]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b7  (
    .clk(clk100m),
    .d(freq1[7]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [7]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b8  (
    .clk(clk100m),
    .d(freq1[8]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [8]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b9  (
    .clk(clk100m),
    .d(freq1[9]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg2_b0  (
    .clk(clk100m),
    .d(\PWM1/n23 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[0]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b1  (
    .clk(clk100m),
    .d(\PWM1/n23 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[1]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b10  (
    .clk(clk100m),
    .d(\PWM1/n23 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[10]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b11  (
    .clk(clk100m),
    .d(\PWM1/n23 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[11]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b12  (
    .clk(clk100m),
    .d(\PWM1/n23 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[12]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b13  (
    .clk(clk100m),
    .d(\PWM1/n23 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[13]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b14  (
    .clk(clk100m),
    .d(\PWM1/n23 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[14]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b15  (
    .clk(clk100m),
    .d(\PWM1/n23 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[15]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b16  (
    .clk(clk100m),
    .d(\PWM1/n23 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[16]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b17  (
    .clk(clk100m),
    .d(\PWM1/n23 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[17]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b18  (
    .clk(clk100m),
    .d(\PWM1/n23 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[18]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b19  (
    .clk(clk100m),
    .d(\PWM1/n23 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[19]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b2  (
    .clk(clk100m),
    .d(\PWM1/n23 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[2]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b20  (
    .clk(clk100m),
    .d(\PWM1/n23 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[20]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b21  (
    .clk(clk100m),
    .d(\PWM1/n23 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[21]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b22  (
    .clk(clk100m),
    .d(\PWM1/n23 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[22]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b23  (
    .clk(clk100m),
    .d(\PWM1/n23 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[23]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b24  (
    .clk(clk100m),
    .d(\PWM1/n23 [24]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[24]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b25  (
    .clk(clk100m),
    .d(\PWM1/n23 [25]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[25]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b26  (
    .clk(clk100m),
    .d(\PWM1/n23 [26]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[26]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b27  (
    .clk(clk100m),
    .d(\PWM1/n23 [27]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[27]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b28  (
    .clk(clk100m),
    .d(\PWM1/n23 [28]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[28]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b29  (
    .clk(clk100m),
    .d(\PWM1/n23 [29]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[29]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b3  (
    .clk(clk100m),
    .d(\PWM1/n23 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[3]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b30  (
    .clk(clk100m),
    .d(\PWM1/n23 [30]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[30]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b31  (
    .clk(clk100m),
    .d(\PWM1/n23 [31]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[31]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b4  (
    .clk(clk100m),
    .d(\PWM1/n23 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[4]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b5  (
    .clk(clk100m),
    .d(\PWM1/n23 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[5]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b6  (
    .clk(clk100m),
    .d(\PWM1/n23 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[6]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b7  (
    .clk(clk100m),
    .d(\PWM1/n23 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[7]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b8  (
    .clk(clk100m),
    .d(\PWM1/n23 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[8]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b9  (
    .clk(clk100m),
    .d(\PWM1/n23 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[9]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg3_b0  (
    .clk(clk100m),
    .d(\PWM1/n31 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[0]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b1  (
    .clk(clk100m),
    .d(\PWM1/n31 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[1]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b10  (
    .clk(clk100m),
    .d(\PWM1/n31 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[10]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b11  (
    .clk(clk100m),
    .d(\PWM1/n31 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[11]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b12  (
    .clk(clk100m),
    .d(\PWM1/n31 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[12]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b13  (
    .clk(clk100m),
    .d(\PWM1/n31 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[13]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b14  (
    .clk(clk100m),
    .d(\PWM1/n31 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[14]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b15  (
    .clk(clk100m),
    .d(\PWM1/n31 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[15]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b16  (
    .clk(clk100m),
    .d(\PWM1/n31 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[16]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b17  (
    .clk(clk100m),
    .d(\PWM1/n31 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[17]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b18  (
    .clk(clk100m),
    .d(\PWM1/n31 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[18]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b19  (
    .clk(clk100m),
    .d(\PWM1/n31 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[19]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b2  (
    .clk(clk100m),
    .d(\PWM1/n31 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[2]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b20  (
    .clk(clk100m),
    .d(\PWM1/n31 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[20]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b21  (
    .clk(clk100m),
    .d(\PWM1/n31 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[21]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b22  (
    .clk(clk100m),
    .d(\PWM1/n31 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[22]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b23  (
    .clk(clk100m),
    .d(\PWM1/n31 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[23]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b3  (
    .clk(clk100m),
    .d(\PWM1/n31 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[3]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b4  (
    .clk(clk100m),
    .d(\PWM1/n31 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[4]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b5  (
    .clk(clk100m),
    .d(\PWM1/n31 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[5]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b6  (
    .clk(clk100m),
    .d(\PWM1/n31 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[6]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b7  (
    .clk(clk100m),
    .d(\PWM1/n31 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[7]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b8  (
    .clk(clk100m),
    .d(\PWM1/n31 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[8]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b9  (
    .clk(clk100m),
    .d(\PWM1/n31 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[9]_keep ));  // src/OnePWM.v(58)
  reg_ar_ss_w1 \PWM1/stopreq_reg  (
    .clk(clk100m),
    .d(\PWM1/n1 ),
    .en(1'b1),
    .reset(1'b0),
    .set(pwm_start_stop[1]),
    .q(\PWM1/stopreq_keep ));  // src/OnePWM.v(15)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub0/u0  (
    .a(\PWM1/FreCnt [0]),
    .b(1'b1),
    .c(\PWM1/sub0/c0 ),
    .o({\PWM1/sub0/c1 ,\PWM1/n12 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub0/u1  (
    .a(\PWM1/FreCnt [1]),
    .b(1'b0),
    .c(\PWM1/sub0/c1 ),
    .o({\PWM1/sub0/c2 ,\PWM1/n12 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub0/u10  (
    .a(\PWM1/FreCnt [10]),
    .b(1'b0),
    .c(\PWM1/sub0/c10 ),
    .o({\PWM1/sub0/c11 ,\PWM1/n12 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub0/u11  (
    .a(\PWM1/FreCnt [11]),
    .b(1'b0),
    .c(\PWM1/sub0/c11 ),
    .o({\PWM1/sub0/c12 ,\PWM1/n12 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub0/u12  (
    .a(\PWM1/FreCnt [12]),
    .b(1'b0),
    .c(\PWM1/sub0/c12 ),
    .o({\PWM1/sub0/c13 ,\PWM1/n12 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub0/u13  (
    .a(\PWM1/FreCnt [13]),
    .b(1'b0),
    .c(\PWM1/sub0/c13 ),
    .o({\PWM1/sub0/c14 ,\PWM1/n12 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub0/u14  (
    .a(\PWM1/FreCnt [14]),
    .b(1'b0),
    .c(\PWM1/sub0/c14 ),
    .o({\PWM1/sub0/c15 ,\PWM1/n12 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub0/u15  (
    .a(\PWM1/FreCnt [15]),
    .b(1'b0),
    .c(\PWM1/sub0/c15 ),
    .o({\PWM1/sub0/c16 ,\PWM1/n12 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub0/u16  (
    .a(\PWM1/FreCnt [16]),
    .b(1'b0),
    .c(\PWM1/sub0/c16 ),
    .o({\PWM1/sub0/c17 ,\PWM1/n12 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub0/u17  (
    .a(\PWM1/FreCnt [17]),
    .b(1'b0),
    .c(\PWM1/sub0/c17 ),
    .o({\PWM1/sub0/c18 ,\PWM1/n12 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub0/u18  (
    .a(\PWM1/FreCnt [18]),
    .b(1'b0),
    .c(\PWM1/sub0/c18 ),
    .o({\PWM1/sub0/c19 ,\PWM1/n12 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub0/u19  (
    .a(\PWM1/FreCnt [19]),
    .b(1'b0),
    .c(\PWM1/sub0/c19 ),
    .o({\PWM1/sub0/c20 ,\PWM1/n12 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub0/u2  (
    .a(\PWM1/FreCnt [2]),
    .b(1'b0),
    .c(\PWM1/sub0/c2 ),
    .o({\PWM1/sub0/c3 ,\PWM1/n12 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub0/u20  (
    .a(\PWM1/FreCnt [20]),
    .b(1'b0),
    .c(\PWM1/sub0/c20 ),
    .o({\PWM1/sub0/c21 ,\PWM1/n12 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub0/u21  (
    .a(\PWM1/FreCnt [21]),
    .b(1'b0),
    .c(\PWM1/sub0/c21 ),
    .o({\PWM1/sub0/c22 ,\PWM1/n12 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub0/u22  (
    .a(\PWM1/FreCnt [22]),
    .b(1'b0),
    .c(\PWM1/sub0/c22 ),
    .o({\PWM1/sub0/c23 ,\PWM1/n12 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub0/u23  (
    .a(\PWM1/FreCnt [23]),
    .b(1'b0),
    .c(\PWM1/sub0/c23 ),
    .o({\PWM1/sub0/c24 ,\PWM1/n12 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub0/u24  (
    .a(\PWM1/FreCnt [24]),
    .b(1'b0),
    .c(\PWM1/sub0/c24 ),
    .o({\PWM1/sub0/c25 ,\PWM1/n12 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub0/u25  (
    .a(\PWM1/FreCnt [25]),
    .b(1'b0),
    .c(\PWM1/sub0/c25 ),
    .o({\PWM1/sub0/c26 ,\PWM1/n12 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub0/u26  (
    .a(\PWM1/FreCnt [26]),
    .b(1'b0),
    .c(\PWM1/sub0/c26 ),
    .o({open_n8,\PWM1/n12 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub0/u3  (
    .a(\PWM1/FreCnt [3]),
    .b(1'b0),
    .c(\PWM1/sub0/c3 ),
    .o({\PWM1/sub0/c4 ,\PWM1/n12 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub0/u4  (
    .a(\PWM1/FreCnt [4]),
    .b(1'b0),
    .c(\PWM1/sub0/c4 ),
    .o({\PWM1/sub0/c5 ,\PWM1/n12 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub0/u5  (
    .a(\PWM1/FreCnt [5]),
    .b(1'b0),
    .c(\PWM1/sub0/c5 ),
    .o({\PWM1/sub0/c6 ,\PWM1/n12 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub0/u6  (
    .a(\PWM1/FreCnt [6]),
    .b(1'b0),
    .c(\PWM1/sub0/c6 ),
    .o({\PWM1/sub0/c7 ,\PWM1/n12 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub0/u7  (
    .a(\PWM1/FreCnt [7]),
    .b(1'b0),
    .c(\PWM1/sub0/c7 ),
    .o({\PWM1/sub0/c8 ,\PWM1/n12 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub0/u8  (
    .a(\PWM1/FreCnt [8]),
    .b(1'b0),
    .c(\PWM1/sub0/c8 ),
    .o({\PWM1/sub0/c9 ,\PWM1/n12 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub0/u9  (
    .a(\PWM1/FreCnt [9]),
    .b(1'b0),
    .c(\PWM1/sub0/c9 ),
    .o({\PWM1/sub0/c10 ,\PWM1/n12 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \PWM1/sub0/ucin  (
    .a(1'b0),
    .o({\PWM1/sub0/c0 ,open_n11}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub1/u0  (
    .a(pnumcnt1[0]),
    .b(1'b1),
    .c(\PWM1/sub1/c0 ),
    .o({\PWM1/sub1/c1 ,\PWM1/n26 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub1/u1  (
    .a(pnumcnt1[1]),
    .b(1'b0),
    .c(\PWM1/sub1/c1 ),
    .o({\PWM1/sub1/c2 ,\PWM1/n26 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub1/u10  (
    .a(pnumcnt1[10]),
    .b(1'b0),
    .c(\PWM1/sub1/c10 ),
    .o({\PWM1/sub1/c11 ,\PWM1/n26 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub1/u11  (
    .a(pnumcnt1[11]),
    .b(1'b0),
    .c(\PWM1/sub1/c11 ),
    .o({\PWM1/sub1/c12 ,\PWM1/n26 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub1/u12  (
    .a(pnumcnt1[12]),
    .b(1'b0),
    .c(\PWM1/sub1/c12 ),
    .o({\PWM1/sub1/c13 ,\PWM1/n26 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub1/u13  (
    .a(pnumcnt1[13]),
    .b(1'b0),
    .c(\PWM1/sub1/c13 ),
    .o({\PWM1/sub1/c14 ,\PWM1/n26 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub1/u14  (
    .a(pnumcnt1[14]),
    .b(1'b0),
    .c(\PWM1/sub1/c14 ),
    .o({\PWM1/sub1/c15 ,\PWM1/n26 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub1/u15  (
    .a(pnumcnt1[15]),
    .b(1'b0),
    .c(\PWM1/sub1/c15 ),
    .o({\PWM1/sub1/c16 ,\PWM1/n26 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub1/u16  (
    .a(pnumcnt1[16]),
    .b(1'b0),
    .c(\PWM1/sub1/c16 ),
    .o({\PWM1/sub1/c17 ,\PWM1/n26 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub1/u17  (
    .a(pnumcnt1[17]),
    .b(1'b0),
    .c(\PWM1/sub1/c17 ),
    .o({\PWM1/sub1/c18 ,\PWM1/n26 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub1/u18  (
    .a(pnumcnt1[18]),
    .b(1'b0),
    .c(\PWM1/sub1/c18 ),
    .o({\PWM1/sub1/c19 ,\PWM1/n26 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub1/u19  (
    .a(pnumcnt1[19]),
    .b(1'b0),
    .c(\PWM1/sub1/c19 ),
    .o({\PWM1/sub1/c20 ,\PWM1/n26 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub1/u2  (
    .a(pnumcnt1[2]),
    .b(1'b0),
    .c(\PWM1/sub1/c2 ),
    .o({\PWM1/sub1/c3 ,\PWM1/n26 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub1/u20  (
    .a(pnumcnt1[20]),
    .b(1'b0),
    .c(\PWM1/sub1/c20 ),
    .o({\PWM1/sub1/c21 ,\PWM1/n26 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub1/u21  (
    .a(pnumcnt1[21]),
    .b(1'b0),
    .c(\PWM1/sub1/c21 ),
    .o({\PWM1/sub1/c22 ,\PWM1/n26 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub1/u22  (
    .a(pnumcnt1[22]),
    .b(1'b0),
    .c(\PWM1/sub1/c22 ),
    .o({\PWM1/sub1/c23 ,\PWM1/n26 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub1/u23  (
    .a(pnumcnt1[23]),
    .b(1'b0),
    .c(\PWM1/sub1/c23 ),
    .o({open_n12,\PWM1/n26 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub1/u3  (
    .a(pnumcnt1[3]),
    .b(1'b0),
    .c(\PWM1/sub1/c3 ),
    .o({\PWM1/sub1/c4 ,\PWM1/n26 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub1/u4  (
    .a(pnumcnt1[4]),
    .b(1'b0),
    .c(\PWM1/sub1/c4 ),
    .o({\PWM1/sub1/c5 ,\PWM1/n26 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub1/u5  (
    .a(pnumcnt1[5]),
    .b(1'b0),
    .c(\PWM1/sub1/c5 ),
    .o({\PWM1/sub1/c6 ,\PWM1/n26 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub1/u6  (
    .a(pnumcnt1[6]),
    .b(1'b0),
    .c(\PWM1/sub1/c6 ),
    .o({\PWM1/sub1/c7 ,\PWM1/n26 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub1/u7  (
    .a(pnumcnt1[7]),
    .b(1'b0),
    .c(\PWM1/sub1/c7 ),
    .o({\PWM1/sub1/c8 ,\PWM1/n26 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub1/u8  (
    .a(pnumcnt1[8]),
    .b(1'b0),
    .c(\PWM1/sub1/c8 ),
    .o({\PWM1/sub1/c9 ,\PWM1/n26 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM1/sub1/u9  (
    .a(pnumcnt1[9]),
    .b(1'b0),
    .c(\PWM1/sub1/c9 ),
    .o({\PWM1/sub1/c10 ,\PWM1/n26 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \PWM1/sub1/ucin  (
    .a(1'b0),
    .o({\PWM1/sub1/c0 ,open_n15}));
  reg_ar_as_w1 \PWM2/State_reg  (
    .clk(clk100m),
    .d(\PWM2/n10 ),
    .en(1'b1),
    .reset(~rstn),
    .set(1'b0),
    .q(pwm_state_read[2]));  // src/OnePWM.v(26)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[0]  (
    .i(\PWM2/RemaTxNum[0]_keep ),
    .o(pnumcnt2[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[10]  (
    .i(\PWM2/RemaTxNum[10]_keep ),
    .o(pnumcnt2[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[11]  (
    .i(\PWM2/RemaTxNum[11]_keep ),
    .o(pnumcnt2[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[12]  (
    .i(\PWM2/RemaTxNum[12]_keep ),
    .o(pnumcnt2[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[13]  (
    .i(\PWM2/RemaTxNum[13]_keep ),
    .o(pnumcnt2[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[14]  (
    .i(\PWM2/RemaTxNum[14]_keep ),
    .o(pnumcnt2[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[15]  (
    .i(\PWM2/RemaTxNum[15]_keep ),
    .o(pnumcnt2[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[16]  (
    .i(\PWM2/RemaTxNum[16]_keep ),
    .o(pnumcnt2[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[17]  (
    .i(\PWM2/RemaTxNum[17]_keep ),
    .o(pnumcnt2[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[18]  (
    .i(\PWM2/RemaTxNum[18]_keep ),
    .o(pnumcnt2[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[19]  (
    .i(\PWM2/RemaTxNum[19]_keep ),
    .o(pnumcnt2[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[1]  (
    .i(\PWM2/RemaTxNum[1]_keep ),
    .o(pnumcnt2[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[20]  (
    .i(\PWM2/RemaTxNum[20]_keep ),
    .o(pnumcnt2[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[21]  (
    .i(\PWM2/RemaTxNum[21]_keep ),
    .o(pnumcnt2[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[22]  (
    .i(\PWM2/RemaTxNum[22]_keep ),
    .o(pnumcnt2[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[23]  (
    .i(\PWM2/RemaTxNum[23]_keep ),
    .o(pnumcnt2[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[2]  (
    .i(\PWM2/RemaTxNum[2]_keep ),
    .o(pnumcnt2[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[3]  (
    .i(\PWM2/RemaTxNum[3]_keep ),
    .o(pnumcnt2[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[4]  (
    .i(\PWM2/RemaTxNum[4]_keep ),
    .o(pnumcnt2[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[5]  (
    .i(\PWM2/RemaTxNum[5]_keep ),
    .o(pnumcnt2[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[6]  (
    .i(\PWM2/RemaTxNum[6]_keep ),
    .o(pnumcnt2[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[7]  (
    .i(\PWM2/RemaTxNum[7]_keep ),
    .o(pnumcnt2[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[8]  (
    .i(\PWM2/RemaTxNum[8]_keep ),
    .o(pnumcnt2[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[9]  (
    .i(\PWM2/RemaTxNum[9]_keep ),
    .o(pnumcnt2[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_dir  (
    .i(\PWM2/dir_keep ),
    .o(dir_pad[2]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[0]  (
    .i(\PWM2/pnumr[0]_keep ),
    .o(\PWM2/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[10]  (
    .i(\PWM2/pnumr[10]_keep ),
    .o(\PWM2/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[11]  (
    .i(\PWM2/pnumr[11]_keep ),
    .o(\PWM2/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[12]  (
    .i(\PWM2/pnumr[12]_keep ),
    .o(\PWM2/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[13]  (
    .i(\PWM2/pnumr[13]_keep ),
    .o(\PWM2/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[14]  (
    .i(\PWM2/pnumr[14]_keep ),
    .o(\PWM2/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[15]  (
    .i(\PWM2/pnumr[15]_keep ),
    .o(\PWM2/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[16]  (
    .i(\PWM2/pnumr[16]_keep ),
    .o(\PWM2/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[17]  (
    .i(\PWM2/pnumr[17]_keep ),
    .o(\PWM2/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[18]  (
    .i(\PWM2/pnumr[18]_keep ),
    .o(\PWM2/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[19]  (
    .i(\PWM2/pnumr[19]_keep ),
    .o(\PWM2/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[1]  (
    .i(\PWM2/pnumr[1]_keep ),
    .o(\PWM2/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[20]  (
    .i(\PWM2/pnumr[20]_keep ),
    .o(\PWM2/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[21]  (
    .i(\PWM2/pnumr[21]_keep ),
    .o(\PWM2/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[22]  (
    .i(\PWM2/pnumr[22]_keep ),
    .o(\PWM2/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[23]  (
    .i(\PWM2/pnumr[23]_keep ),
    .o(\PWM2/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[24]  (
    .i(\PWM2/pnumr[24]_keep ),
    .o(\PWM2/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[25]  (
    .i(\PWM2/pnumr[25]_keep ),
    .o(\PWM2/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[26]  (
    .i(\PWM2/pnumr[26]_keep ),
    .o(\PWM2/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[27]  (
    .i(\PWM2/pnumr[27]_keep ),
    .o(\PWM2/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[28]  (
    .i(\PWM2/pnumr[28]_keep ),
    .o(\PWM2/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[29]  (
    .i(\PWM2/pnumr[29]_keep ),
    .o(\PWM2/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[2]  (
    .i(\PWM2/pnumr[2]_keep ),
    .o(\PWM2/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[30]  (
    .i(\PWM2/pnumr[30]_keep ),
    .o(\PWM2/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[31]  (
    .i(\PWM2/pnumr[31]_keep ),
    .o(\PWM2/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[3]  (
    .i(\PWM2/pnumr[3]_keep ),
    .o(\PWM2/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[4]  (
    .i(\PWM2/pnumr[4]_keep ),
    .o(\PWM2/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[5]  (
    .i(\PWM2/pnumr[5]_keep ),
    .o(\PWM2/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[6]  (
    .i(\PWM2/pnumr[6]_keep ),
    .o(\PWM2/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[7]  (
    .i(\PWM2/pnumr[7]_keep ),
    .o(\PWM2/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[8]  (
    .i(\PWM2/pnumr[8]_keep ),
    .o(\PWM2/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[9]  (
    .i(\PWM2/pnumr[9]_keep ),
    .o(\PWM2/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pwm  (
    .i(\PWM2/pwm_keep ),
    .o(pwm_pad[2]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_stopreq  (
    .i(\PWM2/stopreq_keep ),
    .o(\PWM2/stopreq ));  // src/OnePWM.v(14)
  reg_ar_as_w1 \PWM2/dir_reg  (
    .clk(clk100m),
    .d(\PWM2/n32 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/dir_keep ));  // src/OnePWM.v(58)
  reg_sr_as_w1 \PWM2/pwm_reg  (
    .clk(clk100m),
    .d(\pwm[2]_d ),
    .en(1'b1),
    .reset(~\PWM2/u14_sel_is_1_o ),
    .set(1'b0),
    .q(\PWM2/pwm_keep ));  // src/OnePWM.v(45)
  reg_sr_as_w1 \PWM2/reg0_b0  (
    .clk(clk100m),
    .d(\PWM2/n13 [0]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [0]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b1  (
    .clk(clk100m),
    .d(\PWM2/n13 [1]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [1]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b10  (
    .clk(clk100m),
    .d(\PWM2/n13 [10]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [10]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b11  (
    .clk(clk100m),
    .d(\PWM2/n13 [11]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [11]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b12  (
    .clk(clk100m),
    .d(\PWM2/n13 [12]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [12]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b13  (
    .clk(clk100m),
    .d(\PWM2/n13 [13]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [13]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b14  (
    .clk(clk100m),
    .d(\PWM2/n13 [14]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [14]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b15  (
    .clk(clk100m),
    .d(\PWM2/n13 [15]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [15]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b16  (
    .clk(clk100m),
    .d(\PWM2/n13 [16]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [16]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b17  (
    .clk(clk100m),
    .d(\PWM2/n13 [17]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [17]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b18  (
    .clk(clk100m),
    .d(\PWM2/n13 [18]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [18]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b19  (
    .clk(clk100m),
    .d(\PWM2/n13 [19]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [19]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b2  (
    .clk(clk100m),
    .d(\PWM2/n13 [2]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [2]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b20  (
    .clk(clk100m),
    .d(\PWM2/n13 [20]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [20]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b21  (
    .clk(clk100m),
    .d(\PWM2/n13 [21]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [21]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b22  (
    .clk(clk100m),
    .d(\PWM2/n13 [22]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [22]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b23  (
    .clk(clk100m),
    .d(\PWM2/n13 [23]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [23]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b24  (
    .clk(clk100m),
    .d(\PWM2/n13 [24]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [24]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b25  (
    .clk(clk100m),
    .d(\PWM2/n13 [25]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [25]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b26  (
    .clk(clk100m),
    .d(\PWM2/n13 [26]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [26]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b3  (
    .clk(clk100m),
    .d(\PWM2/n13 [3]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [3]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b4  (
    .clk(clk100m),
    .d(\PWM2/n13 [4]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [4]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b5  (
    .clk(clk100m),
    .d(\PWM2/n13 [5]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [5]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b6  (
    .clk(clk100m),
    .d(\PWM2/n13 [6]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [6]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b7  (
    .clk(clk100m),
    .d(\PWM2/n13 [7]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [7]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b8  (
    .clk(clk100m),
    .d(\PWM2/n13 [8]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [8]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b9  (
    .clk(clk100m),
    .d(\PWM2/n13 [9]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b0  (
    .clk(clk100m),
    .d(freq2[0]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [0]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b1  (
    .clk(clk100m),
    .d(freq2[1]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [1]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b10  (
    .clk(clk100m),
    .d(freq2[10]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [10]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b11  (
    .clk(clk100m),
    .d(freq2[11]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [11]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b12  (
    .clk(clk100m),
    .d(freq2[12]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [12]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b13  (
    .clk(clk100m),
    .d(freq2[13]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [13]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b14  (
    .clk(clk100m),
    .d(freq2[14]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [14]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b15  (
    .clk(clk100m),
    .d(freq2[15]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [15]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b16  (
    .clk(clk100m),
    .d(freq2[16]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [16]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b17  (
    .clk(clk100m),
    .d(freq2[17]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [17]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b18  (
    .clk(clk100m),
    .d(freq2[18]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [18]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b19  (
    .clk(clk100m),
    .d(freq2[19]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [19]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b2  (
    .clk(clk100m),
    .d(freq2[2]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [2]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b20  (
    .clk(clk100m),
    .d(freq2[20]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [20]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b21  (
    .clk(clk100m),
    .d(freq2[21]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [21]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b22  (
    .clk(clk100m),
    .d(freq2[22]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [22]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b23  (
    .clk(clk100m),
    .d(freq2[23]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [23]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b24  (
    .clk(clk100m),
    .d(freq2[24]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [24]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b25  (
    .clk(clk100m),
    .d(freq2[25]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [25]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b26  (
    .clk(clk100m),
    .d(freq2[26]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [26]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b3  (
    .clk(clk100m),
    .d(freq2[3]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [3]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b4  (
    .clk(clk100m),
    .d(freq2[4]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [4]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b5  (
    .clk(clk100m),
    .d(freq2[5]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [5]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b6  (
    .clk(clk100m),
    .d(freq2[6]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [6]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b7  (
    .clk(clk100m),
    .d(freq2[7]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [7]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b8  (
    .clk(clk100m),
    .d(freq2[8]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [8]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b9  (
    .clk(clk100m),
    .d(freq2[9]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg2_b0  (
    .clk(clk100m),
    .d(\PWM2/n23 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[0]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b1  (
    .clk(clk100m),
    .d(\PWM2/n23 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[1]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b10  (
    .clk(clk100m),
    .d(\PWM2/n23 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[10]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b11  (
    .clk(clk100m),
    .d(\PWM2/n23 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[11]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b12  (
    .clk(clk100m),
    .d(\PWM2/n23 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[12]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b13  (
    .clk(clk100m),
    .d(\PWM2/n23 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[13]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b14  (
    .clk(clk100m),
    .d(\PWM2/n23 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[14]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b15  (
    .clk(clk100m),
    .d(\PWM2/n23 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[15]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b16  (
    .clk(clk100m),
    .d(\PWM2/n23 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[16]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b17  (
    .clk(clk100m),
    .d(\PWM2/n23 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[17]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b18  (
    .clk(clk100m),
    .d(\PWM2/n23 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[18]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b19  (
    .clk(clk100m),
    .d(\PWM2/n23 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[19]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b2  (
    .clk(clk100m),
    .d(\PWM2/n23 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[2]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b20  (
    .clk(clk100m),
    .d(\PWM2/n23 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[20]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b21  (
    .clk(clk100m),
    .d(\PWM2/n23 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[21]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b22  (
    .clk(clk100m),
    .d(\PWM2/n23 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[22]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b23  (
    .clk(clk100m),
    .d(\PWM2/n23 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[23]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b24  (
    .clk(clk100m),
    .d(\PWM2/n23 [24]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[24]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b25  (
    .clk(clk100m),
    .d(\PWM2/n23 [25]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[25]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b26  (
    .clk(clk100m),
    .d(\PWM2/n23 [26]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[26]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b27  (
    .clk(clk100m),
    .d(\PWM2/n23 [27]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[27]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b28  (
    .clk(clk100m),
    .d(\PWM2/n23 [28]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[28]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b29  (
    .clk(clk100m),
    .d(\PWM2/n23 [29]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[29]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b3  (
    .clk(clk100m),
    .d(\PWM2/n23 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[3]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b30  (
    .clk(clk100m),
    .d(\PWM2/n23 [30]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[30]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b31  (
    .clk(clk100m),
    .d(\PWM2/n23 [31]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[31]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b4  (
    .clk(clk100m),
    .d(\PWM2/n23 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[4]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b5  (
    .clk(clk100m),
    .d(\PWM2/n23 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[5]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b6  (
    .clk(clk100m),
    .d(\PWM2/n23 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[6]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b7  (
    .clk(clk100m),
    .d(\PWM2/n23 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[7]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b8  (
    .clk(clk100m),
    .d(\PWM2/n23 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[8]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b9  (
    .clk(clk100m),
    .d(\PWM2/n23 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[9]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg3_b0  (
    .clk(clk100m),
    .d(\PWM2/n31 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[0]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b1  (
    .clk(clk100m),
    .d(\PWM2/n31 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[1]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b10  (
    .clk(clk100m),
    .d(\PWM2/n31 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[10]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b11  (
    .clk(clk100m),
    .d(\PWM2/n31 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[11]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b12  (
    .clk(clk100m),
    .d(\PWM2/n31 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[12]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b13  (
    .clk(clk100m),
    .d(\PWM2/n31 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[13]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b14  (
    .clk(clk100m),
    .d(\PWM2/n31 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[14]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b15  (
    .clk(clk100m),
    .d(\PWM2/n31 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[15]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b16  (
    .clk(clk100m),
    .d(\PWM2/n31 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[16]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b17  (
    .clk(clk100m),
    .d(\PWM2/n31 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[17]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b18  (
    .clk(clk100m),
    .d(\PWM2/n31 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[18]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b19  (
    .clk(clk100m),
    .d(\PWM2/n31 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[19]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b2  (
    .clk(clk100m),
    .d(\PWM2/n31 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[2]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b20  (
    .clk(clk100m),
    .d(\PWM2/n31 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[20]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b21  (
    .clk(clk100m),
    .d(\PWM2/n31 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[21]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b22  (
    .clk(clk100m),
    .d(\PWM2/n31 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[22]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b23  (
    .clk(clk100m),
    .d(\PWM2/n31 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[23]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b3  (
    .clk(clk100m),
    .d(\PWM2/n31 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[3]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b4  (
    .clk(clk100m),
    .d(\PWM2/n31 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[4]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b5  (
    .clk(clk100m),
    .d(\PWM2/n31 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[5]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b6  (
    .clk(clk100m),
    .d(\PWM2/n31 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[6]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b7  (
    .clk(clk100m),
    .d(\PWM2/n31 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[7]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b8  (
    .clk(clk100m),
    .d(\PWM2/n31 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[8]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b9  (
    .clk(clk100m),
    .d(\PWM2/n31 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[9]_keep ));  // src/OnePWM.v(58)
  reg_ar_ss_w1 \PWM2/stopreq_reg  (
    .clk(clk100m),
    .d(\PWM2/n1 ),
    .en(1'b1),
    .reset(1'b0),
    .set(pwm_start_stop[2]),
    .q(\PWM2/stopreq_keep ));  // src/OnePWM.v(15)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub0/u0  (
    .a(\PWM2/FreCnt [0]),
    .b(1'b1),
    .c(\PWM2/sub0/c0 ),
    .o({\PWM2/sub0/c1 ,\PWM2/n12 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub0/u1  (
    .a(\PWM2/FreCnt [1]),
    .b(1'b0),
    .c(\PWM2/sub0/c1 ),
    .o({\PWM2/sub0/c2 ,\PWM2/n12 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub0/u10  (
    .a(\PWM2/FreCnt [10]),
    .b(1'b0),
    .c(\PWM2/sub0/c10 ),
    .o({\PWM2/sub0/c11 ,\PWM2/n12 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub0/u11  (
    .a(\PWM2/FreCnt [11]),
    .b(1'b0),
    .c(\PWM2/sub0/c11 ),
    .o({\PWM2/sub0/c12 ,\PWM2/n12 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub0/u12  (
    .a(\PWM2/FreCnt [12]),
    .b(1'b0),
    .c(\PWM2/sub0/c12 ),
    .o({\PWM2/sub0/c13 ,\PWM2/n12 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub0/u13  (
    .a(\PWM2/FreCnt [13]),
    .b(1'b0),
    .c(\PWM2/sub0/c13 ),
    .o({\PWM2/sub0/c14 ,\PWM2/n12 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub0/u14  (
    .a(\PWM2/FreCnt [14]),
    .b(1'b0),
    .c(\PWM2/sub0/c14 ),
    .o({\PWM2/sub0/c15 ,\PWM2/n12 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub0/u15  (
    .a(\PWM2/FreCnt [15]),
    .b(1'b0),
    .c(\PWM2/sub0/c15 ),
    .o({\PWM2/sub0/c16 ,\PWM2/n12 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub0/u16  (
    .a(\PWM2/FreCnt [16]),
    .b(1'b0),
    .c(\PWM2/sub0/c16 ),
    .o({\PWM2/sub0/c17 ,\PWM2/n12 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub0/u17  (
    .a(\PWM2/FreCnt [17]),
    .b(1'b0),
    .c(\PWM2/sub0/c17 ),
    .o({\PWM2/sub0/c18 ,\PWM2/n12 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub0/u18  (
    .a(\PWM2/FreCnt [18]),
    .b(1'b0),
    .c(\PWM2/sub0/c18 ),
    .o({\PWM2/sub0/c19 ,\PWM2/n12 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub0/u19  (
    .a(\PWM2/FreCnt [19]),
    .b(1'b0),
    .c(\PWM2/sub0/c19 ),
    .o({\PWM2/sub0/c20 ,\PWM2/n12 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub0/u2  (
    .a(\PWM2/FreCnt [2]),
    .b(1'b0),
    .c(\PWM2/sub0/c2 ),
    .o({\PWM2/sub0/c3 ,\PWM2/n12 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub0/u20  (
    .a(\PWM2/FreCnt [20]),
    .b(1'b0),
    .c(\PWM2/sub0/c20 ),
    .o({\PWM2/sub0/c21 ,\PWM2/n12 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub0/u21  (
    .a(\PWM2/FreCnt [21]),
    .b(1'b0),
    .c(\PWM2/sub0/c21 ),
    .o({\PWM2/sub0/c22 ,\PWM2/n12 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub0/u22  (
    .a(\PWM2/FreCnt [22]),
    .b(1'b0),
    .c(\PWM2/sub0/c22 ),
    .o({\PWM2/sub0/c23 ,\PWM2/n12 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub0/u23  (
    .a(\PWM2/FreCnt [23]),
    .b(1'b0),
    .c(\PWM2/sub0/c23 ),
    .o({\PWM2/sub0/c24 ,\PWM2/n12 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub0/u24  (
    .a(\PWM2/FreCnt [24]),
    .b(1'b0),
    .c(\PWM2/sub0/c24 ),
    .o({\PWM2/sub0/c25 ,\PWM2/n12 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub0/u25  (
    .a(\PWM2/FreCnt [25]),
    .b(1'b0),
    .c(\PWM2/sub0/c25 ),
    .o({\PWM2/sub0/c26 ,\PWM2/n12 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub0/u26  (
    .a(\PWM2/FreCnt [26]),
    .b(1'b0),
    .c(\PWM2/sub0/c26 ),
    .o({open_n16,\PWM2/n12 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub0/u3  (
    .a(\PWM2/FreCnt [3]),
    .b(1'b0),
    .c(\PWM2/sub0/c3 ),
    .o({\PWM2/sub0/c4 ,\PWM2/n12 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub0/u4  (
    .a(\PWM2/FreCnt [4]),
    .b(1'b0),
    .c(\PWM2/sub0/c4 ),
    .o({\PWM2/sub0/c5 ,\PWM2/n12 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub0/u5  (
    .a(\PWM2/FreCnt [5]),
    .b(1'b0),
    .c(\PWM2/sub0/c5 ),
    .o({\PWM2/sub0/c6 ,\PWM2/n12 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub0/u6  (
    .a(\PWM2/FreCnt [6]),
    .b(1'b0),
    .c(\PWM2/sub0/c6 ),
    .o({\PWM2/sub0/c7 ,\PWM2/n12 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub0/u7  (
    .a(\PWM2/FreCnt [7]),
    .b(1'b0),
    .c(\PWM2/sub0/c7 ),
    .o({\PWM2/sub0/c8 ,\PWM2/n12 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub0/u8  (
    .a(\PWM2/FreCnt [8]),
    .b(1'b0),
    .c(\PWM2/sub0/c8 ),
    .o({\PWM2/sub0/c9 ,\PWM2/n12 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub0/u9  (
    .a(\PWM2/FreCnt [9]),
    .b(1'b0),
    .c(\PWM2/sub0/c9 ),
    .o({\PWM2/sub0/c10 ,\PWM2/n12 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \PWM2/sub0/ucin  (
    .a(1'b0),
    .o({\PWM2/sub0/c0 ,open_n19}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub1/u0  (
    .a(pnumcnt2[0]),
    .b(1'b1),
    .c(\PWM2/sub1/c0 ),
    .o({\PWM2/sub1/c1 ,\PWM2/n26 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub1/u1  (
    .a(pnumcnt2[1]),
    .b(1'b0),
    .c(\PWM2/sub1/c1 ),
    .o({\PWM2/sub1/c2 ,\PWM2/n26 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub1/u10  (
    .a(pnumcnt2[10]),
    .b(1'b0),
    .c(\PWM2/sub1/c10 ),
    .o({\PWM2/sub1/c11 ,\PWM2/n26 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub1/u11  (
    .a(pnumcnt2[11]),
    .b(1'b0),
    .c(\PWM2/sub1/c11 ),
    .o({\PWM2/sub1/c12 ,\PWM2/n26 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub1/u12  (
    .a(pnumcnt2[12]),
    .b(1'b0),
    .c(\PWM2/sub1/c12 ),
    .o({\PWM2/sub1/c13 ,\PWM2/n26 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub1/u13  (
    .a(pnumcnt2[13]),
    .b(1'b0),
    .c(\PWM2/sub1/c13 ),
    .o({\PWM2/sub1/c14 ,\PWM2/n26 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub1/u14  (
    .a(pnumcnt2[14]),
    .b(1'b0),
    .c(\PWM2/sub1/c14 ),
    .o({\PWM2/sub1/c15 ,\PWM2/n26 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub1/u15  (
    .a(pnumcnt2[15]),
    .b(1'b0),
    .c(\PWM2/sub1/c15 ),
    .o({\PWM2/sub1/c16 ,\PWM2/n26 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub1/u16  (
    .a(pnumcnt2[16]),
    .b(1'b0),
    .c(\PWM2/sub1/c16 ),
    .o({\PWM2/sub1/c17 ,\PWM2/n26 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub1/u17  (
    .a(pnumcnt2[17]),
    .b(1'b0),
    .c(\PWM2/sub1/c17 ),
    .o({\PWM2/sub1/c18 ,\PWM2/n26 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub1/u18  (
    .a(pnumcnt2[18]),
    .b(1'b0),
    .c(\PWM2/sub1/c18 ),
    .o({\PWM2/sub1/c19 ,\PWM2/n26 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub1/u19  (
    .a(pnumcnt2[19]),
    .b(1'b0),
    .c(\PWM2/sub1/c19 ),
    .o({\PWM2/sub1/c20 ,\PWM2/n26 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub1/u2  (
    .a(pnumcnt2[2]),
    .b(1'b0),
    .c(\PWM2/sub1/c2 ),
    .o({\PWM2/sub1/c3 ,\PWM2/n26 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub1/u20  (
    .a(pnumcnt2[20]),
    .b(1'b0),
    .c(\PWM2/sub1/c20 ),
    .o({\PWM2/sub1/c21 ,\PWM2/n26 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub1/u21  (
    .a(pnumcnt2[21]),
    .b(1'b0),
    .c(\PWM2/sub1/c21 ),
    .o({\PWM2/sub1/c22 ,\PWM2/n26 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub1/u22  (
    .a(pnumcnt2[22]),
    .b(1'b0),
    .c(\PWM2/sub1/c22 ),
    .o({\PWM2/sub1/c23 ,\PWM2/n26 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub1/u23  (
    .a(pnumcnt2[23]),
    .b(1'b0),
    .c(\PWM2/sub1/c23 ),
    .o({open_n20,\PWM2/n26 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub1/u3  (
    .a(pnumcnt2[3]),
    .b(1'b0),
    .c(\PWM2/sub1/c3 ),
    .o({\PWM2/sub1/c4 ,\PWM2/n26 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub1/u4  (
    .a(pnumcnt2[4]),
    .b(1'b0),
    .c(\PWM2/sub1/c4 ),
    .o({\PWM2/sub1/c5 ,\PWM2/n26 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub1/u5  (
    .a(pnumcnt2[5]),
    .b(1'b0),
    .c(\PWM2/sub1/c5 ),
    .o({\PWM2/sub1/c6 ,\PWM2/n26 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub1/u6  (
    .a(pnumcnt2[6]),
    .b(1'b0),
    .c(\PWM2/sub1/c6 ),
    .o({\PWM2/sub1/c7 ,\PWM2/n26 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub1/u7  (
    .a(pnumcnt2[7]),
    .b(1'b0),
    .c(\PWM2/sub1/c7 ),
    .o({\PWM2/sub1/c8 ,\PWM2/n26 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub1/u8  (
    .a(pnumcnt2[8]),
    .b(1'b0),
    .c(\PWM2/sub1/c8 ),
    .o({\PWM2/sub1/c9 ,\PWM2/n26 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM2/sub1/u9  (
    .a(pnumcnt2[9]),
    .b(1'b0),
    .c(\PWM2/sub1/c9 ),
    .o({\PWM2/sub1/c10 ,\PWM2/n26 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \PWM2/sub1/ucin  (
    .a(1'b0),
    .o({\PWM2/sub1/c0 ,open_n23}));
  reg_ar_as_w1 \PWM3/State_reg  (
    .clk(clk100m),
    .d(\PWM3/n10 ),
    .en(1'b1),
    .reset(~rstn),
    .set(1'b0),
    .q(pwm_state_read[3]));  // src/OnePWM.v(26)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[0]  (
    .i(\PWM3/RemaTxNum[0]_keep ),
    .o(pnumcnt3[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[10]  (
    .i(\PWM3/RemaTxNum[10]_keep ),
    .o(pnumcnt3[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[11]  (
    .i(\PWM3/RemaTxNum[11]_keep ),
    .o(pnumcnt3[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[12]  (
    .i(\PWM3/RemaTxNum[12]_keep ),
    .o(pnumcnt3[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[13]  (
    .i(\PWM3/RemaTxNum[13]_keep ),
    .o(pnumcnt3[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[14]  (
    .i(\PWM3/RemaTxNum[14]_keep ),
    .o(pnumcnt3[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[15]  (
    .i(\PWM3/RemaTxNum[15]_keep ),
    .o(pnumcnt3[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[16]  (
    .i(\PWM3/RemaTxNum[16]_keep ),
    .o(pnumcnt3[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[17]  (
    .i(\PWM3/RemaTxNum[17]_keep ),
    .o(pnumcnt3[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[18]  (
    .i(\PWM3/RemaTxNum[18]_keep ),
    .o(pnumcnt3[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[19]  (
    .i(\PWM3/RemaTxNum[19]_keep ),
    .o(pnumcnt3[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[1]  (
    .i(\PWM3/RemaTxNum[1]_keep ),
    .o(pnumcnt3[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[20]  (
    .i(\PWM3/RemaTxNum[20]_keep ),
    .o(pnumcnt3[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[21]  (
    .i(\PWM3/RemaTxNum[21]_keep ),
    .o(pnumcnt3[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[22]  (
    .i(\PWM3/RemaTxNum[22]_keep ),
    .o(pnumcnt3[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[23]  (
    .i(\PWM3/RemaTxNum[23]_keep ),
    .o(pnumcnt3[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[2]  (
    .i(\PWM3/RemaTxNum[2]_keep ),
    .o(pnumcnt3[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[3]  (
    .i(\PWM3/RemaTxNum[3]_keep ),
    .o(pnumcnt3[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[4]  (
    .i(\PWM3/RemaTxNum[4]_keep ),
    .o(pnumcnt3[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[5]  (
    .i(\PWM3/RemaTxNum[5]_keep ),
    .o(pnumcnt3[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[6]  (
    .i(\PWM3/RemaTxNum[6]_keep ),
    .o(pnumcnt3[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[7]  (
    .i(\PWM3/RemaTxNum[7]_keep ),
    .o(pnumcnt3[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[8]  (
    .i(\PWM3/RemaTxNum[8]_keep ),
    .o(pnumcnt3[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[9]  (
    .i(\PWM3/RemaTxNum[9]_keep ),
    .o(pnumcnt3[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_dir  (
    .i(\PWM3/dir_keep ),
    .o(dir_pad[3]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[0]  (
    .i(\PWM3/pnumr[0]_keep ),
    .o(\PWM3/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[10]  (
    .i(\PWM3/pnumr[10]_keep ),
    .o(\PWM3/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[11]  (
    .i(\PWM3/pnumr[11]_keep ),
    .o(\PWM3/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[12]  (
    .i(\PWM3/pnumr[12]_keep ),
    .o(\PWM3/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[13]  (
    .i(\PWM3/pnumr[13]_keep ),
    .o(\PWM3/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[14]  (
    .i(\PWM3/pnumr[14]_keep ),
    .o(\PWM3/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[15]  (
    .i(\PWM3/pnumr[15]_keep ),
    .o(\PWM3/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[16]  (
    .i(\PWM3/pnumr[16]_keep ),
    .o(\PWM3/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[17]  (
    .i(\PWM3/pnumr[17]_keep ),
    .o(\PWM3/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[18]  (
    .i(\PWM3/pnumr[18]_keep ),
    .o(\PWM3/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[19]  (
    .i(\PWM3/pnumr[19]_keep ),
    .o(\PWM3/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[1]  (
    .i(\PWM3/pnumr[1]_keep ),
    .o(\PWM3/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[20]  (
    .i(\PWM3/pnumr[20]_keep ),
    .o(\PWM3/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[21]  (
    .i(\PWM3/pnumr[21]_keep ),
    .o(\PWM3/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[22]  (
    .i(\PWM3/pnumr[22]_keep ),
    .o(\PWM3/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[23]  (
    .i(\PWM3/pnumr[23]_keep ),
    .o(\PWM3/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[24]  (
    .i(\PWM3/pnumr[24]_keep ),
    .o(\PWM3/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[25]  (
    .i(\PWM3/pnumr[25]_keep ),
    .o(\PWM3/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[26]  (
    .i(\PWM3/pnumr[26]_keep ),
    .o(\PWM3/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[27]  (
    .i(\PWM3/pnumr[27]_keep ),
    .o(\PWM3/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[28]  (
    .i(\PWM3/pnumr[28]_keep ),
    .o(\PWM3/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[29]  (
    .i(\PWM3/pnumr[29]_keep ),
    .o(\PWM3/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[2]  (
    .i(\PWM3/pnumr[2]_keep ),
    .o(\PWM3/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[30]  (
    .i(\PWM3/pnumr[30]_keep ),
    .o(\PWM3/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[31]  (
    .i(\PWM3/pnumr[31]_keep ),
    .o(\PWM3/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[3]  (
    .i(\PWM3/pnumr[3]_keep ),
    .o(\PWM3/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[4]  (
    .i(\PWM3/pnumr[4]_keep ),
    .o(\PWM3/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[5]  (
    .i(\PWM3/pnumr[5]_keep ),
    .o(\PWM3/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[6]  (
    .i(\PWM3/pnumr[6]_keep ),
    .o(\PWM3/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[7]  (
    .i(\PWM3/pnumr[7]_keep ),
    .o(\PWM3/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[8]  (
    .i(\PWM3/pnumr[8]_keep ),
    .o(\PWM3/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[9]  (
    .i(\PWM3/pnumr[9]_keep ),
    .o(\PWM3/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pwm  (
    .i(\PWM3/pwm_keep ),
    .o(pwm_pad[3]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_stopreq  (
    .i(\PWM3/stopreq_keep ),
    .o(\PWM3/stopreq ));  // src/OnePWM.v(14)
  reg_ar_as_w1 \PWM3/dir_reg  (
    .clk(clk100m),
    .d(\PWM3/n32 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/dir_keep ));  // src/OnePWM.v(58)
  reg_sr_as_w1 \PWM3/pwm_reg  (
    .clk(clk100m),
    .d(\pwm[3]_d ),
    .en(1'b1),
    .reset(~\PWM3/u14_sel_is_1_o ),
    .set(1'b0),
    .q(\PWM3/pwm_keep ));  // src/OnePWM.v(45)
  reg_sr_as_w1 \PWM3/reg0_b0  (
    .clk(clk100m),
    .d(\PWM3/n13 [0]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [0]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b1  (
    .clk(clk100m),
    .d(\PWM3/n13 [1]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [1]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b10  (
    .clk(clk100m),
    .d(\PWM3/n13 [10]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [10]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b11  (
    .clk(clk100m),
    .d(\PWM3/n13 [11]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [11]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b12  (
    .clk(clk100m),
    .d(\PWM3/n13 [12]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [12]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b13  (
    .clk(clk100m),
    .d(\PWM3/n13 [13]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [13]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b14  (
    .clk(clk100m),
    .d(\PWM3/n13 [14]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [14]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b15  (
    .clk(clk100m),
    .d(\PWM3/n13 [15]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [15]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b16  (
    .clk(clk100m),
    .d(\PWM3/n13 [16]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [16]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b17  (
    .clk(clk100m),
    .d(\PWM3/n13 [17]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [17]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b18  (
    .clk(clk100m),
    .d(\PWM3/n13 [18]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [18]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b19  (
    .clk(clk100m),
    .d(\PWM3/n13 [19]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [19]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b2  (
    .clk(clk100m),
    .d(\PWM3/n13 [2]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [2]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b20  (
    .clk(clk100m),
    .d(\PWM3/n13 [20]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [20]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b21  (
    .clk(clk100m),
    .d(\PWM3/n13 [21]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [21]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b22  (
    .clk(clk100m),
    .d(\PWM3/n13 [22]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [22]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b23  (
    .clk(clk100m),
    .d(\PWM3/n13 [23]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [23]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b24  (
    .clk(clk100m),
    .d(\PWM3/n13 [24]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [24]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b25  (
    .clk(clk100m),
    .d(\PWM3/n13 [25]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [25]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b26  (
    .clk(clk100m),
    .d(\PWM3/n13 [26]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [26]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b3  (
    .clk(clk100m),
    .d(\PWM3/n13 [3]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [3]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b4  (
    .clk(clk100m),
    .d(\PWM3/n13 [4]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [4]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b5  (
    .clk(clk100m),
    .d(\PWM3/n13 [5]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [5]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b6  (
    .clk(clk100m),
    .d(\PWM3/n13 [6]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [6]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b7  (
    .clk(clk100m),
    .d(\PWM3/n13 [7]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [7]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b8  (
    .clk(clk100m),
    .d(\PWM3/n13 [8]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [8]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b9  (
    .clk(clk100m),
    .d(\PWM3/n13 [9]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b0  (
    .clk(clk100m),
    .d(freq3[0]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [0]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b1  (
    .clk(clk100m),
    .d(freq3[1]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [1]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b10  (
    .clk(clk100m),
    .d(freq3[10]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [10]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b11  (
    .clk(clk100m),
    .d(freq3[11]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [11]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b12  (
    .clk(clk100m),
    .d(freq3[12]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [12]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b13  (
    .clk(clk100m),
    .d(freq3[13]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [13]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b14  (
    .clk(clk100m),
    .d(freq3[14]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [14]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b15  (
    .clk(clk100m),
    .d(freq3[15]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [15]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b16  (
    .clk(clk100m),
    .d(freq3[16]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [16]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b17  (
    .clk(clk100m),
    .d(freq3[17]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [17]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b18  (
    .clk(clk100m),
    .d(freq3[18]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [18]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b19  (
    .clk(clk100m),
    .d(freq3[19]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [19]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b2  (
    .clk(clk100m),
    .d(freq3[2]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [2]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b20  (
    .clk(clk100m),
    .d(freq3[20]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [20]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b21  (
    .clk(clk100m),
    .d(freq3[21]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [21]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b22  (
    .clk(clk100m),
    .d(freq3[22]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [22]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b23  (
    .clk(clk100m),
    .d(freq3[23]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [23]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b24  (
    .clk(clk100m),
    .d(freq3[24]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [24]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b25  (
    .clk(clk100m),
    .d(freq3[25]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [25]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b26  (
    .clk(clk100m),
    .d(freq3[26]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [26]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b3  (
    .clk(clk100m),
    .d(freq3[3]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [3]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b4  (
    .clk(clk100m),
    .d(freq3[4]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [4]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b5  (
    .clk(clk100m),
    .d(freq3[5]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [5]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b6  (
    .clk(clk100m),
    .d(freq3[6]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [6]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b7  (
    .clk(clk100m),
    .d(freq3[7]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [7]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b8  (
    .clk(clk100m),
    .d(freq3[8]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [8]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b9  (
    .clk(clk100m),
    .d(freq3[9]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg2_b0  (
    .clk(clk100m),
    .d(\PWM3/n23 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[0]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b1  (
    .clk(clk100m),
    .d(\PWM3/n23 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[1]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b10  (
    .clk(clk100m),
    .d(\PWM3/n23 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[10]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b11  (
    .clk(clk100m),
    .d(\PWM3/n23 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[11]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b12  (
    .clk(clk100m),
    .d(\PWM3/n23 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[12]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b13  (
    .clk(clk100m),
    .d(\PWM3/n23 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[13]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b14  (
    .clk(clk100m),
    .d(\PWM3/n23 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[14]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b15  (
    .clk(clk100m),
    .d(\PWM3/n23 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[15]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b16  (
    .clk(clk100m),
    .d(\PWM3/n23 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[16]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b17  (
    .clk(clk100m),
    .d(\PWM3/n23 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[17]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b18  (
    .clk(clk100m),
    .d(\PWM3/n23 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[18]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b19  (
    .clk(clk100m),
    .d(\PWM3/n23 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[19]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b2  (
    .clk(clk100m),
    .d(\PWM3/n23 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[2]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b20  (
    .clk(clk100m),
    .d(\PWM3/n23 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[20]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b21  (
    .clk(clk100m),
    .d(\PWM3/n23 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[21]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b22  (
    .clk(clk100m),
    .d(\PWM3/n23 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[22]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b23  (
    .clk(clk100m),
    .d(\PWM3/n23 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[23]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b24  (
    .clk(clk100m),
    .d(\PWM3/n23 [24]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[24]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b25  (
    .clk(clk100m),
    .d(\PWM3/n23 [25]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[25]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b26  (
    .clk(clk100m),
    .d(\PWM3/n23 [26]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[26]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b27  (
    .clk(clk100m),
    .d(\PWM3/n23 [27]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[27]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b28  (
    .clk(clk100m),
    .d(\PWM3/n23 [28]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[28]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b29  (
    .clk(clk100m),
    .d(\PWM3/n23 [29]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[29]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b3  (
    .clk(clk100m),
    .d(\PWM3/n23 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[3]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b30  (
    .clk(clk100m),
    .d(\PWM3/n23 [30]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[30]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b31  (
    .clk(clk100m),
    .d(\PWM3/n23 [31]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[31]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b4  (
    .clk(clk100m),
    .d(\PWM3/n23 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[4]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b5  (
    .clk(clk100m),
    .d(\PWM3/n23 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[5]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b6  (
    .clk(clk100m),
    .d(\PWM3/n23 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[6]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b7  (
    .clk(clk100m),
    .d(\PWM3/n23 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[7]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b8  (
    .clk(clk100m),
    .d(\PWM3/n23 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[8]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b9  (
    .clk(clk100m),
    .d(\PWM3/n23 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[9]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg3_b0  (
    .clk(clk100m),
    .d(\PWM3/n31 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[0]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b1  (
    .clk(clk100m),
    .d(\PWM3/n31 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[1]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b10  (
    .clk(clk100m),
    .d(\PWM3/n31 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[10]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b11  (
    .clk(clk100m),
    .d(\PWM3/n31 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[11]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b12  (
    .clk(clk100m),
    .d(\PWM3/n31 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[12]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b13  (
    .clk(clk100m),
    .d(\PWM3/n31 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[13]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b14  (
    .clk(clk100m),
    .d(\PWM3/n31 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[14]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b15  (
    .clk(clk100m),
    .d(\PWM3/n31 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[15]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b16  (
    .clk(clk100m),
    .d(\PWM3/n31 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[16]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b17  (
    .clk(clk100m),
    .d(\PWM3/n31 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[17]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b18  (
    .clk(clk100m),
    .d(\PWM3/n31 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[18]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b19  (
    .clk(clk100m),
    .d(\PWM3/n31 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[19]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b2  (
    .clk(clk100m),
    .d(\PWM3/n31 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[2]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b20  (
    .clk(clk100m),
    .d(\PWM3/n31 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[20]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b21  (
    .clk(clk100m),
    .d(\PWM3/n31 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[21]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b22  (
    .clk(clk100m),
    .d(\PWM3/n31 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[22]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b23  (
    .clk(clk100m),
    .d(\PWM3/n31 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[23]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b3  (
    .clk(clk100m),
    .d(\PWM3/n31 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[3]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b4  (
    .clk(clk100m),
    .d(\PWM3/n31 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[4]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b5  (
    .clk(clk100m),
    .d(\PWM3/n31 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[5]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b6  (
    .clk(clk100m),
    .d(\PWM3/n31 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[6]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b7  (
    .clk(clk100m),
    .d(\PWM3/n31 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[7]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b8  (
    .clk(clk100m),
    .d(\PWM3/n31 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[8]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b9  (
    .clk(clk100m),
    .d(\PWM3/n31 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[9]_keep ));  // src/OnePWM.v(58)
  reg_ar_ss_w1 \PWM3/stopreq_reg  (
    .clk(clk100m),
    .d(\PWM3/n1 ),
    .en(1'b1),
    .reset(1'b0),
    .set(pwm_start_stop[3]),
    .q(\PWM3/stopreq_keep ));  // src/OnePWM.v(15)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub0/u0  (
    .a(\PWM3/FreCnt [0]),
    .b(1'b1),
    .c(\PWM3/sub0/c0 ),
    .o({\PWM3/sub0/c1 ,\PWM3/n12 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub0/u1  (
    .a(\PWM3/FreCnt [1]),
    .b(1'b0),
    .c(\PWM3/sub0/c1 ),
    .o({\PWM3/sub0/c2 ,\PWM3/n12 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub0/u10  (
    .a(\PWM3/FreCnt [10]),
    .b(1'b0),
    .c(\PWM3/sub0/c10 ),
    .o({\PWM3/sub0/c11 ,\PWM3/n12 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub0/u11  (
    .a(\PWM3/FreCnt [11]),
    .b(1'b0),
    .c(\PWM3/sub0/c11 ),
    .o({\PWM3/sub0/c12 ,\PWM3/n12 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub0/u12  (
    .a(\PWM3/FreCnt [12]),
    .b(1'b0),
    .c(\PWM3/sub0/c12 ),
    .o({\PWM3/sub0/c13 ,\PWM3/n12 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub0/u13  (
    .a(\PWM3/FreCnt [13]),
    .b(1'b0),
    .c(\PWM3/sub0/c13 ),
    .o({\PWM3/sub0/c14 ,\PWM3/n12 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub0/u14  (
    .a(\PWM3/FreCnt [14]),
    .b(1'b0),
    .c(\PWM3/sub0/c14 ),
    .o({\PWM3/sub0/c15 ,\PWM3/n12 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub0/u15  (
    .a(\PWM3/FreCnt [15]),
    .b(1'b0),
    .c(\PWM3/sub0/c15 ),
    .o({\PWM3/sub0/c16 ,\PWM3/n12 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub0/u16  (
    .a(\PWM3/FreCnt [16]),
    .b(1'b0),
    .c(\PWM3/sub0/c16 ),
    .o({\PWM3/sub0/c17 ,\PWM3/n12 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub0/u17  (
    .a(\PWM3/FreCnt [17]),
    .b(1'b0),
    .c(\PWM3/sub0/c17 ),
    .o({\PWM3/sub0/c18 ,\PWM3/n12 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub0/u18  (
    .a(\PWM3/FreCnt [18]),
    .b(1'b0),
    .c(\PWM3/sub0/c18 ),
    .o({\PWM3/sub0/c19 ,\PWM3/n12 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub0/u19  (
    .a(\PWM3/FreCnt [19]),
    .b(1'b0),
    .c(\PWM3/sub0/c19 ),
    .o({\PWM3/sub0/c20 ,\PWM3/n12 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub0/u2  (
    .a(\PWM3/FreCnt [2]),
    .b(1'b0),
    .c(\PWM3/sub0/c2 ),
    .o({\PWM3/sub0/c3 ,\PWM3/n12 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub0/u20  (
    .a(\PWM3/FreCnt [20]),
    .b(1'b0),
    .c(\PWM3/sub0/c20 ),
    .o({\PWM3/sub0/c21 ,\PWM3/n12 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub0/u21  (
    .a(\PWM3/FreCnt [21]),
    .b(1'b0),
    .c(\PWM3/sub0/c21 ),
    .o({\PWM3/sub0/c22 ,\PWM3/n12 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub0/u22  (
    .a(\PWM3/FreCnt [22]),
    .b(1'b0),
    .c(\PWM3/sub0/c22 ),
    .o({\PWM3/sub0/c23 ,\PWM3/n12 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub0/u23  (
    .a(\PWM3/FreCnt [23]),
    .b(1'b0),
    .c(\PWM3/sub0/c23 ),
    .o({\PWM3/sub0/c24 ,\PWM3/n12 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub0/u24  (
    .a(\PWM3/FreCnt [24]),
    .b(1'b0),
    .c(\PWM3/sub0/c24 ),
    .o({\PWM3/sub0/c25 ,\PWM3/n12 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub0/u25  (
    .a(\PWM3/FreCnt [25]),
    .b(1'b0),
    .c(\PWM3/sub0/c25 ),
    .o({\PWM3/sub0/c26 ,\PWM3/n12 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub0/u26  (
    .a(\PWM3/FreCnt [26]),
    .b(1'b0),
    .c(\PWM3/sub0/c26 ),
    .o({open_n24,\PWM3/n12 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub0/u3  (
    .a(\PWM3/FreCnt [3]),
    .b(1'b0),
    .c(\PWM3/sub0/c3 ),
    .o({\PWM3/sub0/c4 ,\PWM3/n12 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub0/u4  (
    .a(\PWM3/FreCnt [4]),
    .b(1'b0),
    .c(\PWM3/sub0/c4 ),
    .o({\PWM3/sub0/c5 ,\PWM3/n12 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub0/u5  (
    .a(\PWM3/FreCnt [5]),
    .b(1'b0),
    .c(\PWM3/sub0/c5 ),
    .o({\PWM3/sub0/c6 ,\PWM3/n12 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub0/u6  (
    .a(\PWM3/FreCnt [6]),
    .b(1'b0),
    .c(\PWM3/sub0/c6 ),
    .o({\PWM3/sub0/c7 ,\PWM3/n12 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub0/u7  (
    .a(\PWM3/FreCnt [7]),
    .b(1'b0),
    .c(\PWM3/sub0/c7 ),
    .o({\PWM3/sub0/c8 ,\PWM3/n12 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub0/u8  (
    .a(\PWM3/FreCnt [8]),
    .b(1'b0),
    .c(\PWM3/sub0/c8 ),
    .o({\PWM3/sub0/c9 ,\PWM3/n12 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub0/u9  (
    .a(\PWM3/FreCnt [9]),
    .b(1'b0),
    .c(\PWM3/sub0/c9 ),
    .o({\PWM3/sub0/c10 ,\PWM3/n12 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \PWM3/sub0/ucin  (
    .a(1'b0),
    .o({\PWM3/sub0/c0 ,open_n27}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub1/u0  (
    .a(pnumcnt3[0]),
    .b(1'b1),
    .c(\PWM3/sub1/c0 ),
    .o({\PWM3/sub1/c1 ,\PWM3/n26 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub1/u1  (
    .a(pnumcnt3[1]),
    .b(1'b0),
    .c(\PWM3/sub1/c1 ),
    .o({\PWM3/sub1/c2 ,\PWM3/n26 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub1/u10  (
    .a(pnumcnt3[10]),
    .b(1'b0),
    .c(\PWM3/sub1/c10 ),
    .o({\PWM3/sub1/c11 ,\PWM3/n26 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub1/u11  (
    .a(pnumcnt3[11]),
    .b(1'b0),
    .c(\PWM3/sub1/c11 ),
    .o({\PWM3/sub1/c12 ,\PWM3/n26 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub1/u12  (
    .a(pnumcnt3[12]),
    .b(1'b0),
    .c(\PWM3/sub1/c12 ),
    .o({\PWM3/sub1/c13 ,\PWM3/n26 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub1/u13  (
    .a(pnumcnt3[13]),
    .b(1'b0),
    .c(\PWM3/sub1/c13 ),
    .o({\PWM3/sub1/c14 ,\PWM3/n26 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub1/u14  (
    .a(pnumcnt3[14]),
    .b(1'b0),
    .c(\PWM3/sub1/c14 ),
    .o({\PWM3/sub1/c15 ,\PWM3/n26 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub1/u15  (
    .a(pnumcnt3[15]),
    .b(1'b0),
    .c(\PWM3/sub1/c15 ),
    .o({\PWM3/sub1/c16 ,\PWM3/n26 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub1/u16  (
    .a(pnumcnt3[16]),
    .b(1'b0),
    .c(\PWM3/sub1/c16 ),
    .o({\PWM3/sub1/c17 ,\PWM3/n26 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub1/u17  (
    .a(pnumcnt3[17]),
    .b(1'b0),
    .c(\PWM3/sub1/c17 ),
    .o({\PWM3/sub1/c18 ,\PWM3/n26 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub1/u18  (
    .a(pnumcnt3[18]),
    .b(1'b0),
    .c(\PWM3/sub1/c18 ),
    .o({\PWM3/sub1/c19 ,\PWM3/n26 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub1/u19  (
    .a(pnumcnt3[19]),
    .b(1'b0),
    .c(\PWM3/sub1/c19 ),
    .o({\PWM3/sub1/c20 ,\PWM3/n26 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub1/u2  (
    .a(pnumcnt3[2]),
    .b(1'b0),
    .c(\PWM3/sub1/c2 ),
    .o({\PWM3/sub1/c3 ,\PWM3/n26 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub1/u20  (
    .a(pnumcnt3[20]),
    .b(1'b0),
    .c(\PWM3/sub1/c20 ),
    .o({\PWM3/sub1/c21 ,\PWM3/n26 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub1/u21  (
    .a(pnumcnt3[21]),
    .b(1'b0),
    .c(\PWM3/sub1/c21 ),
    .o({\PWM3/sub1/c22 ,\PWM3/n26 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub1/u22  (
    .a(pnumcnt3[22]),
    .b(1'b0),
    .c(\PWM3/sub1/c22 ),
    .o({\PWM3/sub1/c23 ,\PWM3/n26 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub1/u23  (
    .a(pnumcnt3[23]),
    .b(1'b0),
    .c(\PWM3/sub1/c23 ),
    .o({open_n28,\PWM3/n26 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub1/u3  (
    .a(pnumcnt3[3]),
    .b(1'b0),
    .c(\PWM3/sub1/c3 ),
    .o({\PWM3/sub1/c4 ,\PWM3/n26 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub1/u4  (
    .a(pnumcnt3[4]),
    .b(1'b0),
    .c(\PWM3/sub1/c4 ),
    .o({\PWM3/sub1/c5 ,\PWM3/n26 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub1/u5  (
    .a(pnumcnt3[5]),
    .b(1'b0),
    .c(\PWM3/sub1/c5 ),
    .o({\PWM3/sub1/c6 ,\PWM3/n26 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub1/u6  (
    .a(pnumcnt3[6]),
    .b(1'b0),
    .c(\PWM3/sub1/c6 ),
    .o({\PWM3/sub1/c7 ,\PWM3/n26 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub1/u7  (
    .a(pnumcnt3[7]),
    .b(1'b0),
    .c(\PWM3/sub1/c7 ),
    .o({\PWM3/sub1/c8 ,\PWM3/n26 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub1/u8  (
    .a(pnumcnt3[8]),
    .b(1'b0),
    .c(\PWM3/sub1/c8 ),
    .o({\PWM3/sub1/c9 ,\PWM3/n26 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM3/sub1/u9  (
    .a(pnumcnt3[9]),
    .b(1'b0),
    .c(\PWM3/sub1/c9 ),
    .o({\PWM3/sub1/c10 ,\PWM3/n26 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \PWM3/sub1/ucin  (
    .a(1'b0),
    .o({\PWM3/sub1/c0 ,open_n31}));
  reg_ar_as_w1 \PWM4/State_reg  (
    .clk(clk100m),
    .d(\PWM4/n10 ),
    .en(1'b1),
    .reset(~rstn),
    .set(1'b0),
    .q(pwm_state_read[4]));  // src/OnePWM.v(26)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[0]  (
    .i(\PWM4/RemaTxNum[0]_keep ),
    .o(pnumcnt4[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[10]  (
    .i(\PWM4/RemaTxNum[10]_keep ),
    .o(pnumcnt4[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[11]  (
    .i(\PWM4/RemaTxNum[11]_keep ),
    .o(pnumcnt4[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[12]  (
    .i(\PWM4/RemaTxNum[12]_keep ),
    .o(pnumcnt4[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[13]  (
    .i(\PWM4/RemaTxNum[13]_keep ),
    .o(pnumcnt4[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[14]  (
    .i(\PWM4/RemaTxNum[14]_keep ),
    .o(pnumcnt4[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[15]  (
    .i(\PWM4/RemaTxNum[15]_keep ),
    .o(pnumcnt4[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[16]  (
    .i(\PWM4/RemaTxNum[16]_keep ),
    .o(pnumcnt4[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[17]  (
    .i(\PWM4/RemaTxNum[17]_keep ),
    .o(pnumcnt4[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[18]  (
    .i(\PWM4/RemaTxNum[18]_keep ),
    .o(pnumcnt4[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[19]  (
    .i(\PWM4/RemaTxNum[19]_keep ),
    .o(pnumcnt4[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[1]  (
    .i(\PWM4/RemaTxNum[1]_keep ),
    .o(pnumcnt4[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[20]  (
    .i(\PWM4/RemaTxNum[20]_keep ),
    .o(pnumcnt4[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[21]  (
    .i(\PWM4/RemaTxNum[21]_keep ),
    .o(pnumcnt4[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[22]  (
    .i(\PWM4/RemaTxNum[22]_keep ),
    .o(pnumcnt4[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[23]  (
    .i(\PWM4/RemaTxNum[23]_keep ),
    .o(pnumcnt4[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[2]  (
    .i(\PWM4/RemaTxNum[2]_keep ),
    .o(pnumcnt4[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[3]  (
    .i(\PWM4/RemaTxNum[3]_keep ),
    .o(pnumcnt4[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[4]  (
    .i(\PWM4/RemaTxNum[4]_keep ),
    .o(pnumcnt4[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[5]  (
    .i(\PWM4/RemaTxNum[5]_keep ),
    .o(pnumcnt4[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[6]  (
    .i(\PWM4/RemaTxNum[6]_keep ),
    .o(pnumcnt4[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[7]  (
    .i(\PWM4/RemaTxNum[7]_keep ),
    .o(pnumcnt4[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[8]  (
    .i(\PWM4/RemaTxNum[8]_keep ),
    .o(pnumcnt4[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[9]  (
    .i(\PWM4/RemaTxNum[9]_keep ),
    .o(pnumcnt4[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_dir  (
    .i(\PWM4/dir_keep ),
    .o(dir_pad[4]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[0]  (
    .i(\PWM4/pnumr[0]_keep ),
    .o(\PWM4/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[10]  (
    .i(\PWM4/pnumr[10]_keep ),
    .o(\PWM4/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[11]  (
    .i(\PWM4/pnumr[11]_keep ),
    .o(\PWM4/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[12]  (
    .i(\PWM4/pnumr[12]_keep ),
    .o(\PWM4/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[13]  (
    .i(\PWM4/pnumr[13]_keep ),
    .o(\PWM4/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[14]  (
    .i(\PWM4/pnumr[14]_keep ),
    .o(\PWM4/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[15]  (
    .i(\PWM4/pnumr[15]_keep ),
    .o(\PWM4/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[16]  (
    .i(\PWM4/pnumr[16]_keep ),
    .o(\PWM4/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[17]  (
    .i(\PWM4/pnumr[17]_keep ),
    .o(\PWM4/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[18]  (
    .i(\PWM4/pnumr[18]_keep ),
    .o(\PWM4/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[19]  (
    .i(\PWM4/pnumr[19]_keep ),
    .o(\PWM4/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[1]  (
    .i(\PWM4/pnumr[1]_keep ),
    .o(\PWM4/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[20]  (
    .i(\PWM4/pnumr[20]_keep ),
    .o(\PWM4/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[21]  (
    .i(\PWM4/pnumr[21]_keep ),
    .o(\PWM4/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[22]  (
    .i(\PWM4/pnumr[22]_keep ),
    .o(\PWM4/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[23]  (
    .i(\PWM4/pnumr[23]_keep ),
    .o(\PWM4/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[24]  (
    .i(\PWM4/pnumr[24]_keep ),
    .o(\PWM4/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[25]  (
    .i(\PWM4/pnumr[25]_keep ),
    .o(\PWM4/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[26]  (
    .i(\PWM4/pnumr[26]_keep ),
    .o(\PWM4/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[27]  (
    .i(\PWM4/pnumr[27]_keep ),
    .o(\PWM4/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[28]  (
    .i(\PWM4/pnumr[28]_keep ),
    .o(\PWM4/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[29]  (
    .i(\PWM4/pnumr[29]_keep ),
    .o(\PWM4/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[2]  (
    .i(\PWM4/pnumr[2]_keep ),
    .o(\PWM4/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[30]  (
    .i(\PWM4/pnumr[30]_keep ),
    .o(\PWM4/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[31]  (
    .i(\PWM4/pnumr[31]_keep ),
    .o(\PWM4/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[3]  (
    .i(\PWM4/pnumr[3]_keep ),
    .o(\PWM4/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[4]  (
    .i(\PWM4/pnumr[4]_keep ),
    .o(\PWM4/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[5]  (
    .i(\PWM4/pnumr[5]_keep ),
    .o(\PWM4/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[6]  (
    .i(\PWM4/pnumr[6]_keep ),
    .o(\PWM4/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[7]  (
    .i(\PWM4/pnumr[7]_keep ),
    .o(\PWM4/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[8]  (
    .i(\PWM4/pnumr[8]_keep ),
    .o(\PWM4/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[9]  (
    .i(\PWM4/pnumr[9]_keep ),
    .o(\PWM4/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pwm  (
    .i(\PWM4/pwm_keep ),
    .o(pwm_pad[4]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_stopreq  (
    .i(\PWM4/stopreq_keep ),
    .o(\PWM4/stopreq ));  // src/OnePWM.v(14)
  reg_ar_as_w1 \PWM4/dir_reg  (
    .clk(clk100m),
    .d(\PWM4/n32 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/dir_keep ));  // src/OnePWM.v(58)
  reg_sr_as_w1 \PWM4/pwm_reg  (
    .clk(clk100m),
    .d(\pwm[4]_d ),
    .en(1'b1),
    .reset(~\PWM4/u14_sel_is_1_o ),
    .set(1'b0),
    .q(\PWM4/pwm_keep ));  // src/OnePWM.v(45)
  reg_sr_as_w1 \PWM4/reg0_b0  (
    .clk(clk100m),
    .d(\PWM4/n13 [0]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [0]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b1  (
    .clk(clk100m),
    .d(\PWM4/n13 [1]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [1]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b10  (
    .clk(clk100m),
    .d(\PWM4/n13 [10]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [10]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b11  (
    .clk(clk100m),
    .d(\PWM4/n13 [11]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [11]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b12  (
    .clk(clk100m),
    .d(\PWM4/n13 [12]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [12]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b13  (
    .clk(clk100m),
    .d(\PWM4/n13 [13]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [13]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b14  (
    .clk(clk100m),
    .d(\PWM4/n13 [14]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [14]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b15  (
    .clk(clk100m),
    .d(\PWM4/n13 [15]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [15]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b16  (
    .clk(clk100m),
    .d(\PWM4/n13 [16]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [16]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b17  (
    .clk(clk100m),
    .d(\PWM4/n13 [17]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [17]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b18  (
    .clk(clk100m),
    .d(\PWM4/n13 [18]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [18]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b19  (
    .clk(clk100m),
    .d(\PWM4/n13 [19]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [19]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b2  (
    .clk(clk100m),
    .d(\PWM4/n13 [2]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [2]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b20  (
    .clk(clk100m),
    .d(\PWM4/n13 [20]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [20]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b21  (
    .clk(clk100m),
    .d(\PWM4/n13 [21]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [21]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b22  (
    .clk(clk100m),
    .d(\PWM4/n13 [22]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [22]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b23  (
    .clk(clk100m),
    .d(\PWM4/n13 [23]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [23]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b24  (
    .clk(clk100m),
    .d(\PWM4/n13 [24]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [24]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b25  (
    .clk(clk100m),
    .d(\PWM4/n13 [25]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [25]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b26  (
    .clk(clk100m),
    .d(\PWM4/n13 [26]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [26]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b3  (
    .clk(clk100m),
    .d(\PWM4/n13 [3]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [3]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b4  (
    .clk(clk100m),
    .d(\PWM4/n13 [4]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [4]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b5  (
    .clk(clk100m),
    .d(\PWM4/n13 [5]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [5]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b6  (
    .clk(clk100m),
    .d(\PWM4/n13 [6]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [6]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b7  (
    .clk(clk100m),
    .d(\PWM4/n13 [7]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [7]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b8  (
    .clk(clk100m),
    .d(\PWM4/n13 [8]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [8]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b9  (
    .clk(clk100m),
    .d(\PWM4/n13 [9]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b0  (
    .clk(clk100m),
    .d(freq4[0]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [0]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b1  (
    .clk(clk100m),
    .d(freq4[1]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [1]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b10  (
    .clk(clk100m),
    .d(freq4[10]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [10]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b11  (
    .clk(clk100m),
    .d(freq4[11]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [11]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b12  (
    .clk(clk100m),
    .d(freq4[12]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [12]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b13  (
    .clk(clk100m),
    .d(freq4[13]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [13]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b14  (
    .clk(clk100m),
    .d(freq4[14]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [14]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b15  (
    .clk(clk100m),
    .d(freq4[15]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [15]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b16  (
    .clk(clk100m),
    .d(freq4[16]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [16]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b17  (
    .clk(clk100m),
    .d(freq4[17]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [17]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b18  (
    .clk(clk100m),
    .d(freq4[18]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [18]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b19  (
    .clk(clk100m),
    .d(freq4[19]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [19]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b2  (
    .clk(clk100m),
    .d(freq4[2]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [2]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b20  (
    .clk(clk100m),
    .d(freq4[20]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [20]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b21  (
    .clk(clk100m),
    .d(freq4[21]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [21]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b22  (
    .clk(clk100m),
    .d(freq4[22]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [22]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b23  (
    .clk(clk100m),
    .d(freq4[23]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [23]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b24  (
    .clk(clk100m),
    .d(freq4[24]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [24]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b25  (
    .clk(clk100m),
    .d(freq4[25]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [25]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b26  (
    .clk(clk100m),
    .d(freq4[26]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [26]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b3  (
    .clk(clk100m),
    .d(freq4[3]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [3]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b4  (
    .clk(clk100m),
    .d(freq4[4]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [4]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b5  (
    .clk(clk100m),
    .d(freq4[5]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [5]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b6  (
    .clk(clk100m),
    .d(freq4[6]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [6]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b7  (
    .clk(clk100m),
    .d(freq4[7]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [7]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b8  (
    .clk(clk100m),
    .d(freq4[8]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [8]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b9  (
    .clk(clk100m),
    .d(freq4[9]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg2_b0  (
    .clk(clk100m),
    .d(\PWM4/n23 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[0]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b1  (
    .clk(clk100m),
    .d(\PWM4/n23 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[1]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b10  (
    .clk(clk100m),
    .d(\PWM4/n23 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[10]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b11  (
    .clk(clk100m),
    .d(\PWM4/n23 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[11]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b12  (
    .clk(clk100m),
    .d(\PWM4/n23 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[12]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b13  (
    .clk(clk100m),
    .d(\PWM4/n23 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[13]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b14  (
    .clk(clk100m),
    .d(\PWM4/n23 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[14]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b15  (
    .clk(clk100m),
    .d(\PWM4/n23 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[15]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b16  (
    .clk(clk100m),
    .d(\PWM4/n23 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[16]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b17  (
    .clk(clk100m),
    .d(\PWM4/n23 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[17]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b18  (
    .clk(clk100m),
    .d(\PWM4/n23 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[18]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b19  (
    .clk(clk100m),
    .d(\PWM4/n23 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[19]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b2  (
    .clk(clk100m),
    .d(\PWM4/n23 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[2]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b20  (
    .clk(clk100m),
    .d(\PWM4/n23 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[20]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b21  (
    .clk(clk100m),
    .d(\PWM4/n23 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[21]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b22  (
    .clk(clk100m),
    .d(\PWM4/n23 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[22]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b23  (
    .clk(clk100m),
    .d(\PWM4/n23 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[23]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b24  (
    .clk(clk100m),
    .d(\PWM4/n23 [24]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[24]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b25  (
    .clk(clk100m),
    .d(\PWM4/n23 [25]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[25]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b26  (
    .clk(clk100m),
    .d(\PWM4/n23 [26]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[26]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b27  (
    .clk(clk100m),
    .d(\PWM4/n23 [27]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[27]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b28  (
    .clk(clk100m),
    .d(\PWM4/n23 [28]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[28]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b29  (
    .clk(clk100m),
    .d(\PWM4/n23 [29]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[29]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b3  (
    .clk(clk100m),
    .d(\PWM4/n23 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[3]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b30  (
    .clk(clk100m),
    .d(\PWM4/n23 [30]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[30]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b31  (
    .clk(clk100m),
    .d(\PWM4/n23 [31]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[31]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b4  (
    .clk(clk100m),
    .d(\PWM4/n23 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[4]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b5  (
    .clk(clk100m),
    .d(\PWM4/n23 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[5]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b6  (
    .clk(clk100m),
    .d(\PWM4/n23 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[6]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b7  (
    .clk(clk100m),
    .d(\PWM4/n23 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[7]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b8  (
    .clk(clk100m),
    .d(\PWM4/n23 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[8]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b9  (
    .clk(clk100m),
    .d(\PWM4/n23 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[9]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg3_b0  (
    .clk(clk100m),
    .d(\PWM4/n31 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[0]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b1  (
    .clk(clk100m),
    .d(\PWM4/n31 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[1]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b10  (
    .clk(clk100m),
    .d(\PWM4/n31 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[10]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b11  (
    .clk(clk100m),
    .d(\PWM4/n31 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[11]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b12  (
    .clk(clk100m),
    .d(\PWM4/n31 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[12]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b13  (
    .clk(clk100m),
    .d(\PWM4/n31 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[13]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b14  (
    .clk(clk100m),
    .d(\PWM4/n31 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[14]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b15  (
    .clk(clk100m),
    .d(\PWM4/n31 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[15]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b16  (
    .clk(clk100m),
    .d(\PWM4/n31 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[16]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b17  (
    .clk(clk100m),
    .d(\PWM4/n31 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[17]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b18  (
    .clk(clk100m),
    .d(\PWM4/n31 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[18]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b19  (
    .clk(clk100m),
    .d(\PWM4/n31 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[19]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b2  (
    .clk(clk100m),
    .d(\PWM4/n31 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[2]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b20  (
    .clk(clk100m),
    .d(\PWM4/n31 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[20]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b21  (
    .clk(clk100m),
    .d(\PWM4/n31 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[21]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b22  (
    .clk(clk100m),
    .d(\PWM4/n31 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[22]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b23  (
    .clk(clk100m),
    .d(\PWM4/n31 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[23]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b3  (
    .clk(clk100m),
    .d(\PWM4/n31 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[3]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b4  (
    .clk(clk100m),
    .d(\PWM4/n31 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[4]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b5  (
    .clk(clk100m),
    .d(\PWM4/n31 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[5]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b6  (
    .clk(clk100m),
    .d(\PWM4/n31 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[6]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b7  (
    .clk(clk100m),
    .d(\PWM4/n31 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[7]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b8  (
    .clk(clk100m),
    .d(\PWM4/n31 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[8]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b9  (
    .clk(clk100m),
    .d(\PWM4/n31 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[9]_keep ));  // src/OnePWM.v(58)
  reg_ar_ss_w1 \PWM4/stopreq_reg  (
    .clk(clk100m),
    .d(\PWM4/n1 ),
    .en(1'b1),
    .reset(1'b0),
    .set(pwm_start_stop[4]),
    .q(\PWM4/stopreq_keep ));  // src/OnePWM.v(15)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub0/u0  (
    .a(\PWM4/FreCnt [0]),
    .b(1'b1),
    .c(\PWM4/sub0/c0 ),
    .o({\PWM4/sub0/c1 ,\PWM4/n12 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub0/u1  (
    .a(\PWM4/FreCnt [1]),
    .b(1'b0),
    .c(\PWM4/sub0/c1 ),
    .o({\PWM4/sub0/c2 ,\PWM4/n12 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub0/u10  (
    .a(\PWM4/FreCnt [10]),
    .b(1'b0),
    .c(\PWM4/sub0/c10 ),
    .o({\PWM4/sub0/c11 ,\PWM4/n12 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub0/u11  (
    .a(\PWM4/FreCnt [11]),
    .b(1'b0),
    .c(\PWM4/sub0/c11 ),
    .o({\PWM4/sub0/c12 ,\PWM4/n12 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub0/u12  (
    .a(\PWM4/FreCnt [12]),
    .b(1'b0),
    .c(\PWM4/sub0/c12 ),
    .o({\PWM4/sub0/c13 ,\PWM4/n12 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub0/u13  (
    .a(\PWM4/FreCnt [13]),
    .b(1'b0),
    .c(\PWM4/sub0/c13 ),
    .o({\PWM4/sub0/c14 ,\PWM4/n12 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub0/u14  (
    .a(\PWM4/FreCnt [14]),
    .b(1'b0),
    .c(\PWM4/sub0/c14 ),
    .o({\PWM4/sub0/c15 ,\PWM4/n12 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub0/u15  (
    .a(\PWM4/FreCnt [15]),
    .b(1'b0),
    .c(\PWM4/sub0/c15 ),
    .o({\PWM4/sub0/c16 ,\PWM4/n12 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub0/u16  (
    .a(\PWM4/FreCnt [16]),
    .b(1'b0),
    .c(\PWM4/sub0/c16 ),
    .o({\PWM4/sub0/c17 ,\PWM4/n12 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub0/u17  (
    .a(\PWM4/FreCnt [17]),
    .b(1'b0),
    .c(\PWM4/sub0/c17 ),
    .o({\PWM4/sub0/c18 ,\PWM4/n12 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub0/u18  (
    .a(\PWM4/FreCnt [18]),
    .b(1'b0),
    .c(\PWM4/sub0/c18 ),
    .o({\PWM4/sub0/c19 ,\PWM4/n12 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub0/u19  (
    .a(\PWM4/FreCnt [19]),
    .b(1'b0),
    .c(\PWM4/sub0/c19 ),
    .o({\PWM4/sub0/c20 ,\PWM4/n12 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub0/u2  (
    .a(\PWM4/FreCnt [2]),
    .b(1'b0),
    .c(\PWM4/sub0/c2 ),
    .o({\PWM4/sub0/c3 ,\PWM4/n12 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub0/u20  (
    .a(\PWM4/FreCnt [20]),
    .b(1'b0),
    .c(\PWM4/sub0/c20 ),
    .o({\PWM4/sub0/c21 ,\PWM4/n12 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub0/u21  (
    .a(\PWM4/FreCnt [21]),
    .b(1'b0),
    .c(\PWM4/sub0/c21 ),
    .o({\PWM4/sub0/c22 ,\PWM4/n12 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub0/u22  (
    .a(\PWM4/FreCnt [22]),
    .b(1'b0),
    .c(\PWM4/sub0/c22 ),
    .o({\PWM4/sub0/c23 ,\PWM4/n12 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub0/u23  (
    .a(\PWM4/FreCnt [23]),
    .b(1'b0),
    .c(\PWM4/sub0/c23 ),
    .o({\PWM4/sub0/c24 ,\PWM4/n12 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub0/u24  (
    .a(\PWM4/FreCnt [24]),
    .b(1'b0),
    .c(\PWM4/sub0/c24 ),
    .o({\PWM4/sub0/c25 ,\PWM4/n12 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub0/u25  (
    .a(\PWM4/FreCnt [25]),
    .b(1'b0),
    .c(\PWM4/sub0/c25 ),
    .o({\PWM4/sub0/c26 ,\PWM4/n12 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub0/u26  (
    .a(\PWM4/FreCnt [26]),
    .b(1'b0),
    .c(\PWM4/sub0/c26 ),
    .o({open_n32,\PWM4/n12 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub0/u3  (
    .a(\PWM4/FreCnt [3]),
    .b(1'b0),
    .c(\PWM4/sub0/c3 ),
    .o({\PWM4/sub0/c4 ,\PWM4/n12 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub0/u4  (
    .a(\PWM4/FreCnt [4]),
    .b(1'b0),
    .c(\PWM4/sub0/c4 ),
    .o({\PWM4/sub0/c5 ,\PWM4/n12 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub0/u5  (
    .a(\PWM4/FreCnt [5]),
    .b(1'b0),
    .c(\PWM4/sub0/c5 ),
    .o({\PWM4/sub0/c6 ,\PWM4/n12 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub0/u6  (
    .a(\PWM4/FreCnt [6]),
    .b(1'b0),
    .c(\PWM4/sub0/c6 ),
    .o({\PWM4/sub0/c7 ,\PWM4/n12 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub0/u7  (
    .a(\PWM4/FreCnt [7]),
    .b(1'b0),
    .c(\PWM4/sub0/c7 ),
    .o({\PWM4/sub0/c8 ,\PWM4/n12 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub0/u8  (
    .a(\PWM4/FreCnt [8]),
    .b(1'b0),
    .c(\PWM4/sub0/c8 ),
    .o({\PWM4/sub0/c9 ,\PWM4/n12 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub0/u9  (
    .a(\PWM4/FreCnt [9]),
    .b(1'b0),
    .c(\PWM4/sub0/c9 ),
    .o({\PWM4/sub0/c10 ,\PWM4/n12 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \PWM4/sub0/ucin  (
    .a(1'b0),
    .o({\PWM4/sub0/c0 ,open_n35}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub1/u0  (
    .a(pnumcnt4[0]),
    .b(1'b1),
    .c(\PWM4/sub1/c0 ),
    .o({\PWM4/sub1/c1 ,\PWM4/n26 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub1/u1  (
    .a(pnumcnt4[1]),
    .b(1'b0),
    .c(\PWM4/sub1/c1 ),
    .o({\PWM4/sub1/c2 ,\PWM4/n26 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub1/u10  (
    .a(pnumcnt4[10]),
    .b(1'b0),
    .c(\PWM4/sub1/c10 ),
    .o({\PWM4/sub1/c11 ,\PWM4/n26 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub1/u11  (
    .a(pnumcnt4[11]),
    .b(1'b0),
    .c(\PWM4/sub1/c11 ),
    .o({\PWM4/sub1/c12 ,\PWM4/n26 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub1/u12  (
    .a(pnumcnt4[12]),
    .b(1'b0),
    .c(\PWM4/sub1/c12 ),
    .o({\PWM4/sub1/c13 ,\PWM4/n26 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub1/u13  (
    .a(pnumcnt4[13]),
    .b(1'b0),
    .c(\PWM4/sub1/c13 ),
    .o({\PWM4/sub1/c14 ,\PWM4/n26 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub1/u14  (
    .a(pnumcnt4[14]),
    .b(1'b0),
    .c(\PWM4/sub1/c14 ),
    .o({\PWM4/sub1/c15 ,\PWM4/n26 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub1/u15  (
    .a(pnumcnt4[15]),
    .b(1'b0),
    .c(\PWM4/sub1/c15 ),
    .o({\PWM4/sub1/c16 ,\PWM4/n26 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub1/u16  (
    .a(pnumcnt4[16]),
    .b(1'b0),
    .c(\PWM4/sub1/c16 ),
    .o({\PWM4/sub1/c17 ,\PWM4/n26 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub1/u17  (
    .a(pnumcnt4[17]),
    .b(1'b0),
    .c(\PWM4/sub1/c17 ),
    .o({\PWM4/sub1/c18 ,\PWM4/n26 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub1/u18  (
    .a(pnumcnt4[18]),
    .b(1'b0),
    .c(\PWM4/sub1/c18 ),
    .o({\PWM4/sub1/c19 ,\PWM4/n26 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub1/u19  (
    .a(pnumcnt4[19]),
    .b(1'b0),
    .c(\PWM4/sub1/c19 ),
    .o({\PWM4/sub1/c20 ,\PWM4/n26 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub1/u2  (
    .a(pnumcnt4[2]),
    .b(1'b0),
    .c(\PWM4/sub1/c2 ),
    .o({\PWM4/sub1/c3 ,\PWM4/n26 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub1/u20  (
    .a(pnumcnt4[20]),
    .b(1'b0),
    .c(\PWM4/sub1/c20 ),
    .o({\PWM4/sub1/c21 ,\PWM4/n26 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub1/u21  (
    .a(pnumcnt4[21]),
    .b(1'b0),
    .c(\PWM4/sub1/c21 ),
    .o({\PWM4/sub1/c22 ,\PWM4/n26 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub1/u22  (
    .a(pnumcnt4[22]),
    .b(1'b0),
    .c(\PWM4/sub1/c22 ),
    .o({\PWM4/sub1/c23 ,\PWM4/n26 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub1/u23  (
    .a(pnumcnt4[23]),
    .b(1'b0),
    .c(\PWM4/sub1/c23 ),
    .o({open_n36,\PWM4/n26 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub1/u3  (
    .a(pnumcnt4[3]),
    .b(1'b0),
    .c(\PWM4/sub1/c3 ),
    .o({\PWM4/sub1/c4 ,\PWM4/n26 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub1/u4  (
    .a(pnumcnt4[4]),
    .b(1'b0),
    .c(\PWM4/sub1/c4 ),
    .o({\PWM4/sub1/c5 ,\PWM4/n26 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub1/u5  (
    .a(pnumcnt4[5]),
    .b(1'b0),
    .c(\PWM4/sub1/c5 ),
    .o({\PWM4/sub1/c6 ,\PWM4/n26 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub1/u6  (
    .a(pnumcnt4[6]),
    .b(1'b0),
    .c(\PWM4/sub1/c6 ),
    .o({\PWM4/sub1/c7 ,\PWM4/n26 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub1/u7  (
    .a(pnumcnt4[7]),
    .b(1'b0),
    .c(\PWM4/sub1/c7 ),
    .o({\PWM4/sub1/c8 ,\PWM4/n26 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub1/u8  (
    .a(pnumcnt4[8]),
    .b(1'b0),
    .c(\PWM4/sub1/c8 ),
    .o({\PWM4/sub1/c9 ,\PWM4/n26 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM4/sub1/u9  (
    .a(pnumcnt4[9]),
    .b(1'b0),
    .c(\PWM4/sub1/c9 ),
    .o({\PWM4/sub1/c10 ,\PWM4/n26 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \PWM4/sub1/ucin  (
    .a(1'b0),
    .o({\PWM4/sub1/c0 ,open_n39}));
  reg_ar_as_w1 \PWM5/State_reg  (
    .clk(clk100m),
    .d(\PWM5/n10 ),
    .en(1'b1),
    .reset(~rstn),
    .set(1'b0),
    .q(pwm_state_read[5]));  // src/OnePWM.v(26)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[0]  (
    .i(\PWM5/RemaTxNum[0]_keep ),
    .o(pnumcnt5[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[10]  (
    .i(\PWM5/RemaTxNum[10]_keep ),
    .o(pnumcnt5[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[11]  (
    .i(\PWM5/RemaTxNum[11]_keep ),
    .o(pnumcnt5[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[12]  (
    .i(\PWM5/RemaTxNum[12]_keep ),
    .o(pnumcnt5[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[13]  (
    .i(\PWM5/RemaTxNum[13]_keep ),
    .o(pnumcnt5[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[14]  (
    .i(\PWM5/RemaTxNum[14]_keep ),
    .o(pnumcnt5[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[15]  (
    .i(\PWM5/RemaTxNum[15]_keep ),
    .o(pnumcnt5[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[16]  (
    .i(\PWM5/RemaTxNum[16]_keep ),
    .o(pnumcnt5[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[17]  (
    .i(\PWM5/RemaTxNum[17]_keep ),
    .o(pnumcnt5[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[18]  (
    .i(\PWM5/RemaTxNum[18]_keep ),
    .o(pnumcnt5[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[19]  (
    .i(\PWM5/RemaTxNum[19]_keep ),
    .o(pnumcnt5[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[1]  (
    .i(\PWM5/RemaTxNum[1]_keep ),
    .o(pnumcnt5[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[20]  (
    .i(\PWM5/RemaTxNum[20]_keep ),
    .o(pnumcnt5[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[21]  (
    .i(\PWM5/RemaTxNum[21]_keep ),
    .o(pnumcnt5[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[22]  (
    .i(\PWM5/RemaTxNum[22]_keep ),
    .o(pnumcnt5[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[23]  (
    .i(\PWM5/RemaTxNum[23]_keep ),
    .o(pnumcnt5[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[2]  (
    .i(\PWM5/RemaTxNum[2]_keep ),
    .o(pnumcnt5[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[3]  (
    .i(\PWM5/RemaTxNum[3]_keep ),
    .o(pnumcnt5[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[4]  (
    .i(\PWM5/RemaTxNum[4]_keep ),
    .o(pnumcnt5[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[5]  (
    .i(\PWM5/RemaTxNum[5]_keep ),
    .o(pnumcnt5[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[6]  (
    .i(\PWM5/RemaTxNum[6]_keep ),
    .o(pnumcnt5[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[7]  (
    .i(\PWM5/RemaTxNum[7]_keep ),
    .o(pnumcnt5[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[8]  (
    .i(\PWM5/RemaTxNum[8]_keep ),
    .o(pnumcnt5[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[9]  (
    .i(\PWM5/RemaTxNum[9]_keep ),
    .o(pnumcnt5[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_dir  (
    .i(\PWM5/dir_keep ),
    .o(dir_pad[5]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[0]  (
    .i(\PWM5/pnumr[0]_keep ),
    .o(\PWM5/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[10]  (
    .i(\PWM5/pnumr[10]_keep ),
    .o(\PWM5/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[11]  (
    .i(\PWM5/pnumr[11]_keep ),
    .o(\PWM5/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[12]  (
    .i(\PWM5/pnumr[12]_keep ),
    .o(\PWM5/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[13]  (
    .i(\PWM5/pnumr[13]_keep ),
    .o(\PWM5/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[14]  (
    .i(\PWM5/pnumr[14]_keep ),
    .o(\PWM5/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[15]  (
    .i(\PWM5/pnumr[15]_keep ),
    .o(\PWM5/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[16]  (
    .i(\PWM5/pnumr[16]_keep ),
    .o(\PWM5/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[17]  (
    .i(\PWM5/pnumr[17]_keep ),
    .o(\PWM5/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[18]  (
    .i(\PWM5/pnumr[18]_keep ),
    .o(\PWM5/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[19]  (
    .i(\PWM5/pnumr[19]_keep ),
    .o(\PWM5/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[1]  (
    .i(\PWM5/pnumr[1]_keep ),
    .o(\PWM5/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[20]  (
    .i(\PWM5/pnumr[20]_keep ),
    .o(\PWM5/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[21]  (
    .i(\PWM5/pnumr[21]_keep ),
    .o(\PWM5/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[22]  (
    .i(\PWM5/pnumr[22]_keep ),
    .o(\PWM5/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[23]  (
    .i(\PWM5/pnumr[23]_keep ),
    .o(\PWM5/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[24]  (
    .i(\PWM5/pnumr[24]_keep ),
    .o(\PWM5/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[25]  (
    .i(\PWM5/pnumr[25]_keep ),
    .o(\PWM5/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[26]  (
    .i(\PWM5/pnumr[26]_keep ),
    .o(\PWM5/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[27]  (
    .i(\PWM5/pnumr[27]_keep ),
    .o(\PWM5/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[28]  (
    .i(\PWM5/pnumr[28]_keep ),
    .o(\PWM5/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[29]  (
    .i(\PWM5/pnumr[29]_keep ),
    .o(\PWM5/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[2]  (
    .i(\PWM5/pnumr[2]_keep ),
    .o(\PWM5/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[30]  (
    .i(\PWM5/pnumr[30]_keep ),
    .o(\PWM5/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[31]  (
    .i(\PWM5/pnumr[31]_keep ),
    .o(\PWM5/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[3]  (
    .i(\PWM5/pnumr[3]_keep ),
    .o(\PWM5/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[4]  (
    .i(\PWM5/pnumr[4]_keep ),
    .o(\PWM5/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[5]  (
    .i(\PWM5/pnumr[5]_keep ),
    .o(\PWM5/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[6]  (
    .i(\PWM5/pnumr[6]_keep ),
    .o(\PWM5/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[7]  (
    .i(\PWM5/pnumr[7]_keep ),
    .o(\PWM5/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[8]  (
    .i(\PWM5/pnumr[8]_keep ),
    .o(\PWM5/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[9]  (
    .i(\PWM5/pnumr[9]_keep ),
    .o(\PWM5/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pwm  (
    .i(\PWM5/pwm_keep ),
    .o(pwm_pad[5]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_stopreq  (
    .i(\PWM5/stopreq_keep ),
    .o(\PWM5/stopreq ));  // src/OnePWM.v(14)
  reg_ar_as_w1 \PWM5/dir_reg  (
    .clk(clk100m),
    .d(\PWM5/n32 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/dir_keep ));  // src/OnePWM.v(58)
  reg_sr_as_w1 \PWM5/pwm_reg  (
    .clk(clk100m),
    .d(\pwm[5]_d ),
    .en(1'b1),
    .reset(~\PWM5/u14_sel_is_1_o ),
    .set(1'b0),
    .q(\PWM5/pwm_keep ));  // src/OnePWM.v(45)
  reg_sr_as_w1 \PWM5/reg0_b0  (
    .clk(clk100m),
    .d(\PWM5/n13 [0]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [0]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b1  (
    .clk(clk100m),
    .d(\PWM5/n13 [1]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [1]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b10  (
    .clk(clk100m),
    .d(\PWM5/n13 [10]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [10]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b11  (
    .clk(clk100m),
    .d(\PWM5/n13 [11]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [11]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b12  (
    .clk(clk100m),
    .d(\PWM5/n13 [12]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [12]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b13  (
    .clk(clk100m),
    .d(\PWM5/n13 [13]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [13]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b14  (
    .clk(clk100m),
    .d(\PWM5/n13 [14]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [14]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b15  (
    .clk(clk100m),
    .d(\PWM5/n13 [15]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [15]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b16  (
    .clk(clk100m),
    .d(\PWM5/n13 [16]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [16]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b17  (
    .clk(clk100m),
    .d(\PWM5/n13 [17]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [17]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b18  (
    .clk(clk100m),
    .d(\PWM5/n13 [18]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [18]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b19  (
    .clk(clk100m),
    .d(\PWM5/n13 [19]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [19]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b2  (
    .clk(clk100m),
    .d(\PWM5/n13 [2]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [2]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b20  (
    .clk(clk100m),
    .d(\PWM5/n13 [20]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [20]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b21  (
    .clk(clk100m),
    .d(\PWM5/n13 [21]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [21]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b22  (
    .clk(clk100m),
    .d(\PWM5/n13 [22]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [22]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b23  (
    .clk(clk100m),
    .d(\PWM5/n13 [23]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [23]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b24  (
    .clk(clk100m),
    .d(\PWM5/n13 [24]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [24]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b25  (
    .clk(clk100m),
    .d(\PWM5/n13 [25]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [25]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b26  (
    .clk(clk100m),
    .d(\PWM5/n13 [26]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [26]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b3  (
    .clk(clk100m),
    .d(\PWM5/n13 [3]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [3]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b4  (
    .clk(clk100m),
    .d(\PWM5/n13 [4]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [4]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b5  (
    .clk(clk100m),
    .d(\PWM5/n13 [5]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [5]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b6  (
    .clk(clk100m),
    .d(\PWM5/n13 [6]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [6]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b7  (
    .clk(clk100m),
    .d(\PWM5/n13 [7]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [7]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b8  (
    .clk(clk100m),
    .d(\PWM5/n13 [8]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [8]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b9  (
    .clk(clk100m),
    .d(\PWM5/n13 [9]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b0  (
    .clk(clk100m),
    .d(freq5[0]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [0]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b1  (
    .clk(clk100m),
    .d(freq5[1]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [1]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b10  (
    .clk(clk100m),
    .d(freq5[10]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [10]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b11  (
    .clk(clk100m),
    .d(freq5[11]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [11]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b12  (
    .clk(clk100m),
    .d(freq5[12]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [12]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b13  (
    .clk(clk100m),
    .d(freq5[13]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [13]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b14  (
    .clk(clk100m),
    .d(freq5[14]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [14]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b15  (
    .clk(clk100m),
    .d(freq5[15]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [15]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b16  (
    .clk(clk100m),
    .d(freq5[16]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [16]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b17  (
    .clk(clk100m),
    .d(freq5[17]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [17]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b18  (
    .clk(clk100m),
    .d(freq5[18]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [18]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b19  (
    .clk(clk100m),
    .d(freq5[19]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [19]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b2  (
    .clk(clk100m),
    .d(freq5[2]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [2]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b20  (
    .clk(clk100m),
    .d(freq5[20]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [20]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b21  (
    .clk(clk100m),
    .d(freq5[21]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [21]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b22  (
    .clk(clk100m),
    .d(freq5[22]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [22]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b23  (
    .clk(clk100m),
    .d(freq5[23]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [23]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b24  (
    .clk(clk100m),
    .d(freq5[24]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [24]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b25  (
    .clk(clk100m),
    .d(freq5[25]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [25]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b26  (
    .clk(clk100m),
    .d(freq5[26]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [26]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b3  (
    .clk(clk100m),
    .d(freq5[3]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [3]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b4  (
    .clk(clk100m),
    .d(freq5[4]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [4]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b5  (
    .clk(clk100m),
    .d(freq5[5]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [5]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b6  (
    .clk(clk100m),
    .d(freq5[6]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [6]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b7  (
    .clk(clk100m),
    .d(freq5[7]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [7]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b8  (
    .clk(clk100m),
    .d(freq5[8]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [8]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b9  (
    .clk(clk100m),
    .d(freq5[9]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg2_b0  (
    .clk(clk100m),
    .d(\PWM5/n23 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[0]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b1  (
    .clk(clk100m),
    .d(\PWM5/n23 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[1]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b10  (
    .clk(clk100m),
    .d(\PWM5/n23 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[10]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b11  (
    .clk(clk100m),
    .d(\PWM5/n23 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[11]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b12  (
    .clk(clk100m),
    .d(\PWM5/n23 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[12]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b13  (
    .clk(clk100m),
    .d(\PWM5/n23 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[13]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b14  (
    .clk(clk100m),
    .d(\PWM5/n23 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[14]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b15  (
    .clk(clk100m),
    .d(\PWM5/n23 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[15]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b16  (
    .clk(clk100m),
    .d(\PWM5/n23 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[16]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b17  (
    .clk(clk100m),
    .d(\PWM5/n23 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[17]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b18  (
    .clk(clk100m),
    .d(\PWM5/n23 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[18]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b19  (
    .clk(clk100m),
    .d(\PWM5/n23 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[19]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b2  (
    .clk(clk100m),
    .d(\PWM5/n23 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[2]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b20  (
    .clk(clk100m),
    .d(\PWM5/n23 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[20]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b21  (
    .clk(clk100m),
    .d(\PWM5/n23 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[21]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b22  (
    .clk(clk100m),
    .d(\PWM5/n23 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[22]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b23  (
    .clk(clk100m),
    .d(\PWM5/n23 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[23]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b24  (
    .clk(clk100m),
    .d(\PWM5/n23 [24]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[24]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b25  (
    .clk(clk100m),
    .d(\PWM5/n23 [25]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[25]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b26  (
    .clk(clk100m),
    .d(\PWM5/n23 [26]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[26]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b27  (
    .clk(clk100m),
    .d(\PWM5/n23 [27]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[27]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b28  (
    .clk(clk100m),
    .d(\PWM5/n23 [28]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[28]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b29  (
    .clk(clk100m),
    .d(\PWM5/n23 [29]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[29]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b3  (
    .clk(clk100m),
    .d(\PWM5/n23 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[3]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b30  (
    .clk(clk100m),
    .d(\PWM5/n23 [30]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[30]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b31  (
    .clk(clk100m),
    .d(\PWM5/n23 [31]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[31]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b4  (
    .clk(clk100m),
    .d(\PWM5/n23 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[4]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b5  (
    .clk(clk100m),
    .d(\PWM5/n23 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[5]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b6  (
    .clk(clk100m),
    .d(\PWM5/n23 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[6]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b7  (
    .clk(clk100m),
    .d(\PWM5/n23 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[7]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b8  (
    .clk(clk100m),
    .d(\PWM5/n23 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[8]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b9  (
    .clk(clk100m),
    .d(\PWM5/n23 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[9]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg3_b0  (
    .clk(clk100m),
    .d(\PWM5/n31 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[0]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b1  (
    .clk(clk100m),
    .d(\PWM5/n31 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[1]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b10  (
    .clk(clk100m),
    .d(\PWM5/n31 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[10]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b11  (
    .clk(clk100m),
    .d(\PWM5/n31 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[11]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b12  (
    .clk(clk100m),
    .d(\PWM5/n31 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[12]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b13  (
    .clk(clk100m),
    .d(\PWM5/n31 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[13]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b14  (
    .clk(clk100m),
    .d(\PWM5/n31 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[14]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b15  (
    .clk(clk100m),
    .d(\PWM5/n31 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[15]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b16  (
    .clk(clk100m),
    .d(\PWM5/n31 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[16]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b17  (
    .clk(clk100m),
    .d(\PWM5/n31 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[17]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b18  (
    .clk(clk100m),
    .d(\PWM5/n31 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[18]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b19  (
    .clk(clk100m),
    .d(\PWM5/n31 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[19]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b2  (
    .clk(clk100m),
    .d(\PWM5/n31 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[2]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b20  (
    .clk(clk100m),
    .d(\PWM5/n31 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[20]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b21  (
    .clk(clk100m),
    .d(\PWM5/n31 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[21]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b22  (
    .clk(clk100m),
    .d(\PWM5/n31 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[22]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b23  (
    .clk(clk100m),
    .d(\PWM5/n31 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[23]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b3  (
    .clk(clk100m),
    .d(\PWM5/n31 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[3]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b4  (
    .clk(clk100m),
    .d(\PWM5/n31 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[4]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b5  (
    .clk(clk100m),
    .d(\PWM5/n31 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[5]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b6  (
    .clk(clk100m),
    .d(\PWM5/n31 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[6]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b7  (
    .clk(clk100m),
    .d(\PWM5/n31 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[7]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b8  (
    .clk(clk100m),
    .d(\PWM5/n31 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[8]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b9  (
    .clk(clk100m),
    .d(\PWM5/n31 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[9]_keep ));  // src/OnePWM.v(58)
  reg_ar_ss_w1 \PWM5/stopreq_reg  (
    .clk(clk100m),
    .d(\PWM5/n1 ),
    .en(1'b1),
    .reset(1'b0),
    .set(pwm_start_stop[5]),
    .q(\PWM5/stopreq_keep ));  // src/OnePWM.v(15)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub0/u0  (
    .a(\PWM5/FreCnt [0]),
    .b(1'b1),
    .c(\PWM5/sub0/c0 ),
    .o({\PWM5/sub0/c1 ,\PWM5/n12 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub0/u1  (
    .a(\PWM5/FreCnt [1]),
    .b(1'b0),
    .c(\PWM5/sub0/c1 ),
    .o({\PWM5/sub0/c2 ,\PWM5/n12 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub0/u10  (
    .a(\PWM5/FreCnt [10]),
    .b(1'b0),
    .c(\PWM5/sub0/c10 ),
    .o({\PWM5/sub0/c11 ,\PWM5/n12 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub0/u11  (
    .a(\PWM5/FreCnt [11]),
    .b(1'b0),
    .c(\PWM5/sub0/c11 ),
    .o({\PWM5/sub0/c12 ,\PWM5/n12 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub0/u12  (
    .a(\PWM5/FreCnt [12]),
    .b(1'b0),
    .c(\PWM5/sub0/c12 ),
    .o({\PWM5/sub0/c13 ,\PWM5/n12 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub0/u13  (
    .a(\PWM5/FreCnt [13]),
    .b(1'b0),
    .c(\PWM5/sub0/c13 ),
    .o({\PWM5/sub0/c14 ,\PWM5/n12 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub0/u14  (
    .a(\PWM5/FreCnt [14]),
    .b(1'b0),
    .c(\PWM5/sub0/c14 ),
    .o({\PWM5/sub0/c15 ,\PWM5/n12 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub0/u15  (
    .a(\PWM5/FreCnt [15]),
    .b(1'b0),
    .c(\PWM5/sub0/c15 ),
    .o({\PWM5/sub0/c16 ,\PWM5/n12 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub0/u16  (
    .a(\PWM5/FreCnt [16]),
    .b(1'b0),
    .c(\PWM5/sub0/c16 ),
    .o({\PWM5/sub0/c17 ,\PWM5/n12 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub0/u17  (
    .a(\PWM5/FreCnt [17]),
    .b(1'b0),
    .c(\PWM5/sub0/c17 ),
    .o({\PWM5/sub0/c18 ,\PWM5/n12 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub0/u18  (
    .a(\PWM5/FreCnt [18]),
    .b(1'b0),
    .c(\PWM5/sub0/c18 ),
    .o({\PWM5/sub0/c19 ,\PWM5/n12 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub0/u19  (
    .a(\PWM5/FreCnt [19]),
    .b(1'b0),
    .c(\PWM5/sub0/c19 ),
    .o({\PWM5/sub0/c20 ,\PWM5/n12 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub0/u2  (
    .a(\PWM5/FreCnt [2]),
    .b(1'b0),
    .c(\PWM5/sub0/c2 ),
    .o({\PWM5/sub0/c3 ,\PWM5/n12 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub0/u20  (
    .a(\PWM5/FreCnt [20]),
    .b(1'b0),
    .c(\PWM5/sub0/c20 ),
    .o({\PWM5/sub0/c21 ,\PWM5/n12 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub0/u21  (
    .a(\PWM5/FreCnt [21]),
    .b(1'b0),
    .c(\PWM5/sub0/c21 ),
    .o({\PWM5/sub0/c22 ,\PWM5/n12 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub0/u22  (
    .a(\PWM5/FreCnt [22]),
    .b(1'b0),
    .c(\PWM5/sub0/c22 ),
    .o({\PWM5/sub0/c23 ,\PWM5/n12 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub0/u23  (
    .a(\PWM5/FreCnt [23]),
    .b(1'b0),
    .c(\PWM5/sub0/c23 ),
    .o({\PWM5/sub0/c24 ,\PWM5/n12 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub0/u24  (
    .a(\PWM5/FreCnt [24]),
    .b(1'b0),
    .c(\PWM5/sub0/c24 ),
    .o({\PWM5/sub0/c25 ,\PWM5/n12 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub0/u25  (
    .a(\PWM5/FreCnt [25]),
    .b(1'b0),
    .c(\PWM5/sub0/c25 ),
    .o({\PWM5/sub0/c26 ,\PWM5/n12 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub0/u26  (
    .a(\PWM5/FreCnt [26]),
    .b(1'b0),
    .c(\PWM5/sub0/c26 ),
    .o({open_n40,\PWM5/n12 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub0/u3  (
    .a(\PWM5/FreCnt [3]),
    .b(1'b0),
    .c(\PWM5/sub0/c3 ),
    .o({\PWM5/sub0/c4 ,\PWM5/n12 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub0/u4  (
    .a(\PWM5/FreCnt [4]),
    .b(1'b0),
    .c(\PWM5/sub0/c4 ),
    .o({\PWM5/sub0/c5 ,\PWM5/n12 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub0/u5  (
    .a(\PWM5/FreCnt [5]),
    .b(1'b0),
    .c(\PWM5/sub0/c5 ),
    .o({\PWM5/sub0/c6 ,\PWM5/n12 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub0/u6  (
    .a(\PWM5/FreCnt [6]),
    .b(1'b0),
    .c(\PWM5/sub0/c6 ),
    .o({\PWM5/sub0/c7 ,\PWM5/n12 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub0/u7  (
    .a(\PWM5/FreCnt [7]),
    .b(1'b0),
    .c(\PWM5/sub0/c7 ),
    .o({\PWM5/sub0/c8 ,\PWM5/n12 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub0/u8  (
    .a(\PWM5/FreCnt [8]),
    .b(1'b0),
    .c(\PWM5/sub0/c8 ),
    .o({\PWM5/sub0/c9 ,\PWM5/n12 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub0/u9  (
    .a(\PWM5/FreCnt [9]),
    .b(1'b0),
    .c(\PWM5/sub0/c9 ),
    .o({\PWM5/sub0/c10 ,\PWM5/n12 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \PWM5/sub0/ucin  (
    .a(1'b0),
    .o({\PWM5/sub0/c0 ,open_n43}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub1/u0  (
    .a(pnumcnt5[0]),
    .b(1'b1),
    .c(\PWM5/sub1/c0 ),
    .o({\PWM5/sub1/c1 ,\PWM5/n26 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub1/u1  (
    .a(pnumcnt5[1]),
    .b(1'b0),
    .c(\PWM5/sub1/c1 ),
    .o({\PWM5/sub1/c2 ,\PWM5/n26 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub1/u10  (
    .a(pnumcnt5[10]),
    .b(1'b0),
    .c(\PWM5/sub1/c10 ),
    .o({\PWM5/sub1/c11 ,\PWM5/n26 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub1/u11  (
    .a(pnumcnt5[11]),
    .b(1'b0),
    .c(\PWM5/sub1/c11 ),
    .o({\PWM5/sub1/c12 ,\PWM5/n26 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub1/u12  (
    .a(pnumcnt5[12]),
    .b(1'b0),
    .c(\PWM5/sub1/c12 ),
    .o({\PWM5/sub1/c13 ,\PWM5/n26 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub1/u13  (
    .a(pnumcnt5[13]),
    .b(1'b0),
    .c(\PWM5/sub1/c13 ),
    .o({\PWM5/sub1/c14 ,\PWM5/n26 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub1/u14  (
    .a(pnumcnt5[14]),
    .b(1'b0),
    .c(\PWM5/sub1/c14 ),
    .o({\PWM5/sub1/c15 ,\PWM5/n26 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub1/u15  (
    .a(pnumcnt5[15]),
    .b(1'b0),
    .c(\PWM5/sub1/c15 ),
    .o({\PWM5/sub1/c16 ,\PWM5/n26 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub1/u16  (
    .a(pnumcnt5[16]),
    .b(1'b0),
    .c(\PWM5/sub1/c16 ),
    .o({\PWM5/sub1/c17 ,\PWM5/n26 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub1/u17  (
    .a(pnumcnt5[17]),
    .b(1'b0),
    .c(\PWM5/sub1/c17 ),
    .o({\PWM5/sub1/c18 ,\PWM5/n26 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub1/u18  (
    .a(pnumcnt5[18]),
    .b(1'b0),
    .c(\PWM5/sub1/c18 ),
    .o({\PWM5/sub1/c19 ,\PWM5/n26 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub1/u19  (
    .a(pnumcnt5[19]),
    .b(1'b0),
    .c(\PWM5/sub1/c19 ),
    .o({\PWM5/sub1/c20 ,\PWM5/n26 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub1/u2  (
    .a(pnumcnt5[2]),
    .b(1'b0),
    .c(\PWM5/sub1/c2 ),
    .o({\PWM5/sub1/c3 ,\PWM5/n26 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub1/u20  (
    .a(pnumcnt5[20]),
    .b(1'b0),
    .c(\PWM5/sub1/c20 ),
    .o({\PWM5/sub1/c21 ,\PWM5/n26 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub1/u21  (
    .a(pnumcnt5[21]),
    .b(1'b0),
    .c(\PWM5/sub1/c21 ),
    .o({\PWM5/sub1/c22 ,\PWM5/n26 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub1/u22  (
    .a(pnumcnt5[22]),
    .b(1'b0),
    .c(\PWM5/sub1/c22 ),
    .o({\PWM5/sub1/c23 ,\PWM5/n26 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub1/u23  (
    .a(pnumcnt5[23]),
    .b(1'b0),
    .c(\PWM5/sub1/c23 ),
    .o({open_n44,\PWM5/n26 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub1/u3  (
    .a(pnumcnt5[3]),
    .b(1'b0),
    .c(\PWM5/sub1/c3 ),
    .o({\PWM5/sub1/c4 ,\PWM5/n26 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub1/u4  (
    .a(pnumcnt5[4]),
    .b(1'b0),
    .c(\PWM5/sub1/c4 ),
    .o({\PWM5/sub1/c5 ,\PWM5/n26 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub1/u5  (
    .a(pnumcnt5[5]),
    .b(1'b0),
    .c(\PWM5/sub1/c5 ),
    .o({\PWM5/sub1/c6 ,\PWM5/n26 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub1/u6  (
    .a(pnumcnt5[6]),
    .b(1'b0),
    .c(\PWM5/sub1/c6 ),
    .o({\PWM5/sub1/c7 ,\PWM5/n26 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub1/u7  (
    .a(pnumcnt5[7]),
    .b(1'b0),
    .c(\PWM5/sub1/c7 ),
    .o({\PWM5/sub1/c8 ,\PWM5/n26 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub1/u8  (
    .a(pnumcnt5[8]),
    .b(1'b0),
    .c(\PWM5/sub1/c8 ),
    .o({\PWM5/sub1/c9 ,\PWM5/n26 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM5/sub1/u9  (
    .a(pnumcnt5[9]),
    .b(1'b0),
    .c(\PWM5/sub1/c9 ),
    .o({\PWM5/sub1/c10 ,\PWM5/n26 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \PWM5/sub1/ucin  (
    .a(1'b0),
    .o({\PWM5/sub1/c0 ,open_n47}));
  reg_ar_as_w1 \PWM6/State_reg  (
    .clk(clk100m),
    .d(\PWM6/n10 ),
    .en(1'b1),
    .reset(~rstn),
    .set(1'b0),
    .q(pwm_state_read[6]));  // src/OnePWM.v(26)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[0]  (
    .i(\PWM6/RemaTxNum[0]_keep ),
    .o(pnumcnt6[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[10]  (
    .i(\PWM6/RemaTxNum[10]_keep ),
    .o(pnumcnt6[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[11]  (
    .i(\PWM6/RemaTxNum[11]_keep ),
    .o(pnumcnt6[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[12]  (
    .i(\PWM6/RemaTxNum[12]_keep ),
    .o(pnumcnt6[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[13]  (
    .i(\PWM6/RemaTxNum[13]_keep ),
    .o(pnumcnt6[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[14]  (
    .i(\PWM6/RemaTxNum[14]_keep ),
    .o(pnumcnt6[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[15]  (
    .i(\PWM6/RemaTxNum[15]_keep ),
    .o(pnumcnt6[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[16]  (
    .i(\PWM6/RemaTxNum[16]_keep ),
    .o(pnumcnt6[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[17]  (
    .i(\PWM6/RemaTxNum[17]_keep ),
    .o(pnumcnt6[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[18]  (
    .i(\PWM6/RemaTxNum[18]_keep ),
    .o(pnumcnt6[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[19]  (
    .i(\PWM6/RemaTxNum[19]_keep ),
    .o(pnumcnt6[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[1]  (
    .i(\PWM6/RemaTxNum[1]_keep ),
    .o(pnumcnt6[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[20]  (
    .i(\PWM6/RemaTxNum[20]_keep ),
    .o(pnumcnt6[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[21]  (
    .i(\PWM6/RemaTxNum[21]_keep ),
    .o(pnumcnt6[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[22]  (
    .i(\PWM6/RemaTxNum[22]_keep ),
    .o(pnumcnt6[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[23]  (
    .i(\PWM6/RemaTxNum[23]_keep ),
    .o(pnumcnt6[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[2]  (
    .i(\PWM6/RemaTxNum[2]_keep ),
    .o(pnumcnt6[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[3]  (
    .i(\PWM6/RemaTxNum[3]_keep ),
    .o(pnumcnt6[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[4]  (
    .i(\PWM6/RemaTxNum[4]_keep ),
    .o(pnumcnt6[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[5]  (
    .i(\PWM6/RemaTxNum[5]_keep ),
    .o(pnumcnt6[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[6]  (
    .i(\PWM6/RemaTxNum[6]_keep ),
    .o(pnumcnt6[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[7]  (
    .i(\PWM6/RemaTxNum[7]_keep ),
    .o(pnumcnt6[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[8]  (
    .i(\PWM6/RemaTxNum[8]_keep ),
    .o(pnumcnt6[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[9]  (
    .i(\PWM6/RemaTxNum[9]_keep ),
    .o(pnumcnt6[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_dir  (
    .i(\PWM6/dir_keep ),
    .o(dir_pad[6]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[0]  (
    .i(\PWM6/pnumr[0]_keep ),
    .o(\PWM6/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[10]  (
    .i(\PWM6/pnumr[10]_keep ),
    .o(\PWM6/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[11]  (
    .i(\PWM6/pnumr[11]_keep ),
    .o(\PWM6/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[12]  (
    .i(\PWM6/pnumr[12]_keep ),
    .o(\PWM6/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[13]  (
    .i(\PWM6/pnumr[13]_keep ),
    .o(\PWM6/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[14]  (
    .i(\PWM6/pnumr[14]_keep ),
    .o(\PWM6/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[15]  (
    .i(\PWM6/pnumr[15]_keep ),
    .o(\PWM6/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[16]  (
    .i(\PWM6/pnumr[16]_keep ),
    .o(\PWM6/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[17]  (
    .i(\PWM6/pnumr[17]_keep ),
    .o(\PWM6/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[18]  (
    .i(\PWM6/pnumr[18]_keep ),
    .o(\PWM6/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[19]  (
    .i(\PWM6/pnumr[19]_keep ),
    .o(\PWM6/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[1]  (
    .i(\PWM6/pnumr[1]_keep ),
    .o(\PWM6/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[20]  (
    .i(\PWM6/pnumr[20]_keep ),
    .o(\PWM6/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[21]  (
    .i(\PWM6/pnumr[21]_keep ),
    .o(\PWM6/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[22]  (
    .i(\PWM6/pnumr[22]_keep ),
    .o(\PWM6/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[23]  (
    .i(\PWM6/pnumr[23]_keep ),
    .o(\PWM6/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[24]  (
    .i(\PWM6/pnumr[24]_keep ),
    .o(\PWM6/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[25]  (
    .i(\PWM6/pnumr[25]_keep ),
    .o(\PWM6/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[26]  (
    .i(\PWM6/pnumr[26]_keep ),
    .o(\PWM6/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[27]  (
    .i(\PWM6/pnumr[27]_keep ),
    .o(\PWM6/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[28]  (
    .i(\PWM6/pnumr[28]_keep ),
    .o(\PWM6/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[29]  (
    .i(\PWM6/pnumr[29]_keep ),
    .o(\PWM6/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[2]  (
    .i(\PWM6/pnumr[2]_keep ),
    .o(\PWM6/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[30]  (
    .i(\PWM6/pnumr[30]_keep ),
    .o(\PWM6/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[31]  (
    .i(\PWM6/pnumr[31]_keep ),
    .o(\PWM6/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[3]  (
    .i(\PWM6/pnumr[3]_keep ),
    .o(\PWM6/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[4]  (
    .i(\PWM6/pnumr[4]_keep ),
    .o(\PWM6/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[5]  (
    .i(\PWM6/pnumr[5]_keep ),
    .o(\PWM6/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[6]  (
    .i(\PWM6/pnumr[6]_keep ),
    .o(\PWM6/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[7]  (
    .i(\PWM6/pnumr[7]_keep ),
    .o(\PWM6/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[8]  (
    .i(\PWM6/pnumr[8]_keep ),
    .o(\PWM6/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[9]  (
    .i(\PWM6/pnumr[9]_keep ),
    .o(\PWM6/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pwm  (
    .i(\PWM6/pwm_keep ),
    .o(pwm_pad[6]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_stopreq  (
    .i(\PWM6/stopreq_keep ),
    .o(\PWM6/stopreq ));  // src/OnePWM.v(14)
  reg_ar_as_w1 \PWM6/dir_reg  (
    .clk(clk100m),
    .d(\PWM6/n32 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/dir_keep ));  // src/OnePWM.v(58)
  reg_sr_as_w1 \PWM6/pwm_reg  (
    .clk(clk100m),
    .d(\pwm[6]_d ),
    .en(1'b1),
    .reset(~\PWM6/u14_sel_is_1_o ),
    .set(1'b0),
    .q(\PWM6/pwm_keep ));  // src/OnePWM.v(45)
  reg_sr_as_w1 \PWM6/reg0_b0  (
    .clk(clk100m),
    .d(\PWM6/n13 [0]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [0]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b1  (
    .clk(clk100m),
    .d(\PWM6/n13 [1]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [1]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b10  (
    .clk(clk100m),
    .d(\PWM6/n13 [10]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [10]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b11  (
    .clk(clk100m),
    .d(\PWM6/n13 [11]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [11]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b12  (
    .clk(clk100m),
    .d(\PWM6/n13 [12]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [12]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b13  (
    .clk(clk100m),
    .d(\PWM6/n13 [13]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [13]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b14  (
    .clk(clk100m),
    .d(\PWM6/n13 [14]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [14]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b15  (
    .clk(clk100m),
    .d(\PWM6/n13 [15]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [15]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b16  (
    .clk(clk100m),
    .d(\PWM6/n13 [16]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [16]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b17  (
    .clk(clk100m),
    .d(\PWM6/n13 [17]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [17]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b18  (
    .clk(clk100m),
    .d(\PWM6/n13 [18]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [18]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b19  (
    .clk(clk100m),
    .d(\PWM6/n13 [19]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [19]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b2  (
    .clk(clk100m),
    .d(\PWM6/n13 [2]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [2]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b20  (
    .clk(clk100m),
    .d(\PWM6/n13 [20]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [20]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b21  (
    .clk(clk100m),
    .d(\PWM6/n13 [21]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [21]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b22  (
    .clk(clk100m),
    .d(\PWM6/n13 [22]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [22]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b23  (
    .clk(clk100m),
    .d(\PWM6/n13 [23]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [23]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b24  (
    .clk(clk100m),
    .d(\PWM6/n13 [24]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [24]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b25  (
    .clk(clk100m),
    .d(\PWM6/n13 [25]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [25]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b26  (
    .clk(clk100m),
    .d(\PWM6/n13 [26]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [26]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b3  (
    .clk(clk100m),
    .d(\PWM6/n13 [3]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [3]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b4  (
    .clk(clk100m),
    .d(\PWM6/n13 [4]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [4]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b5  (
    .clk(clk100m),
    .d(\PWM6/n13 [5]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [5]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b6  (
    .clk(clk100m),
    .d(\PWM6/n13 [6]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [6]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b7  (
    .clk(clk100m),
    .d(\PWM6/n13 [7]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [7]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b8  (
    .clk(clk100m),
    .d(\PWM6/n13 [8]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [8]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b9  (
    .clk(clk100m),
    .d(\PWM6/n13 [9]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b0  (
    .clk(clk100m),
    .d(freq6[0]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [0]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b1  (
    .clk(clk100m),
    .d(freq6[1]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [1]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b10  (
    .clk(clk100m),
    .d(freq6[10]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [10]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b11  (
    .clk(clk100m),
    .d(freq6[11]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [11]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b12  (
    .clk(clk100m),
    .d(freq6[12]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [12]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b13  (
    .clk(clk100m),
    .d(freq6[13]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [13]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b14  (
    .clk(clk100m),
    .d(freq6[14]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [14]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b15  (
    .clk(clk100m),
    .d(freq6[15]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [15]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b16  (
    .clk(clk100m),
    .d(freq6[16]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [16]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b17  (
    .clk(clk100m),
    .d(freq6[17]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [17]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b18  (
    .clk(clk100m),
    .d(freq6[18]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [18]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b19  (
    .clk(clk100m),
    .d(freq6[19]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [19]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b2  (
    .clk(clk100m),
    .d(freq6[2]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [2]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b20  (
    .clk(clk100m),
    .d(freq6[20]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [20]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b21  (
    .clk(clk100m),
    .d(freq6[21]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [21]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b22  (
    .clk(clk100m),
    .d(freq6[22]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [22]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b23  (
    .clk(clk100m),
    .d(freq6[23]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [23]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b24  (
    .clk(clk100m),
    .d(freq6[24]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [24]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b25  (
    .clk(clk100m),
    .d(freq6[25]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [25]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b26  (
    .clk(clk100m),
    .d(freq6[26]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [26]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b3  (
    .clk(clk100m),
    .d(freq6[3]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [3]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b4  (
    .clk(clk100m),
    .d(freq6[4]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [4]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b5  (
    .clk(clk100m),
    .d(freq6[5]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [5]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b6  (
    .clk(clk100m),
    .d(freq6[6]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [6]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b7  (
    .clk(clk100m),
    .d(freq6[7]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [7]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b8  (
    .clk(clk100m),
    .d(freq6[8]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [8]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b9  (
    .clk(clk100m),
    .d(freq6[9]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg2_b0  (
    .clk(clk100m),
    .d(\PWM6/n23 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[0]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b1  (
    .clk(clk100m),
    .d(\PWM6/n23 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[1]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b10  (
    .clk(clk100m),
    .d(\PWM6/n23 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[10]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b11  (
    .clk(clk100m),
    .d(\PWM6/n23 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[11]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b12  (
    .clk(clk100m),
    .d(\PWM6/n23 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[12]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b13  (
    .clk(clk100m),
    .d(\PWM6/n23 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[13]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b14  (
    .clk(clk100m),
    .d(\PWM6/n23 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[14]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b15  (
    .clk(clk100m),
    .d(\PWM6/n23 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[15]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b16  (
    .clk(clk100m),
    .d(\PWM6/n23 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[16]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b17  (
    .clk(clk100m),
    .d(\PWM6/n23 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[17]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b18  (
    .clk(clk100m),
    .d(\PWM6/n23 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[18]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b19  (
    .clk(clk100m),
    .d(\PWM6/n23 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[19]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b2  (
    .clk(clk100m),
    .d(\PWM6/n23 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[2]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b20  (
    .clk(clk100m),
    .d(\PWM6/n23 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[20]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b21  (
    .clk(clk100m),
    .d(\PWM6/n23 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[21]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b22  (
    .clk(clk100m),
    .d(\PWM6/n23 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[22]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b23  (
    .clk(clk100m),
    .d(\PWM6/n23 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[23]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b24  (
    .clk(clk100m),
    .d(\PWM6/n23 [24]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[24]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b25  (
    .clk(clk100m),
    .d(\PWM6/n23 [25]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[25]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b26  (
    .clk(clk100m),
    .d(\PWM6/n23 [26]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[26]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b27  (
    .clk(clk100m),
    .d(\PWM6/n23 [27]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[27]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b28  (
    .clk(clk100m),
    .d(\PWM6/n23 [28]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[28]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b29  (
    .clk(clk100m),
    .d(\PWM6/n23 [29]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[29]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b3  (
    .clk(clk100m),
    .d(\PWM6/n23 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[3]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b30  (
    .clk(clk100m),
    .d(\PWM6/n23 [30]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[30]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b31  (
    .clk(clk100m),
    .d(\PWM6/n23 [31]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[31]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b4  (
    .clk(clk100m),
    .d(\PWM6/n23 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[4]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b5  (
    .clk(clk100m),
    .d(\PWM6/n23 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[5]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b6  (
    .clk(clk100m),
    .d(\PWM6/n23 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[6]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b7  (
    .clk(clk100m),
    .d(\PWM6/n23 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[7]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b8  (
    .clk(clk100m),
    .d(\PWM6/n23 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[8]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b9  (
    .clk(clk100m),
    .d(\PWM6/n23 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[9]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg3_b0  (
    .clk(clk100m),
    .d(\PWM6/n31 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[0]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b1  (
    .clk(clk100m),
    .d(\PWM6/n31 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[1]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b10  (
    .clk(clk100m),
    .d(\PWM6/n31 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[10]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b11  (
    .clk(clk100m),
    .d(\PWM6/n31 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[11]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b12  (
    .clk(clk100m),
    .d(\PWM6/n31 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[12]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b13  (
    .clk(clk100m),
    .d(\PWM6/n31 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[13]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b14  (
    .clk(clk100m),
    .d(\PWM6/n31 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[14]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b15  (
    .clk(clk100m),
    .d(\PWM6/n31 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[15]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b16  (
    .clk(clk100m),
    .d(\PWM6/n31 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[16]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b17  (
    .clk(clk100m),
    .d(\PWM6/n31 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[17]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b18  (
    .clk(clk100m),
    .d(\PWM6/n31 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[18]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b19  (
    .clk(clk100m),
    .d(\PWM6/n31 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[19]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b2  (
    .clk(clk100m),
    .d(\PWM6/n31 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[2]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b20  (
    .clk(clk100m),
    .d(\PWM6/n31 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[20]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b21  (
    .clk(clk100m),
    .d(\PWM6/n31 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[21]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b22  (
    .clk(clk100m),
    .d(\PWM6/n31 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[22]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b23  (
    .clk(clk100m),
    .d(\PWM6/n31 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[23]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b3  (
    .clk(clk100m),
    .d(\PWM6/n31 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[3]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b4  (
    .clk(clk100m),
    .d(\PWM6/n31 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[4]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b5  (
    .clk(clk100m),
    .d(\PWM6/n31 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[5]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b6  (
    .clk(clk100m),
    .d(\PWM6/n31 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[6]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b7  (
    .clk(clk100m),
    .d(\PWM6/n31 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[7]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b8  (
    .clk(clk100m),
    .d(\PWM6/n31 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[8]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b9  (
    .clk(clk100m),
    .d(\PWM6/n31 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[9]_keep ));  // src/OnePWM.v(58)
  reg_ar_ss_w1 \PWM6/stopreq_reg  (
    .clk(clk100m),
    .d(\PWM6/n1 ),
    .en(1'b1),
    .reset(1'b0),
    .set(pwm_start_stop[6]),
    .q(\PWM6/stopreq_keep ));  // src/OnePWM.v(15)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub0/u0  (
    .a(\PWM6/FreCnt [0]),
    .b(1'b1),
    .c(\PWM6/sub0/c0 ),
    .o({\PWM6/sub0/c1 ,\PWM6/n12 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub0/u1  (
    .a(\PWM6/FreCnt [1]),
    .b(1'b0),
    .c(\PWM6/sub0/c1 ),
    .o({\PWM6/sub0/c2 ,\PWM6/n12 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub0/u10  (
    .a(\PWM6/FreCnt [10]),
    .b(1'b0),
    .c(\PWM6/sub0/c10 ),
    .o({\PWM6/sub0/c11 ,\PWM6/n12 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub0/u11  (
    .a(\PWM6/FreCnt [11]),
    .b(1'b0),
    .c(\PWM6/sub0/c11 ),
    .o({\PWM6/sub0/c12 ,\PWM6/n12 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub0/u12  (
    .a(\PWM6/FreCnt [12]),
    .b(1'b0),
    .c(\PWM6/sub0/c12 ),
    .o({\PWM6/sub0/c13 ,\PWM6/n12 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub0/u13  (
    .a(\PWM6/FreCnt [13]),
    .b(1'b0),
    .c(\PWM6/sub0/c13 ),
    .o({\PWM6/sub0/c14 ,\PWM6/n12 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub0/u14  (
    .a(\PWM6/FreCnt [14]),
    .b(1'b0),
    .c(\PWM6/sub0/c14 ),
    .o({\PWM6/sub0/c15 ,\PWM6/n12 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub0/u15  (
    .a(\PWM6/FreCnt [15]),
    .b(1'b0),
    .c(\PWM6/sub0/c15 ),
    .o({\PWM6/sub0/c16 ,\PWM6/n12 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub0/u16  (
    .a(\PWM6/FreCnt [16]),
    .b(1'b0),
    .c(\PWM6/sub0/c16 ),
    .o({\PWM6/sub0/c17 ,\PWM6/n12 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub0/u17  (
    .a(\PWM6/FreCnt [17]),
    .b(1'b0),
    .c(\PWM6/sub0/c17 ),
    .o({\PWM6/sub0/c18 ,\PWM6/n12 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub0/u18  (
    .a(\PWM6/FreCnt [18]),
    .b(1'b0),
    .c(\PWM6/sub0/c18 ),
    .o({\PWM6/sub0/c19 ,\PWM6/n12 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub0/u19  (
    .a(\PWM6/FreCnt [19]),
    .b(1'b0),
    .c(\PWM6/sub0/c19 ),
    .o({\PWM6/sub0/c20 ,\PWM6/n12 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub0/u2  (
    .a(\PWM6/FreCnt [2]),
    .b(1'b0),
    .c(\PWM6/sub0/c2 ),
    .o({\PWM6/sub0/c3 ,\PWM6/n12 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub0/u20  (
    .a(\PWM6/FreCnt [20]),
    .b(1'b0),
    .c(\PWM6/sub0/c20 ),
    .o({\PWM6/sub0/c21 ,\PWM6/n12 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub0/u21  (
    .a(\PWM6/FreCnt [21]),
    .b(1'b0),
    .c(\PWM6/sub0/c21 ),
    .o({\PWM6/sub0/c22 ,\PWM6/n12 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub0/u22  (
    .a(\PWM6/FreCnt [22]),
    .b(1'b0),
    .c(\PWM6/sub0/c22 ),
    .o({\PWM6/sub0/c23 ,\PWM6/n12 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub0/u23  (
    .a(\PWM6/FreCnt [23]),
    .b(1'b0),
    .c(\PWM6/sub0/c23 ),
    .o({\PWM6/sub0/c24 ,\PWM6/n12 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub0/u24  (
    .a(\PWM6/FreCnt [24]),
    .b(1'b0),
    .c(\PWM6/sub0/c24 ),
    .o({\PWM6/sub0/c25 ,\PWM6/n12 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub0/u25  (
    .a(\PWM6/FreCnt [25]),
    .b(1'b0),
    .c(\PWM6/sub0/c25 ),
    .o({\PWM6/sub0/c26 ,\PWM6/n12 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub0/u26  (
    .a(\PWM6/FreCnt [26]),
    .b(1'b0),
    .c(\PWM6/sub0/c26 ),
    .o({open_n48,\PWM6/n12 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub0/u3  (
    .a(\PWM6/FreCnt [3]),
    .b(1'b0),
    .c(\PWM6/sub0/c3 ),
    .o({\PWM6/sub0/c4 ,\PWM6/n12 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub0/u4  (
    .a(\PWM6/FreCnt [4]),
    .b(1'b0),
    .c(\PWM6/sub0/c4 ),
    .o({\PWM6/sub0/c5 ,\PWM6/n12 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub0/u5  (
    .a(\PWM6/FreCnt [5]),
    .b(1'b0),
    .c(\PWM6/sub0/c5 ),
    .o({\PWM6/sub0/c6 ,\PWM6/n12 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub0/u6  (
    .a(\PWM6/FreCnt [6]),
    .b(1'b0),
    .c(\PWM6/sub0/c6 ),
    .o({\PWM6/sub0/c7 ,\PWM6/n12 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub0/u7  (
    .a(\PWM6/FreCnt [7]),
    .b(1'b0),
    .c(\PWM6/sub0/c7 ),
    .o({\PWM6/sub0/c8 ,\PWM6/n12 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub0/u8  (
    .a(\PWM6/FreCnt [8]),
    .b(1'b0),
    .c(\PWM6/sub0/c8 ),
    .o({\PWM6/sub0/c9 ,\PWM6/n12 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub0/u9  (
    .a(\PWM6/FreCnt [9]),
    .b(1'b0),
    .c(\PWM6/sub0/c9 ),
    .o({\PWM6/sub0/c10 ,\PWM6/n12 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \PWM6/sub0/ucin  (
    .a(1'b0),
    .o({\PWM6/sub0/c0 ,open_n51}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub1/u0  (
    .a(pnumcnt6[0]),
    .b(1'b1),
    .c(\PWM6/sub1/c0 ),
    .o({\PWM6/sub1/c1 ,\PWM6/n26 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub1/u1  (
    .a(pnumcnt6[1]),
    .b(1'b0),
    .c(\PWM6/sub1/c1 ),
    .o({\PWM6/sub1/c2 ,\PWM6/n26 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub1/u10  (
    .a(pnumcnt6[10]),
    .b(1'b0),
    .c(\PWM6/sub1/c10 ),
    .o({\PWM6/sub1/c11 ,\PWM6/n26 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub1/u11  (
    .a(pnumcnt6[11]),
    .b(1'b0),
    .c(\PWM6/sub1/c11 ),
    .o({\PWM6/sub1/c12 ,\PWM6/n26 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub1/u12  (
    .a(pnumcnt6[12]),
    .b(1'b0),
    .c(\PWM6/sub1/c12 ),
    .o({\PWM6/sub1/c13 ,\PWM6/n26 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub1/u13  (
    .a(pnumcnt6[13]),
    .b(1'b0),
    .c(\PWM6/sub1/c13 ),
    .o({\PWM6/sub1/c14 ,\PWM6/n26 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub1/u14  (
    .a(pnumcnt6[14]),
    .b(1'b0),
    .c(\PWM6/sub1/c14 ),
    .o({\PWM6/sub1/c15 ,\PWM6/n26 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub1/u15  (
    .a(pnumcnt6[15]),
    .b(1'b0),
    .c(\PWM6/sub1/c15 ),
    .o({\PWM6/sub1/c16 ,\PWM6/n26 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub1/u16  (
    .a(pnumcnt6[16]),
    .b(1'b0),
    .c(\PWM6/sub1/c16 ),
    .o({\PWM6/sub1/c17 ,\PWM6/n26 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub1/u17  (
    .a(pnumcnt6[17]),
    .b(1'b0),
    .c(\PWM6/sub1/c17 ),
    .o({\PWM6/sub1/c18 ,\PWM6/n26 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub1/u18  (
    .a(pnumcnt6[18]),
    .b(1'b0),
    .c(\PWM6/sub1/c18 ),
    .o({\PWM6/sub1/c19 ,\PWM6/n26 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub1/u19  (
    .a(pnumcnt6[19]),
    .b(1'b0),
    .c(\PWM6/sub1/c19 ),
    .o({\PWM6/sub1/c20 ,\PWM6/n26 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub1/u2  (
    .a(pnumcnt6[2]),
    .b(1'b0),
    .c(\PWM6/sub1/c2 ),
    .o({\PWM6/sub1/c3 ,\PWM6/n26 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub1/u20  (
    .a(pnumcnt6[20]),
    .b(1'b0),
    .c(\PWM6/sub1/c20 ),
    .o({\PWM6/sub1/c21 ,\PWM6/n26 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub1/u21  (
    .a(pnumcnt6[21]),
    .b(1'b0),
    .c(\PWM6/sub1/c21 ),
    .o({\PWM6/sub1/c22 ,\PWM6/n26 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub1/u22  (
    .a(pnumcnt6[22]),
    .b(1'b0),
    .c(\PWM6/sub1/c22 ),
    .o({\PWM6/sub1/c23 ,\PWM6/n26 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub1/u23  (
    .a(pnumcnt6[23]),
    .b(1'b0),
    .c(\PWM6/sub1/c23 ),
    .o({open_n52,\PWM6/n26 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub1/u3  (
    .a(pnumcnt6[3]),
    .b(1'b0),
    .c(\PWM6/sub1/c3 ),
    .o({\PWM6/sub1/c4 ,\PWM6/n26 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub1/u4  (
    .a(pnumcnt6[4]),
    .b(1'b0),
    .c(\PWM6/sub1/c4 ),
    .o({\PWM6/sub1/c5 ,\PWM6/n26 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub1/u5  (
    .a(pnumcnt6[5]),
    .b(1'b0),
    .c(\PWM6/sub1/c5 ),
    .o({\PWM6/sub1/c6 ,\PWM6/n26 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub1/u6  (
    .a(pnumcnt6[6]),
    .b(1'b0),
    .c(\PWM6/sub1/c6 ),
    .o({\PWM6/sub1/c7 ,\PWM6/n26 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub1/u7  (
    .a(pnumcnt6[7]),
    .b(1'b0),
    .c(\PWM6/sub1/c7 ),
    .o({\PWM6/sub1/c8 ,\PWM6/n26 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub1/u8  (
    .a(pnumcnt6[8]),
    .b(1'b0),
    .c(\PWM6/sub1/c8 ),
    .o({\PWM6/sub1/c9 ,\PWM6/n26 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM6/sub1/u9  (
    .a(pnumcnt6[9]),
    .b(1'b0),
    .c(\PWM6/sub1/c9 ),
    .o({\PWM6/sub1/c10 ,\PWM6/n26 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \PWM6/sub1/ucin  (
    .a(1'b0),
    .o({\PWM6/sub1/c0 ,open_n55}));
  reg_ar_as_w1 \PWM7/State_reg  (
    .clk(clk100m),
    .d(\PWM7/n10 ),
    .en(1'b1),
    .reset(~rstn),
    .set(1'b0),
    .q(pwm_state_read[7]));  // src/OnePWM.v(26)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[0]  (
    .i(\PWM7/RemaTxNum[0]_keep ),
    .o(pnumcnt7[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[10]  (
    .i(\PWM7/RemaTxNum[10]_keep ),
    .o(pnumcnt7[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[11]  (
    .i(\PWM7/RemaTxNum[11]_keep ),
    .o(pnumcnt7[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[12]  (
    .i(\PWM7/RemaTxNum[12]_keep ),
    .o(pnumcnt7[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[13]  (
    .i(\PWM7/RemaTxNum[13]_keep ),
    .o(pnumcnt7[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[14]  (
    .i(\PWM7/RemaTxNum[14]_keep ),
    .o(pnumcnt7[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[15]  (
    .i(\PWM7/RemaTxNum[15]_keep ),
    .o(pnumcnt7[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[16]  (
    .i(\PWM7/RemaTxNum[16]_keep ),
    .o(pnumcnt7[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[17]  (
    .i(\PWM7/RemaTxNum[17]_keep ),
    .o(pnumcnt7[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[18]  (
    .i(\PWM7/RemaTxNum[18]_keep ),
    .o(pnumcnt7[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[19]  (
    .i(\PWM7/RemaTxNum[19]_keep ),
    .o(pnumcnt7[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[1]  (
    .i(\PWM7/RemaTxNum[1]_keep ),
    .o(pnumcnt7[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[20]  (
    .i(\PWM7/RemaTxNum[20]_keep ),
    .o(pnumcnt7[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[21]  (
    .i(\PWM7/RemaTxNum[21]_keep ),
    .o(pnumcnt7[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[22]  (
    .i(\PWM7/RemaTxNum[22]_keep ),
    .o(pnumcnt7[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[23]  (
    .i(\PWM7/RemaTxNum[23]_keep ),
    .o(pnumcnt7[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[2]  (
    .i(\PWM7/RemaTxNum[2]_keep ),
    .o(pnumcnt7[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[3]  (
    .i(\PWM7/RemaTxNum[3]_keep ),
    .o(pnumcnt7[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[4]  (
    .i(\PWM7/RemaTxNum[4]_keep ),
    .o(pnumcnt7[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[5]  (
    .i(\PWM7/RemaTxNum[5]_keep ),
    .o(pnumcnt7[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[6]  (
    .i(\PWM7/RemaTxNum[6]_keep ),
    .o(pnumcnt7[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[7]  (
    .i(\PWM7/RemaTxNum[7]_keep ),
    .o(pnumcnt7[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[8]  (
    .i(\PWM7/RemaTxNum[8]_keep ),
    .o(pnumcnt7[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[9]  (
    .i(\PWM7/RemaTxNum[9]_keep ),
    .o(pnumcnt7[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_dir  (
    .i(\PWM7/dir_keep ),
    .o(dir_pad[7]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[0]  (
    .i(\PWM7/pnumr[0]_keep ),
    .o(\PWM7/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[10]  (
    .i(\PWM7/pnumr[10]_keep ),
    .o(\PWM7/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[11]  (
    .i(\PWM7/pnumr[11]_keep ),
    .o(\PWM7/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[12]  (
    .i(\PWM7/pnumr[12]_keep ),
    .o(\PWM7/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[13]  (
    .i(\PWM7/pnumr[13]_keep ),
    .o(\PWM7/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[14]  (
    .i(\PWM7/pnumr[14]_keep ),
    .o(\PWM7/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[15]  (
    .i(\PWM7/pnumr[15]_keep ),
    .o(\PWM7/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[16]  (
    .i(\PWM7/pnumr[16]_keep ),
    .o(\PWM7/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[17]  (
    .i(\PWM7/pnumr[17]_keep ),
    .o(\PWM7/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[18]  (
    .i(\PWM7/pnumr[18]_keep ),
    .o(\PWM7/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[19]  (
    .i(\PWM7/pnumr[19]_keep ),
    .o(\PWM7/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[1]  (
    .i(\PWM7/pnumr[1]_keep ),
    .o(\PWM7/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[20]  (
    .i(\PWM7/pnumr[20]_keep ),
    .o(\PWM7/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[21]  (
    .i(\PWM7/pnumr[21]_keep ),
    .o(\PWM7/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[22]  (
    .i(\PWM7/pnumr[22]_keep ),
    .o(\PWM7/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[23]  (
    .i(\PWM7/pnumr[23]_keep ),
    .o(\PWM7/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[24]  (
    .i(\PWM7/pnumr[24]_keep ),
    .o(\PWM7/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[25]  (
    .i(\PWM7/pnumr[25]_keep ),
    .o(\PWM7/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[26]  (
    .i(\PWM7/pnumr[26]_keep ),
    .o(\PWM7/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[27]  (
    .i(\PWM7/pnumr[27]_keep ),
    .o(\PWM7/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[28]  (
    .i(\PWM7/pnumr[28]_keep ),
    .o(\PWM7/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[29]  (
    .i(\PWM7/pnumr[29]_keep ),
    .o(\PWM7/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[2]  (
    .i(\PWM7/pnumr[2]_keep ),
    .o(\PWM7/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[30]  (
    .i(\PWM7/pnumr[30]_keep ),
    .o(\PWM7/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[31]  (
    .i(\PWM7/pnumr[31]_keep ),
    .o(\PWM7/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[3]  (
    .i(\PWM7/pnumr[3]_keep ),
    .o(\PWM7/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[4]  (
    .i(\PWM7/pnumr[4]_keep ),
    .o(\PWM7/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[5]  (
    .i(\PWM7/pnumr[5]_keep ),
    .o(\PWM7/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[6]  (
    .i(\PWM7/pnumr[6]_keep ),
    .o(\PWM7/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[7]  (
    .i(\PWM7/pnumr[7]_keep ),
    .o(\PWM7/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[8]  (
    .i(\PWM7/pnumr[8]_keep ),
    .o(\PWM7/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[9]  (
    .i(\PWM7/pnumr[9]_keep ),
    .o(\PWM7/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pwm  (
    .i(\PWM7/pwm_keep ),
    .o(pwm_pad[7]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_stopreq  (
    .i(\PWM7/stopreq_keep ),
    .o(\PWM7/stopreq ));  // src/OnePWM.v(14)
  reg_ar_as_w1 \PWM7/dir_reg  (
    .clk(clk100m),
    .d(\PWM7/n32 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/dir_keep ));  // src/OnePWM.v(58)
  reg_sr_as_w1 \PWM7/pwm_reg  (
    .clk(clk100m),
    .d(\pwm[7]_d ),
    .en(1'b1),
    .reset(~\PWM7/u14_sel_is_1_o ),
    .set(1'b0),
    .q(\PWM7/pwm_keep ));  // src/OnePWM.v(45)
  reg_sr_as_w1 \PWM7/reg0_b0  (
    .clk(clk100m),
    .d(\PWM7/n13 [0]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [0]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b1  (
    .clk(clk100m),
    .d(\PWM7/n13 [1]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [1]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b10  (
    .clk(clk100m),
    .d(\PWM7/n13 [10]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [10]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b11  (
    .clk(clk100m),
    .d(\PWM7/n13 [11]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [11]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b12  (
    .clk(clk100m),
    .d(\PWM7/n13 [12]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [12]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b13  (
    .clk(clk100m),
    .d(\PWM7/n13 [13]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [13]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b14  (
    .clk(clk100m),
    .d(\PWM7/n13 [14]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [14]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b15  (
    .clk(clk100m),
    .d(\PWM7/n13 [15]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [15]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b16  (
    .clk(clk100m),
    .d(\PWM7/n13 [16]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [16]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b17  (
    .clk(clk100m),
    .d(\PWM7/n13 [17]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [17]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b18  (
    .clk(clk100m),
    .d(\PWM7/n13 [18]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [18]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b19  (
    .clk(clk100m),
    .d(\PWM7/n13 [19]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [19]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b2  (
    .clk(clk100m),
    .d(\PWM7/n13 [2]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [2]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b20  (
    .clk(clk100m),
    .d(\PWM7/n13 [20]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [20]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b21  (
    .clk(clk100m),
    .d(\PWM7/n13 [21]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [21]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b22  (
    .clk(clk100m),
    .d(\PWM7/n13 [22]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [22]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b23  (
    .clk(clk100m),
    .d(\PWM7/n13 [23]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [23]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b24  (
    .clk(clk100m),
    .d(\PWM7/n13 [24]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [24]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b25  (
    .clk(clk100m),
    .d(\PWM7/n13 [25]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [25]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b26  (
    .clk(clk100m),
    .d(\PWM7/n13 [26]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [26]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b3  (
    .clk(clk100m),
    .d(\PWM7/n13 [3]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [3]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b4  (
    .clk(clk100m),
    .d(\PWM7/n13 [4]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [4]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b5  (
    .clk(clk100m),
    .d(\PWM7/n13 [5]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [5]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b6  (
    .clk(clk100m),
    .d(\PWM7/n13 [6]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [6]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b7  (
    .clk(clk100m),
    .d(\PWM7/n13 [7]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [7]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b8  (
    .clk(clk100m),
    .d(\PWM7/n13 [8]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [8]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b9  (
    .clk(clk100m),
    .d(\PWM7/n13 [9]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b0  (
    .clk(clk100m),
    .d(freq7[0]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [0]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b1  (
    .clk(clk100m),
    .d(freq7[1]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [1]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b10  (
    .clk(clk100m),
    .d(freq7[10]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [10]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b11  (
    .clk(clk100m),
    .d(freq7[11]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [11]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b12  (
    .clk(clk100m),
    .d(freq7[12]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [12]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b13  (
    .clk(clk100m),
    .d(freq7[13]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [13]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b14  (
    .clk(clk100m),
    .d(freq7[14]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [14]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b15  (
    .clk(clk100m),
    .d(freq7[15]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [15]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b16  (
    .clk(clk100m),
    .d(freq7[16]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [16]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b17  (
    .clk(clk100m),
    .d(freq7[17]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [17]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b18  (
    .clk(clk100m),
    .d(freq7[18]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [18]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b19  (
    .clk(clk100m),
    .d(freq7[19]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [19]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b2  (
    .clk(clk100m),
    .d(freq7[2]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [2]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b20  (
    .clk(clk100m),
    .d(freq7[20]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [20]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b21  (
    .clk(clk100m),
    .d(freq7[21]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [21]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b22  (
    .clk(clk100m),
    .d(freq7[22]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [22]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b23  (
    .clk(clk100m),
    .d(freq7[23]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [23]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b24  (
    .clk(clk100m),
    .d(freq7[24]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [24]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b25  (
    .clk(clk100m),
    .d(freq7[25]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [25]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b26  (
    .clk(clk100m),
    .d(freq7[26]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [26]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b3  (
    .clk(clk100m),
    .d(freq7[3]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [3]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b4  (
    .clk(clk100m),
    .d(freq7[4]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [4]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b5  (
    .clk(clk100m),
    .d(freq7[5]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [5]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b6  (
    .clk(clk100m),
    .d(freq7[6]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [6]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b7  (
    .clk(clk100m),
    .d(freq7[7]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [7]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b8  (
    .clk(clk100m),
    .d(freq7[8]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [8]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b9  (
    .clk(clk100m),
    .d(freq7[9]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg2_b0  (
    .clk(clk100m),
    .d(\PWM7/n23 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[0]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b1  (
    .clk(clk100m),
    .d(\PWM7/n23 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[1]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b10  (
    .clk(clk100m),
    .d(\PWM7/n23 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[10]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b11  (
    .clk(clk100m),
    .d(\PWM7/n23 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[11]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b12  (
    .clk(clk100m),
    .d(\PWM7/n23 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[12]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b13  (
    .clk(clk100m),
    .d(\PWM7/n23 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[13]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b14  (
    .clk(clk100m),
    .d(\PWM7/n23 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[14]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b15  (
    .clk(clk100m),
    .d(\PWM7/n23 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[15]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b16  (
    .clk(clk100m),
    .d(\PWM7/n23 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[16]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b17  (
    .clk(clk100m),
    .d(\PWM7/n23 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[17]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b18  (
    .clk(clk100m),
    .d(\PWM7/n23 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[18]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b19  (
    .clk(clk100m),
    .d(\PWM7/n23 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[19]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b2  (
    .clk(clk100m),
    .d(\PWM7/n23 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[2]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b20  (
    .clk(clk100m),
    .d(\PWM7/n23 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[20]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b21  (
    .clk(clk100m),
    .d(\PWM7/n23 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[21]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b22  (
    .clk(clk100m),
    .d(\PWM7/n23 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[22]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b23  (
    .clk(clk100m),
    .d(\PWM7/n23 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[23]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b24  (
    .clk(clk100m),
    .d(\PWM7/n23 [24]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[24]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b25  (
    .clk(clk100m),
    .d(\PWM7/n23 [25]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[25]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b26  (
    .clk(clk100m),
    .d(\PWM7/n23 [26]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[26]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b27  (
    .clk(clk100m),
    .d(\PWM7/n23 [27]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[27]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b28  (
    .clk(clk100m),
    .d(\PWM7/n23 [28]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[28]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b29  (
    .clk(clk100m),
    .d(\PWM7/n23 [29]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[29]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b3  (
    .clk(clk100m),
    .d(\PWM7/n23 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[3]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b30  (
    .clk(clk100m),
    .d(\PWM7/n23 [30]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[30]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b31  (
    .clk(clk100m),
    .d(\PWM7/n23 [31]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[31]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b4  (
    .clk(clk100m),
    .d(\PWM7/n23 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[4]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b5  (
    .clk(clk100m),
    .d(\PWM7/n23 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[5]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b6  (
    .clk(clk100m),
    .d(\PWM7/n23 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[6]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b7  (
    .clk(clk100m),
    .d(\PWM7/n23 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[7]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b8  (
    .clk(clk100m),
    .d(\PWM7/n23 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[8]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b9  (
    .clk(clk100m),
    .d(\PWM7/n23 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[9]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg3_b0  (
    .clk(clk100m),
    .d(\PWM7/n31 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[0]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b1  (
    .clk(clk100m),
    .d(\PWM7/n31 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[1]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b10  (
    .clk(clk100m),
    .d(\PWM7/n31 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[10]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b11  (
    .clk(clk100m),
    .d(\PWM7/n31 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[11]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b12  (
    .clk(clk100m),
    .d(\PWM7/n31 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[12]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b13  (
    .clk(clk100m),
    .d(\PWM7/n31 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[13]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b14  (
    .clk(clk100m),
    .d(\PWM7/n31 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[14]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b15  (
    .clk(clk100m),
    .d(\PWM7/n31 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[15]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b16  (
    .clk(clk100m),
    .d(\PWM7/n31 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[16]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b17  (
    .clk(clk100m),
    .d(\PWM7/n31 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[17]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b18  (
    .clk(clk100m),
    .d(\PWM7/n31 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[18]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b19  (
    .clk(clk100m),
    .d(\PWM7/n31 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[19]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b2  (
    .clk(clk100m),
    .d(\PWM7/n31 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[2]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b20  (
    .clk(clk100m),
    .d(\PWM7/n31 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[20]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b21  (
    .clk(clk100m),
    .d(\PWM7/n31 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[21]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b22  (
    .clk(clk100m),
    .d(\PWM7/n31 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[22]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b23  (
    .clk(clk100m),
    .d(\PWM7/n31 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[23]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b3  (
    .clk(clk100m),
    .d(\PWM7/n31 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[3]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b4  (
    .clk(clk100m),
    .d(\PWM7/n31 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[4]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b5  (
    .clk(clk100m),
    .d(\PWM7/n31 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[5]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b6  (
    .clk(clk100m),
    .d(\PWM7/n31 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[6]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b7  (
    .clk(clk100m),
    .d(\PWM7/n31 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[7]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b8  (
    .clk(clk100m),
    .d(\PWM7/n31 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[8]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b9  (
    .clk(clk100m),
    .d(\PWM7/n31 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[9]_keep ));  // src/OnePWM.v(58)
  reg_ar_ss_w1 \PWM7/stopreq_reg  (
    .clk(clk100m),
    .d(\PWM7/n1 ),
    .en(1'b1),
    .reset(1'b0),
    .set(pwm_start_stop[7]),
    .q(\PWM7/stopreq_keep ));  // src/OnePWM.v(15)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub0/u0  (
    .a(\PWM7/FreCnt [0]),
    .b(1'b1),
    .c(\PWM7/sub0/c0 ),
    .o({\PWM7/sub0/c1 ,\PWM7/n12 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub0/u1  (
    .a(\PWM7/FreCnt [1]),
    .b(1'b0),
    .c(\PWM7/sub0/c1 ),
    .o({\PWM7/sub0/c2 ,\PWM7/n12 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub0/u10  (
    .a(\PWM7/FreCnt [10]),
    .b(1'b0),
    .c(\PWM7/sub0/c10 ),
    .o({\PWM7/sub0/c11 ,\PWM7/n12 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub0/u11  (
    .a(\PWM7/FreCnt [11]),
    .b(1'b0),
    .c(\PWM7/sub0/c11 ),
    .o({\PWM7/sub0/c12 ,\PWM7/n12 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub0/u12  (
    .a(\PWM7/FreCnt [12]),
    .b(1'b0),
    .c(\PWM7/sub0/c12 ),
    .o({\PWM7/sub0/c13 ,\PWM7/n12 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub0/u13  (
    .a(\PWM7/FreCnt [13]),
    .b(1'b0),
    .c(\PWM7/sub0/c13 ),
    .o({\PWM7/sub0/c14 ,\PWM7/n12 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub0/u14  (
    .a(\PWM7/FreCnt [14]),
    .b(1'b0),
    .c(\PWM7/sub0/c14 ),
    .o({\PWM7/sub0/c15 ,\PWM7/n12 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub0/u15  (
    .a(\PWM7/FreCnt [15]),
    .b(1'b0),
    .c(\PWM7/sub0/c15 ),
    .o({\PWM7/sub0/c16 ,\PWM7/n12 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub0/u16  (
    .a(\PWM7/FreCnt [16]),
    .b(1'b0),
    .c(\PWM7/sub0/c16 ),
    .o({\PWM7/sub0/c17 ,\PWM7/n12 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub0/u17  (
    .a(\PWM7/FreCnt [17]),
    .b(1'b0),
    .c(\PWM7/sub0/c17 ),
    .o({\PWM7/sub0/c18 ,\PWM7/n12 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub0/u18  (
    .a(\PWM7/FreCnt [18]),
    .b(1'b0),
    .c(\PWM7/sub0/c18 ),
    .o({\PWM7/sub0/c19 ,\PWM7/n12 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub0/u19  (
    .a(\PWM7/FreCnt [19]),
    .b(1'b0),
    .c(\PWM7/sub0/c19 ),
    .o({\PWM7/sub0/c20 ,\PWM7/n12 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub0/u2  (
    .a(\PWM7/FreCnt [2]),
    .b(1'b0),
    .c(\PWM7/sub0/c2 ),
    .o({\PWM7/sub0/c3 ,\PWM7/n12 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub0/u20  (
    .a(\PWM7/FreCnt [20]),
    .b(1'b0),
    .c(\PWM7/sub0/c20 ),
    .o({\PWM7/sub0/c21 ,\PWM7/n12 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub0/u21  (
    .a(\PWM7/FreCnt [21]),
    .b(1'b0),
    .c(\PWM7/sub0/c21 ),
    .o({\PWM7/sub0/c22 ,\PWM7/n12 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub0/u22  (
    .a(\PWM7/FreCnt [22]),
    .b(1'b0),
    .c(\PWM7/sub0/c22 ),
    .o({\PWM7/sub0/c23 ,\PWM7/n12 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub0/u23  (
    .a(\PWM7/FreCnt [23]),
    .b(1'b0),
    .c(\PWM7/sub0/c23 ),
    .o({\PWM7/sub0/c24 ,\PWM7/n12 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub0/u24  (
    .a(\PWM7/FreCnt [24]),
    .b(1'b0),
    .c(\PWM7/sub0/c24 ),
    .o({\PWM7/sub0/c25 ,\PWM7/n12 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub0/u25  (
    .a(\PWM7/FreCnt [25]),
    .b(1'b0),
    .c(\PWM7/sub0/c25 ),
    .o({\PWM7/sub0/c26 ,\PWM7/n12 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub0/u26  (
    .a(\PWM7/FreCnt [26]),
    .b(1'b0),
    .c(\PWM7/sub0/c26 ),
    .o({open_n56,\PWM7/n12 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub0/u3  (
    .a(\PWM7/FreCnt [3]),
    .b(1'b0),
    .c(\PWM7/sub0/c3 ),
    .o({\PWM7/sub0/c4 ,\PWM7/n12 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub0/u4  (
    .a(\PWM7/FreCnt [4]),
    .b(1'b0),
    .c(\PWM7/sub0/c4 ),
    .o({\PWM7/sub0/c5 ,\PWM7/n12 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub0/u5  (
    .a(\PWM7/FreCnt [5]),
    .b(1'b0),
    .c(\PWM7/sub0/c5 ),
    .o({\PWM7/sub0/c6 ,\PWM7/n12 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub0/u6  (
    .a(\PWM7/FreCnt [6]),
    .b(1'b0),
    .c(\PWM7/sub0/c6 ),
    .o({\PWM7/sub0/c7 ,\PWM7/n12 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub0/u7  (
    .a(\PWM7/FreCnt [7]),
    .b(1'b0),
    .c(\PWM7/sub0/c7 ),
    .o({\PWM7/sub0/c8 ,\PWM7/n12 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub0/u8  (
    .a(\PWM7/FreCnt [8]),
    .b(1'b0),
    .c(\PWM7/sub0/c8 ),
    .o({\PWM7/sub0/c9 ,\PWM7/n12 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub0/u9  (
    .a(\PWM7/FreCnt [9]),
    .b(1'b0),
    .c(\PWM7/sub0/c9 ),
    .o({\PWM7/sub0/c10 ,\PWM7/n12 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \PWM7/sub0/ucin  (
    .a(1'b0),
    .o({\PWM7/sub0/c0 ,open_n59}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub1/u0  (
    .a(pnumcnt7[0]),
    .b(1'b1),
    .c(\PWM7/sub1/c0 ),
    .o({\PWM7/sub1/c1 ,\PWM7/n26 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub1/u1  (
    .a(pnumcnt7[1]),
    .b(1'b0),
    .c(\PWM7/sub1/c1 ),
    .o({\PWM7/sub1/c2 ,\PWM7/n26 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub1/u10  (
    .a(pnumcnt7[10]),
    .b(1'b0),
    .c(\PWM7/sub1/c10 ),
    .o({\PWM7/sub1/c11 ,\PWM7/n26 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub1/u11  (
    .a(pnumcnt7[11]),
    .b(1'b0),
    .c(\PWM7/sub1/c11 ),
    .o({\PWM7/sub1/c12 ,\PWM7/n26 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub1/u12  (
    .a(pnumcnt7[12]),
    .b(1'b0),
    .c(\PWM7/sub1/c12 ),
    .o({\PWM7/sub1/c13 ,\PWM7/n26 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub1/u13  (
    .a(pnumcnt7[13]),
    .b(1'b0),
    .c(\PWM7/sub1/c13 ),
    .o({\PWM7/sub1/c14 ,\PWM7/n26 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub1/u14  (
    .a(pnumcnt7[14]),
    .b(1'b0),
    .c(\PWM7/sub1/c14 ),
    .o({\PWM7/sub1/c15 ,\PWM7/n26 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub1/u15  (
    .a(pnumcnt7[15]),
    .b(1'b0),
    .c(\PWM7/sub1/c15 ),
    .o({\PWM7/sub1/c16 ,\PWM7/n26 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub1/u16  (
    .a(pnumcnt7[16]),
    .b(1'b0),
    .c(\PWM7/sub1/c16 ),
    .o({\PWM7/sub1/c17 ,\PWM7/n26 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub1/u17  (
    .a(pnumcnt7[17]),
    .b(1'b0),
    .c(\PWM7/sub1/c17 ),
    .o({\PWM7/sub1/c18 ,\PWM7/n26 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub1/u18  (
    .a(pnumcnt7[18]),
    .b(1'b0),
    .c(\PWM7/sub1/c18 ),
    .o({\PWM7/sub1/c19 ,\PWM7/n26 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub1/u19  (
    .a(pnumcnt7[19]),
    .b(1'b0),
    .c(\PWM7/sub1/c19 ),
    .o({\PWM7/sub1/c20 ,\PWM7/n26 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub1/u2  (
    .a(pnumcnt7[2]),
    .b(1'b0),
    .c(\PWM7/sub1/c2 ),
    .o({\PWM7/sub1/c3 ,\PWM7/n26 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub1/u20  (
    .a(pnumcnt7[20]),
    .b(1'b0),
    .c(\PWM7/sub1/c20 ),
    .o({\PWM7/sub1/c21 ,\PWM7/n26 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub1/u21  (
    .a(pnumcnt7[21]),
    .b(1'b0),
    .c(\PWM7/sub1/c21 ),
    .o({\PWM7/sub1/c22 ,\PWM7/n26 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub1/u22  (
    .a(pnumcnt7[22]),
    .b(1'b0),
    .c(\PWM7/sub1/c22 ),
    .o({\PWM7/sub1/c23 ,\PWM7/n26 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub1/u23  (
    .a(pnumcnt7[23]),
    .b(1'b0),
    .c(\PWM7/sub1/c23 ),
    .o({open_n60,\PWM7/n26 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub1/u3  (
    .a(pnumcnt7[3]),
    .b(1'b0),
    .c(\PWM7/sub1/c3 ),
    .o({\PWM7/sub1/c4 ,\PWM7/n26 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub1/u4  (
    .a(pnumcnt7[4]),
    .b(1'b0),
    .c(\PWM7/sub1/c4 ),
    .o({\PWM7/sub1/c5 ,\PWM7/n26 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub1/u5  (
    .a(pnumcnt7[5]),
    .b(1'b0),
    .c(\PWM7/sub1/c5 ),
    .o({\PWM7/sub1/c6 ,\PWM7/n26 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub1/u6  (
    .a(pnumcnt7[6]),
    .b(1'b0),
    .c(\PWM7/sub1/c6 ),
    .o({\PWM7/sub1/c7 ,\PWM7/n26 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub1/u7  (
    .a(pnumcnt7[7]),
    .b(1'b0),
    .c(\PWM7/sub1/c7 ),
    .o({\PWM7/sub1/c8 ,\PWM7/n26 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub1/u8  (
    .a(pnumcnt7[8]),
    .b(1'b0),
    .c(\PWM7/sub1/c8 ),
    .o({\PWM7/sub1/c9 ,\PWM7/n26 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM7/sub1/u9  (
    .a(pnumcnt7[9]),
    .b(1'b0),
    .c(\PWM7/sub1/c9 ),
    .o({\PWM7/sub1/c10 ,\PWM7/n26 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \PWM7/sub1/ucin  (
    .a(1'b0),
    .o({\PWM7/sub1/c0 ,open_n63}));
  reg_ar_as_w1 \PWM8/State_reg  (
    .clk(clk100m),
    .d(\PWM8/n10 ),
    .en(1'b1),
    .reset(~rstn),
    .set(1'b0),
    .q(pwm_state_read[8]));  // src/OnePWM.v(26)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[0]  (
    .i(\PWM8/RemaTxNum[0]_keep ),
    .o(pnumcnt8[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[10]  (
    .i(\PWM8/RemaTxNum[10]_keep ),
    .o(pnumcnt8[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[11]  (
    .i(\PWM8/RemaTxNum[11]_keep ),
    .o(pnumcnt8[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[12]  (
    .i(\PWM8/RemaTxNum[12]_keep ),
    .o(pnumcnt8[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[13]  (
    .i(\PWM8/RemaTxNum[13]_keep ),
    .o(pnumcnt8[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[14]  (
    .i(\PWM8/RemaTxNum[14]_keep ),
    .o(pnumcnt8[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[15]  (
    .i(\PWM8/RemaTxNum[15]_keep ),
    .o(pnumcnt8[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[16]  (
    .i(\PWM8/RemaTxNum[16]_keep ),
    .o(pnumcnt8[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[17]  (
    .i(\PWM8/RemaTxNum[17]_keep ),
    .o(pnumcnt8[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[18]  (
    .i(\PWM8/RemaTxNum[18]_keep ),
    .o(pnumcnt8[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[19]  (
    .i(\PWM8/RemaTxNum[19]_keep ),
    .o(pnumcnt8[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[1]  (
    .i(\PWM8/RemaTxNum[1]_keep ),
    .o(pnumcnt8[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[20]  (
    .i(\PWM8/RemaTxNum[20]_keep ),
    .o(pnumcnt8[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[21]  (
    .i(\PWM8/RemaTxNum[21]_keep ),
    .o(pnumcnt8[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[22]  (
    .i(\PWM8/RemaTxNum[22]_keep ),
    .o(pnumcnt8[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[23]  (
    .i(\PWM8/RemaTxNum[23]_keep ),
    .o(pnumcnt8[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[2]  (
    .i(\PWM8/RemaTxNum[2]_keep ),
    .o(pnumcnt8[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[3]  (
    .i(\PWM8/RemaTxNum[3]_keep ),
    .o(pnumcnt8[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[4]  (
    .i(\PWM8/RemaTxNum[4]_keep ),
    .o(pnumcnt8[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[5]  (
    .i(\PWM8/RemaTxNum[5]_keep ),
    .o(pnumcnt8[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[6]  (
    .i(\PWM8/RemaTxNum[6]_keep ),
    .o(pnumcnt8[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[7]  (
    .i(\PWM8/RemaTxNum[7]_keep ),
    .o(pnumcnt8[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[8]  (
    .i(\PWM8/RemaTxNum[8]_keep ),
    .o(pnumcnt8[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[9]  (
    .i(\PWM8/RemaTxNum[9]_keep ),
    .o(pnumcnt8[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_dir  (
    .i(\PWM8/dir_keep ),
    .o(dir_pad[8]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[0]  (
    .i(\PWM8/pnumr[0]_keep ),
    .o(\PWM8/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[10]  (
    .i(\PWM8/pnumr[10]_keep ),
    .o(\PWM8/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[11]  (
    .i(\PWM8/pnumr[11]_keep ),
    .o(\PWM8/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[12]  (
    .i(\PWM8/pnumr[12]_keep ),
    .o(\PWM8/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[13]  (
    .i(\PWM8/pnumr[13]_keep ),
    .o(\PWM8/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[14]  (
    .i(\PWM8/pnumr[14]_keep ),
    .o(\PWM8/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[15]  (
    .i(\PWM8/pnumr[15]_keep ),
    .o(\PWM8/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[16]  (
    .i(\PWM8/pnumr[16]_keep ),
    .o(\PWM8/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[17]  (
    .i(\PWM8/pnumr[17]_keep ),
    .o(\PWM8/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[18]  (
    .i(\PWM8/pnumr[18]_keep ),
    .o(\PWM8/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[19]  (
    .i(\PWM8/pnumr[19]_keep ),
    .o(\PWM8/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[1]  (
    .i(\PWM8/pnumr[1]_keep ),
    .o(\PWM8/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[20]  (
    .i(\PWM8/pnumr[20]_keep ),
    .o(\PWM8/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[21]  (
    .i(\PWM8/pnumr[21]_keep ),
    .o(\PWM8/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[22]  (
    .i(\PWM8/pnumr[22]_keep ),
    .o(\PWM8/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[23]  (
    .i(\PWM8/pnumr[23]_keep ),
    .o(\PWM8/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[24]  (
    .i(\PWM8/pnumr[24]_keep ),
    .o(\PWM8/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[25]  (
    .i(\PWM8/pnumr[25]_keep ),
    .o(\PWM8/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[26]  (
    .i(\PWM8/pnumr[26]_keep ),
    .o(\PWM8/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[27]  (
    .i(\PWM8/pnumr[27]_keep ),
    .o(\PWM8/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[28]  (
    .i(\PWM8/pnumr[28]_keep ),
    .o(\PWM8/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[29]  (
    .i(\PWM8/pnumr[29]_keep ),
    .o(\PWM8/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[2]  (
    .i(\PWM8/pnumr[2]_keep ),
    .o(\PWM8/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[30]  (
    .i(\PWM8/pnumr[30]_keep ),
    .o(\PWM8/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[31]  (
    .i(\PWM8/pnumr[31]_keep ),
    .o(\PWM8/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[3]  (
    .i(\PWM8/pnumr[3]_keep ),
    .o(\PWM8/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[4]  (
    .i(\PWM8/pnumr[4]_keep ),
    .o(\PWM8/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[5]  (
    .i(\PWM8/pnumr[5]_keep ),
    .o(\PWM8/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[6]  (
    .i(\PWM8/pnumr[6]_keep ),
    .o(\PWM8/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[7]  (
    .i(\PWM8/pnumr[7]_keep ),
    .o(\PWM8/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[8]  (
    .i(\PWM8/pnumr[8]_keep ),
    .o(\PWM8/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[9]  (
    .i(\PWM8/pnumr[9]_keep ),
    .o(\PWM8/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pwm  (
    .i(\PWM8/pwm_keep ),
    .o(pwm_pad[8]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_stopreq  (
    .i(\PWM8/stopreq_keep ),
    .o(\PWM8/stopreq ));  // src/OnePWM.v(14)
  reg_ar_as_w1 \PWM8/dir_reg  (
    .clk(clk100m),
    .d(\PWM8/n32 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/dir_keep ));  // src/OnePWM.v(58)
  reg_sr_as_w1 \PWM8/pwm_reg  (
    .clk(clk100m),
    .d(\pwm[8]_d ),
    .en(1'b1),
    .reset(~\PWM8/u14_sel_is_1_o ),
    .set(1'b0),
    .q(\PWM8/pwm_keep ));  // src/OnePWM.v(45)
  reg_sr_as_w1 \PWM8/reg0_b0  (
    .clk(clk100m),
    .d(\PWM8/n13 [0]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [0]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b1  (
    .clk(clk100m),
    .d(\PWM8/n13 [1]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [1]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b10  (
    .clk(clk100m),
    .d(\PWM8/n13 [10]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [10]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b11  (
    .clk(clk100m),
    .d(\PWM8/n13 [11]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [11]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b12  (
    .clk(clk100m),
    .d(\PWM8/n13 [12]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [12]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b13  (
    .clk(clk100m),
    .d(\PWM8/n13 [13]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [13]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b14  (
    .clk(clk100m),
    .d(\PWM8/n13 [14]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [14]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b15  (
    .clk(clk100m),
    .d(\PWM8/n13 [15]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [15]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b16  (
    .clk(clk100m),
    .d(\PWM8/n13 [16]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [16]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b17  (
    .clk(clk100m),
    .d(\PWM8/n13 [17]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [17]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b18  (
    .clk(clk100m),
    .d(\PWM8/n13 [18]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [18]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b19  (
    .clk(clk100m),
    .d(\PWM8/n13 [19]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [19]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b2  (
    .clk(clk100m),
    .d(\PWM8/n13 [2]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [2]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b20  (
    .clk(clk100m),
    .d(\PWM8/n13 [20]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [20]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b21  (
    .clk(clk100m),
    .d(\PWM8/n13 [21]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [21]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b22  (
    .clk(clk100m),
    .d(\PWM8/n13 [22]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [22]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b23  (
    .clk(clk100m),
    .d(\PWM8/n13 [23]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [23]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b24  (
    .clk(clk100m),
    .d(\PWM8/n13 [24]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [24]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b25  (
    .clk(clk100m),
    .d(\PWM8/n13 [25]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [25]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b26  (
    .clk(clk100m),
    .d(\PWM8/n13 [26]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [26]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b3  (
    .clk(clk100m),
    .d(\PWM8/n13 [3]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [3]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b4  (
    .clk(clk100m),
    .d(\PWM8/n13 [4]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [4]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b5  (
    .clk(clk100m),
    .d(\PWM8/n13 [5]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [5]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b6  (
    .clk(clk100m),
    .d(\PWM8/n13 [6]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [6]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b7  (
    .clk(clk100m),
    .d(\PWM8/n13 [7]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [7]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b8  (
    .clk(clk100m),
    .d(\PWM8/n13 [8]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [8]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b9  (
    .clk(clk100m),
    .d(\PWM8/n13 [9]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b0  (
    .clk(clk100m),
    .d(freq8[0]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [0]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b1  (
    .clk(clk100m),
    .d(freq8[1]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [1]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b10  (
    .clk(clk100m),
    .d(freq8[10]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [10]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b11  (
    .clk(clk100m),
    .d(freq8[11]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [11]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b12  (
    .clk(clk100m),
    .d(freq8[12]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [12]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b13  (
    .clk(clk100m),
    .d(freq8[13]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [13]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b14  (
    .clk(clk100m),
    .d(freq8[14]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [14]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b15  (
    .clk(clk100m),
    .d(freq8[15]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [15]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b16  (
    .clk(clk100m),
    .d(freq8[16]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [16]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b17  (
    .clk(clk100m),
    .d(freq8[17]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [17]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b18  (
    .clk(clk100m),
    .d(freq8[18]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [18]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b19  (
    .clk(clk100m),
    .d(freq8[19]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [19]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b2  (
    .clk(clk100m),
    .d(freq8[2]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [2]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b20  (
    .clk(clk100m),
    .d(freq8[20]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [20]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b21  (
    .clk(clk100m),
    .d(freq8[21]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [21]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b22  (
    .clk(clk100m),
    .d(freq8[22]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [22]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b23  (
    .clk(clk100m),
    .d(freq8[23]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [23]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b24  (
    .clk(clk100m),
    .d(freq8[24]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [24]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b25  (
    .clk(clk100m),
    .d(freq8[25]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [25]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b26  (
    .clk(clk100m),
    .d(freq8[26]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [26]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b3  (
    .clk(clk100m),
    .d(freq8[3]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [3]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b4  (
    .clk(clk100m),
    .d(freq8[4]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [4]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b5  (
    .clk(clk100m),
    .d(freq8[5]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [5]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b6  (
    .clk(clk100m),
    .d(freq8[6]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [6]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b7  (
    .clk(clk100m),
    .d(freq8[7]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [7]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b8  (
    .clk(clk100m),
    .d(freq8[8]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [8]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b9  (
    .clk(clk100m),
    .d(freq8[9]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg2_b0  (
    .clk(clk100m),
    .d(\PWM8/n23 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[0]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b1  (
    .clk(clk100m),
    .d(\PWM8/n23 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[1]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b10  (
    .clk(clk100m),
    .d(\PWM8/n23 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[10]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b11  (
    .clk(clk100m),
    .d(\PWM8/n23 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[11]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b12  (
    .clk(clk100m),
    .d(\PWM8/n23 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[12]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b13  (
    .clk(clk100m),
    .d(\PWM8/n23 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[13]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b14  (
    .clk(clk100m),
    .d(\PWM8/n23 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[14]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b15  (
    .clk(clk100m),
    .d(\PWM8/n23 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[15]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b16  (
    .clk(clk100m),
    .d(\PWM8/n23 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[16]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b17  (
    .clk(clk100m),
    .d(\PWM8/n23 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[17]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b18  (
    .clk(clk100m),
    .d(\PWM8/n23 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[18]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b19  (
    .clk(clk100m),
    .d(\PWM8/n23 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[19]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b2  (
    .clk(clk100m),
    .d(\PWM8/n23 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[2]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b20  (
    .clk(clk100m),
    .d(\PWM8/n23 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[20]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b21  (
    .clk(clk100m),
    .d(\PWM8/n23 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[21]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b22  (
    .clk(clk100m),
    .d(\PWM8/n23 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[22]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b23  (
    .clk(clk100m),
    .d(\PWM8/n23 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[23]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b24  (
    .clk(clk100m),
    .d(\PWM8/n23 [24]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[24]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b25  (
    .clk(clk100m),
    .d(\PWM8/n23 [25]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[25]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b26  (
    .clk(clk100m),
    .d(\PWM8/n23 [26]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[26]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b27  (
    .clk(clk100m),
    .d(\PWM8/n23 [27]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[27]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b28  (
    .clk(clk100m),
    .d(\PWM8/n23 [28]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[28]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b29  (
    .clk(clk100m),
    .d(\PWM8/n23 [29]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[29]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b3  (
    .clk(clk100m),
    .d(\PWM8/n23 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[3]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b30  (
    .clk(clk100m),
    .d(\PWM8/n23 [30]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[30]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b31  (
    .clk(clk100m),
    .d(\PWM8/n23 [31]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[31]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b4  (
    .clk(clk100m),
    .d(\PWM8/n23 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[4]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b5  (
    .clk(clk100m),
    .d(\PWM8/n23 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[5]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b6  (
    .clk(clk100m),
    .d(\PWM8/n23 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[6]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b7  (
    .clk(clk100m),
    .d(\PWM8/n23 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[7]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b8  (
    .clk(clk100m),
    .d(\PWM8/n23 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[8]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b9  (
    .clk(clk100m),
    .d(\PWM8/n23 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[9]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg3_b0  (
    .clk(clk100m),
    .d(\PWM8/n31 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[0]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b1  (
    .clk(clk100m),
    .d(\PWM8/n31 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[1]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b10  (
    .clk(clk100m),
    .d(\PWM8/n31 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[10]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b11  (
    .clk(clk100m),
    .d(\PWM8/n31 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[11]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b12  (
    .clk(clk100m),
    .d(\PWM8/n31 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[12]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b13  (
    .clk(clk100m),
    .d(\PWM8/n31 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[13]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b14  (
    .clk(clk100m),
    .d(\PWM8/n31 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[14]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b15  (
    .clk(clk100m),
    .d(\PWM8/n31 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[15]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b16  (
    .clk(clk100m),
    .d(\PWM8/n31 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[16]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b17  (
    .clk(clk100m),
    .d(\PWM8/n31 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[17]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b18  (
    .clk(clk100m),
    .d(\PWM8/n31 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[18]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b19  (
    .clk(clk100m),
    .d(\PWM8/n31 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[19]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b2  (
    .clk(clk100m),
    .d(\PWM8/n31 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[2]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b20  (
    .clk(clk100m),
    .d(\PWM8/n31 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[20]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b21  (
    .clk(clk100m),
    .d(\PWM8/n31 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[21]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b22  (
    .clk(clk100m),
    .d(\PWM8/n31 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[22]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b23  (
    .clk(clk100m),
    .d(\PWM8/n31 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[23]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b3  (
    .clk(clk100m),
    .d(\PWM8/n31 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[3]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b4  (
    .clk(clk100m),
    .d(\PWM8/n31 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[4]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b5  (
    .clk(clk100m),
    .d(\PWM8/n31 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[5]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b6  (
    .clk(clk100m),
    .d(\PWM8/n31 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[6]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b7  (
    .clk(clk100m),
    .d(\PWM8/n31 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[7]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b8  (
    .clk(clk100m),
    .d(\PWM8/n31 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[8]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b9  (
    .clk(clk100m),
    .d(\PWM8/n31 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[9]_keep ));  // src/OnePWM.v(58)
  reg_ar_ss_w1 \PWM8/stopreq_reg  (
    .clk(clk100m),
    .d(\PWM8/n1 ),
    .en(1'b1),
    .reset(1'b0),
    .set(pwm_start_stop[8]),
    .q(\PWM8/stopreq_keep ));  // src/OnePWM.v(15)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub0/u0  (
    .a(\PWM8/FreCnt [0]),
    .b(1'b1),
    .c(\PWM8/sub0/c0 ),
    .o({\PWM8/sub0/c1 ,\PWM8/n12 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub0/u1  (
    .a(\PWM8/FreCnt [1]),
    .b(1'b0),
    .c(\PWM8/sub0/c1 ),
    .o({\PWM8/sub0/c2 ,\PWM8/n12 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub0/u10  (
    .a(\PWM8/FreCnt [10]),
    .b(1'b0),
    .c(\PWM8/sub0/c10 ),
    .o({\PWM8/sub0/c11 ,\PWM8/n12 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub0/u11  (
    .a(\PWM8/FreCnt [11]),
    .b(1'b0),
    .c(\PWM8/sub0/c11 ),
    .o({\PWM8/sub0/c12 ,\PWM8/n12 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub0/u12  (
    .a(\PWM8/FreCnt [12]),
    .b(1'b0),
    .c(\PWM8/sub0/c12 ),
    .o({\PWM8/sub0/c13 ,\PWM8/n12 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub0/u13  (
    .a(\PWM8/FreCnt [13]),
    .b(1'b0),
    .c(\PWM8/sub0/c13 ),
    .o({\PWM8/sub0/c14 ,\PWM8/n12 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub0/u14  (
    .a(\PWM8/FreCnt [14]),
    .b(1'b0),
    .c(\PWM8/sub0/c14 ),
    .o({\PWM8/sub0/c15 ,\PWM8/n12 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub0/u15  (
    .a(\PWM8/FreCnt [15]),
    .b(1'b0),
    .c(\PWM8/sub0/c15 ),
    .o({\PWM8/sub0/c16 ,\PWM8/n12 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub0/u16  (
    .a(\PWM8/FreCnt [16]),
    .b(1'b0),
    .c(\PWM8/sub0/c16 ),
    .o({\PWM8/sub0/c17 ,\PWM8/n12 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub0/u17  (
    .a(\PWM8/FreCnt [17]),
    .b(1'b0),
    .c(\PWM8/sub0/c17 ),
    .o({\PWM8/sub0/c18 ,\PWM8/n12 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub0/u18  (
    .a(\PWM8/FreCnt [18]),
    .b(1'b0),
    .c(\PWM8/sub0/c18 ),
    .o({\PWM8/sub0/c19 ,\PWM8/n12 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub0/u19  (
    .a(\PWM8/FreCnt [19]),
    .b(1'b0),
    .c(\PWM8/sub0/c19 ),
    .o({\PWM8/sub0/c20 ,\PWM8/n12 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub0/u2  (
    .a(\PWM8/FreCnt [2]),
    .b(1'b0),
    .c(\PWM8/sub0/c2 ),
    .o({\PWM8/sub0/c3 ,\PWM8/n12 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub0/u20  (
    .a(\PWM8/FreCnt [20]),
    .b(1'b0),
    .c(\PWM8/sub0/c20 ),
    .o({\PWM8/sub0/c21 ,\PWM8/n12 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub0/u21  (
    .a(\PWM8/FreCnt [21]),
    .b(1'b0),
    .c(\PWM8/sub0/c21 ),
    .o({\PWM8/sub0/c22 ,\PWM8/n12 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub0/u22  (
    .a(\PWM8/FreCnt [22]),
    .b(1'b0),
    .c(\PWM8/sub0/c22 ),
    .o({\PWM8/sub0/c23 ,\PWM8/n12 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub0/u23  (
    .a(\PWM8/FreCnt [23]),
    .b(1'b0),
    .c(\PWM8/sub0/c23 ),
    .o({\PWM8/sub0/c24 ,\PWM8/n12 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub0/u24  (
    .a(\PWM8/FreCnt [24]),
    .b(1'b0),
    .c(\PWM8/sub0/c24 ),
    .o({\PWM8/sub0/c25 ,\PWM8/n12 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub0/u25  (
    .a(\PWM8/FreCnt [25]),
    .b(1'b0),
    .c(\PWM8/sub0/c25 ),
    .o({\PWM8/sub0/c26 ,\PWM8/n12 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub0/u26  (
    .a(\PWM8/FreCnt [26]),
    .b(1'b0),
    .c(\PWM8/sub0/c26 ),
    .o({open_n64,\PWM8/n12 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub0/u3  (
    .a(\PWM8/FreCnt [3]),
    .b(1'b0),
    .c(\PWM8/sub0/c3 ),
    .o({\PWM8/sub0/c4 ,\PWM8/n12 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub0/u4  (
    .a(\PWM8/FreCnt [4]),
    .b(1'b0),
    .c(\PWM8/sub0/c4 ),
    .o({\PWM8/sub0/c5 ,\PWM8/n12 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub0/u5  (
    .a(\PWM8/FreCnt [5]),
    .b(1'b0),
    .c(\PWM8/sub0/c5 ),
    .o({\PWM8/sub0/c6 ,\PWM8/n12 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub0/u6  (
    .a(\PWM8/FreCnt [6]),
    .b(1'b0),
    .c(\PWM8/sub0/c6 ),
    .o({\PWM8/sub0/c7 ,\PWM8/n12 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub0/u7  (
    .a(\PWM8/FreCnt [7]),
    .b(1'b0),
    .c(\PWM8/sub0/c7 ),
    .o({\PWM8/sub0/c8 ,\PWM8/n12 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub0/u8  (
    .a(\PWM8/FreCnt [8]),
    .b(1'b0),
    .c(\PWM8/sub0/c8 ),
    .o({\PWM8/sub0/c9 ,\PWM8/n12 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub0/u9  (
    .a(\PWM8/FreCnt [9]),
    .b(1'b0),
    .c(\PWM8/sub0/c9 ),
    .o({\PWM8/sub0/c10 ,\PWM8/n12 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \PWM8/sub0/ucin  (
    .a(1'b0),
    .o({\PWM8/sub0/c0 ,open_n67}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub1/u0  (
    .a(pnumcnt8[0]),
    .b(1'b1),
    .c(\PWM8/sub1/c0 ),
    .o({\PWM8/sub1/c1 ,\PWM8/n26 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub1/u1  (
    .a(pnumcnt8[1]),
    .b(1'b0),
    .c(\PWM8/sub1/c1 ),
    .o({\PWM8/sub1/c2 ,\PWM8/n26 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub1/u10  (
    .a(pnumcnt8[10]),
    .b(1'b0),
    .c(\PWM8/sub1/c10 ),
    .o({\PWM8/sub1/c11 ,\PWM8/n26 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub1/u11  (
    .a(pnumcnt8[11]),
    .b(1'b0),
    .c(\PWM8/sub1/c11 ),
    .o({\PWM8/sub1/c12 ,\PWM8/n26 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub1/u12  (
    .a(pnumcnt8[12]),
    .b(1'b0),
    .c(\PWM8/sub1/c12 ),
    .o({\PWM8/sub1/c13 ,\PWM8/n26 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub1/u13  (
    .a(pnumcnt8[13]),
    .b(1'b0),
    .c(\PWM8/sub1/c13 ),
    .o({\PWM8/sub1/c14 ,\PWM8/n26 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub1/u14  (
    .a(pnumcnt8[14]),
    .b(1'b0),
    .c(\PWM8/sub1/c14 ),
    .o({\PWM8/sub1/c15 ,\PWM8/n26 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub1/u15  (
    .a(pnumcnt8[15]),
    .b(1'b0),
    .c(\PWM8/sub1/c15 ),
    .o({\PWM8/sub1/c16 ,\PWM8/n26 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub1/u16  (
    .a(pnumcnt8[16]),
    .b(1'b0),
    .c(\PWM8/sub1/c16 ),
    .o({\PWM8/sub1/c17 ,\PWM8/n26 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub1/u17  (
    .a(pnumcnt8[17]),
    .b(1'b0),
    .c(\PWM8/sub1/c17 ),
    .o({\PWM8/sub1/c18 ,\PWM8/n26 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub1/u18  (
    .a(pnumcnt8[18]),
    .b(1'b0),
    .c(\PWM8/sub1/c18 ),
    .o({\PWM8/sub1/c19 ,\PWM8/n26 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub1/u19  (
    .a(pnumcnt8[19]),
    .b(1'b0),
    .c(\PWM8/sub1/c19 ),
    .o({\PWM8/sub1/c20 ,\PWM8/n26 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub1/u2  (
    .a(pnumcnt8[2]),
    .b(1'b0),
    .c(\PWM8/sub1/c2 ),
    .o({\PWM8/sub1/c3 ,\PWM8/n26 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub1/u20  (
    .a(pnumcnt8[20]),
    .b(1'b0),
    .c(\PWM8/sub1/c20 ),
    .o({\PWM8/sub1/c21 ,\PWM8/n26 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub1/u21  (
    .a(pnumcnt8[21]),
    .b(1'b0),
    .c(\PWM8/sub1/c21 ),
    .o({\PWM8/sub1/c22 ,\PWM8/n26 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub1/u22  (
    .a(pnumcnt8[22]),
    .b(1'b0),
    .c(\PWM8/sub1/c22 ),
    .o({\PWM8/sub1/c23 ,\PWM8/n26 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub1/u23  (
    .a(pnumcnt8[23]),
    .b(1'b0),
    .c(\PWM8/sub1/c23 ),
    .o({open_n68,\PWM8/n26 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub1/u3  (
    .a(pnumcnt8[3]),
    .b(1'b0),
    .c(\PWM8/sub1/c3 ),
    .o({\PWM8/sub1/c4 ,\PWM8/n26 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub1/u4  (
    .a(pnumcnt8[4]),
    .b(1'b0),
    .c(\PWM8/sub1/c4 ),
    .o({\PWM8/sub1/c5 ,\PWM8/n26 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub1/u5  (
    .a(pnumcnt8[5]),
    .b(1'b0),
    .c(\PWM8/sub1/c5 ),
    .o({\PWM8/sub1/c6 ,\PWM8/n26 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub1/u6  (
    .a(pnumcnt8[6]),
    .b(1'b0),
    .c(\PWM8/sub1/c6 ),
    .o({\PWM8/sub1/c7 ,\PWM8/n26 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub1/u7  (
    .a(pnumcnt8[7]),
    .b(1'b0),
    .c(\PWM8/sub1/c7 ),
    .o({\PWM8/sub1/c8 ,\PWM8/n26 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub1/u8  (
    .a(pnumcnt8[8]),
    .b(1'b0),
    .c(\PWM8/sub1/c8 ),
    .o({\PWM8/sub1/c9 ,\PWM8/n26 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM8/sub1/u9  (
    .a(pnumcnt8[9]),
    .b(1'b0),
    .c(\PWM8/sub1/c9 ),
    .o({\PWM8/sub1/c10 ,\PWM8/n26 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \PWM8/sub1/ucin  (
    .a(1'b0),
    .o({\PWM8/sub1/c0 ,open_n71}));
  reg_ar_as_w1 \PWM9/State_reg  (
    .clk(clk100m),
    .d(\PWM9/n10 ),
    .en(1'b1),
    .reset(~rstn),
    .set(1'b0),
    .q(pwm_state_read[9]));  // src/OnePWM.v(26)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[0]  (
    .i(\PWM9/RemaTxNum[0]_keep ),
    .o(pnumcnt9[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[10]  (
    .i(\PWM9/RemaTxNum[10]_keep ),
    .o(pnumcnt9[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[11]  (
    .i(\PWM9/RemaTxNum[11]_keep ),
    .o(pnumcnt9[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[12]  (
    .i(\PWM9/RemaTxNum[12]_keep ),
    .o(pnumcnt9[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[13]  (
    .i(\PWM9/RemaTxNum[13]_keep ),
    .o(pnumcnt9[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[14]  (
    .i(\PWM9/RemaTxNum[14]_keep ),
    .o(pnumcnt9[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[15]  (
    .i(\PWM9/RemaTxNum[15]_keep ),
    .o(pnumcnt9[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[16]  (
    .i(\PWM9/RemaTxNum[16]_keep ),
    .o(pnumcnt9[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[17]  (
    .i(\PWM9/RemaTxNum[17]_keep ),
    .o(pnumcnt9[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[18]  (
    .i(\PWM9/RemaTxNum[18]_keep ),
    .o(pnumcnt9[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[19]  (
    .i(\PWM9/RemaTxNum[19]_keep ),
    .o(pnumcnt9[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[1]  (
    .i(\PWM9/RemaTxNum[1]_keep ),
    .o(pnumcnt9[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[20]  (
    .i(\PWM9/RemaTxNum[20]_keep ),
    .o(pnumcnt9[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[21]  (
    .i(\PWM9/RemaTxNum[21]_keep ),
    .o(pnumcnt9[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[22]  (
    .i(\PWM9/RemaTxNum[22]_keep ),
    .o(pnumcnt9[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[23]  (
    .i(\PWM9/RemaTxNum[23]_keep ),
    .o(pnumcnt9[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[2]  (
    .i(\PWM9/RemaTxNum[2]_keep ),
    .o(pnumcnt9[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[3]  (
    .i(\PWM9/RemaTxNum[3]_keep ),
    .o(pnumcnt9[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[4]  (
    .i(\PWM9/RemaTxNum[4]_keep ),
    .o(pnumcnt9[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[5]  (
    .i(\PWM9/RemaTxNum[5]_keep ),
    .o(pnumcnt9[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[6]  (
    .i(\PWM9/RemaTxNum[6]_keep ),
    .o(pnumcnt9[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[7]  (
    .i(\PWM9/RemaTxNum[7]_keep ),
    .o(pnumcnt9[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[8]  (
    .i(\PWM9/RemaTxNum[8]_keep ),
    .o(pnumcnt9[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[9]  (
    .i(\PWM9/RemaTxNum[9]_keep ),
    .o(pnumcnt9[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_dir  (
    .i(\PWM9/dir_keep ),
    .o(dir_pad[9]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[0]  (
    .i(\PWM9/pnumr[0]_keep ),
    .o(\PWM9/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[10]  (
    .i(\PWM9/pnumr[10]_keep ),
    .o(\PWM9/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[11]  (
    .i(\PWM9/pnumr[11]_keep ),
    .o(\PWM9/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[12]  (
    .i(\PWM9/pnumr[12]_keep ),
    .o(\PWM9/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[13]  (
    .i(\PWM9/pnumr[13]_keep ),
    .o(\PWM9/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[14]  (
    .i(\PWM9/pnumr[14]_keep ),
    .o(\PWM9/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[15]  (
    .i(\PWM9/pnumr[15]_keep ),
    .o(\PWM9/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[16]  (
    .i(\PWM9/pnumr[16]_keep ),
    .o(\PWM9/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[17]  (
    .i(\PWM9/pnumr[17]_keep ),
    .o(\PWM9/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[18]  (
    .i(\PWM9/pnumr[18]_keep ),
    .o(\PWM9/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[19]  (
    .i(\PWM9/pnumr[19]_keep ),
    .o(\PWM9/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[1]  (
    .i(\PWM9/pnumr[1]_keep ),
    .o(\PWM9/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[20]  (
    .i(\PWM9/pnumr[20]_keep ),
    .o(\PWM9/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[21]  (
    .i(\PWM9/pnumr[21]_keep ),
    .o(\PWM9/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[22]  (
    .i(\PWM9/pnumr[22]_keep ),
    .o(\PWM9/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[23]  (
    .i(\PWM9/pnumr[23]_keep ),
    .o(\PWM9/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[24]  (
    .i(\PWM9/pnumr[24]_keep ),
    .o(\PWM9/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[25]  (
    .i(\PWM9/pnumr[25]_keep ),
    .o(\PWM9/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[26]  (
    .i(\PWM9/pnumr[26]_keep ),
    .o(\PWM9/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[27]  (
    .i(\PWM9/pnumr[27]_keep ),
    .o(\PWM9/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[28]  (
    .i(\PWM9/pnumr[28]_keep ),
    .o(\PWM9/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[29]  (
    .i(\PWM9/pnumr[29]_keep ),
    .o(\PWM9/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[2]  (
    .i(\PWM9/pnumr[2]_keep ),
    .o(\PWM9/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[30]  (
    .i(\PWM9/pnumr[30]_keep ),
    .o(\PWM9/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[31]  (
    .i(\PWM9/pnumr[31]_keep ),
    .o(\PWM9/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[3]  (
    .i(\PWM9/pnumr[3]_keep ),
    .o(\PWM9/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[4]  (
    .i(\PWM9/pnumr[4]_keep ),
    .o(\PWM9/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[5]  (
    .i(\PWM9/pnumr[5]_keep ),
    .o(\PWM9/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[6]  (
    .i(\PWM9/pnumr[6]_keep ),
    .o(\PWM9/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[7]  (
    .i(\PWM9/pnumr[7]_keep ),
    .o(\PWM9/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[8]  (
    .i(\PWM9/pnumr[8]_keep ),
    .o(\PWM9/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[9]  (
    .i(\PWM9/pnumr[9]_keep ),
    .o(\PWM9/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pwm  (
    .i(\PWM9/pwm_keep ),
    .o(pwm_pad[9]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_stopreq  (
    .i(\PWM9/stopreq_keep ),
    .o(\PWM9/stopreq ));  // src/OnePWM.v(14)
  reg_ar_as_w1 \PWM9/dir_reg  (
    .clk(clk100m),
    .d(\PWM9/n32 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/dir_keep ));  // src/OnePWM.v(58)
  reg_sr_as_w1 \PWM9/pwm_reg  (
    .clk(clk100m),
    .d(\pwm[9]_d ),
    .en(1'b1),
    .reset(~\PWM9/u14_sel_is_1_o ),
    .set(1'b0),
    .q(\PWM9/pwm_keep ));  // src/OnePWM.v(45)
  reg_sr_as_w1 \PWM9/reg0_b0  (
    .clk(clk100m),
    .d(\PWM9/n13 [0]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [0]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b1  (
    .clk(clk100m),
    .d(\PWM9/n13 [1]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [1]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b10  (
    .clk(clk100m),
    .d(\PWM9/n13 [10]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [10]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b11  (
    .clk(clk100m),
    .d(\PWM9/n13 [11]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [11]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b12  (
    .clk(clk100m),
    .d(\PWM9/n13 [12]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [12]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b13  (
    .clk(clk100m),
    .d(\PWM9/n13 [13]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [13]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b14  (
    .clk(clk100m),
    .d(\PWM9/n13 [14]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [14]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b15  (
    .clk(clk100m),
    .d(\PWM9/n13 [15]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [15]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b16  (
    .clk(clk100m),
    .d(\PWM9/n13 [16]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [16]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b17  (
    .clk(clk100m),
    .d(\PWM9/n13 [17]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [17]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b18  (
    .clk(clk100m),
    .d(\PWM9/n13 [18]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [18]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b19  (
    .clk(clk100m),
    .d(\PWM9/n13 [19]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [19]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b2  (
    .clk(clk100m),
    .d(\PWM9/n13 [2]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [2]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b20  (
    .clk(clk100m),
    .d(\PWM9/n13 [20]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [20]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b21  (
    .clk(clk100m),
    .d(\PWM9/n13 [21]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [21]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b22  (
    .clk(clk100m),
    .d(\PWM9/n13 [22]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [22]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b23  (
    .clk(clk100m),
    .d(\PWM9/n13 [23]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [23]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b24  (
    .clk(clk100m),
    .d(\PWM9/n13 [24]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [24]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b25  (
    .clk(clk100m),
    .d(\PWM9/n13 [25]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [25]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b26  (
    .clk(clk100m),
    .d(\PWM9/n13 [26]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [26]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b3  (
    .clk(clk100m),
    .d(\PWM9/n13 [3]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [3]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b4  (
    .clk(clk100m),
    .d(\PWM9/n13 [4]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [4]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b5  (
    .clk(clk100m),
    .d(\PWM9/n13 [5]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [5]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b6  (
    .clk(clk100m),
    .d(\PWM9/n13 [6]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [6]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b7  (
    .clk(clk100m),
    .d(\PWM9/n13 [7]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [7]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b8  (
    .clk(clk100m),
    .d(\PWM9/n13 [8]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [8]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b9  (
    .clk(clk100m),
    .d(\PWM9/n13 [9]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b0  (
    .clk(clk100m),
    .d(freq9[0]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [0]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b1  (
    .clk(clk100m),
    .d(freq9[1]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [1]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b10  (
    .clk(clk100m),
    .d(freq9[10]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [10]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b11  (
    .clk(clk100m),
    .d(freq9[11]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [11]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b12  (
    .clk(clk100m),
    .d(freq9[12]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [12]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b13  (
    .clk(clk100m),
    .d(freq9[13]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [13]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b14  (
    .clk(clk100m),
    .d(freq9[14]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [14]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b15  (
    .clk(clk100m),
    .d(freq9[15]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [15]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b16  (
    .clk(clk100m),
    .d(freq9[16]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [16]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b17  (
    .clk(clk100m),
    .d(freq9[17]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [17]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b18  (
    .clk(clk100m),
    .d(freq9[18]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [18]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b19  (
    .clk(clk100m),
    .d(freq9[19]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [19]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b2  (
    .clk(clk100m),
    .d(freq9[2]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [2]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b20  (
    .clk(clk100m),
    .d(freq9[20]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [20]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b21  (
    .clk(clk100m),
    .d(freq9[21]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [21]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b22  (
    .clk(clk100m),
    .d(freq9[22]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [22]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b23  (
    .clk(clk100m),
    .d(freq9[23]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [23]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b24  (
    .clk(clk100m),
    .d(freq9[24]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [24]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b25  (
    .clk(clk100m),
    .d(freq9[25]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [25]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b26  (
    .clk(clk100m),
    .d(freq9[26]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [26]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b3  (
    .clk(clk100m),
    .d(freq9[3]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [3]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b4  (
    .clk(clk100m),
    .d(freq9[4]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [4]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b5  (
    .clk(clk100m),
    .d(freq9[5]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [5]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b6  (
    .clk(clk100m),
    .d(freq9[6]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [6]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b7  (
    .clk(clk100m),
    .d(freq9[7]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [7]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b8  (
    .clk(clk100m),
    .d(freq9[8]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [8]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b9  (
    .clk(clk100m),
    .d(freq9[9]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg2_b0  (
    .clk(clk100m),
    .d(\PWM9/n23 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[0]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b1  (
    .clk(clk100m),
    .d(\PWM9/n23 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[1]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b10  (
    .clk(clk100m),
    .d(\PWM9/n23 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[10]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b11  (
    .clk(clk100m),
    .d(\PWM9/n23 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[11]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b12  (
    .clk(clk100m),
    .d(\PWM9/n23 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[12]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b13  (
    .clk(clk100m),
    .d(\PWM9/n23 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[13]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b14  (
    .clk(clk100m),
    .d(\PWM9/n23 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[14]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b15  (
    .clk(clk100m),
    .d(\PWM9/n23 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[15]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b16  (
    .clk(clk100m),
    .d(\PWM9/n23 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[16]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b17  (
    .clk(clk100m),
    .d(\PWM9/n23 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[17]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b18  (
    .clk(clk100m),
    .d(\PWM9/n23 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[18]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b19  (
    .clk(clk100m),
    .d(\PWM9/n23 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[19]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b2  (
    .clk(clk100m),
    .d(\PWM9/n23 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[2]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b20  (
    .clk(clk100m),
    .d(\PWM9/n23 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[20]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b21  (
    .clk(clk100m),
    .d(\PWM9/n23 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[21]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b22  (
    .clk(clk100m),
    .d(\PWM9/n23 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[22]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b23  (
    .clk(clk100m),
    .d(\PWM9/n23 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[23]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b24  (
    .clk(clk100m),
    .d(\PWM9/n23 [24]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[24]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b25  (
    .clk(clk100m),
    .d(\PWM9/n23 [25]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[25]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b26  (
    .clk(clk100m),
    .d(\PWM9/n23 [26]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[26]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b27  (
    .clk(clk100m),
    .d(\PWM9/n23 [27]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[27]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b28  (
    .clk(clk100m),
    .d(\PWM9/n23 [28]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[28]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b29  (
    .clk(clk100m),
    .d(\PWM9/n23 [29]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[29]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b3  (
    .clk(clk100m),
    .d(\PWM9/n23 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[3]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b30  (
    .clk(clk100m),
    .d(\PWM9/n23 [30]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[30]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b31  (
    .clk(clk100m),
    .d(\PWM9/n23 [31]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[31]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b4  (
    .clk(clk100m),
    .d(\PWM9/n23 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[4]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b5  (
    .clk(clk100m),
    .d(\PWM9/n23 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[5]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b6  (
    .clk(clk100m),
    .d(\PWM9/n23 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[6]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b7  (
    .clk(clk100m),
    .d(\PWM9/n23 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[7]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b8  (
    .clk(clk100m),
    .d(\PWM9/n23 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[8]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b9  (
    .clk(clk100m),
    .d(\PWM9/n23 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[9]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg3_b0  (
    .clk(clk100m),
    .d(\PWM9/n31 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[0]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b1  (
    .clk(clk100m),
    .d(\PWM9/n31 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[1]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b10  (
    .clk(clk100m),
    .d(\PWM9/n31 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[10]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b11  (
    .clk(clk100m),
    .d(\PWM9/n31 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[11]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b12  (
    .clk(clk100m),
    .d(\PWM9/n31 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[12]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b13  (
    .clk(clk100m),
    .d(\PWM9/n31 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[13]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b14  (
    .clk(clk100m),
    .d(\PWM9/n31 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[14]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b15  (
    .clk(clk100m),
    .d(\PWM9/n31 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[15]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b16  (
    .clk(clk100m),
    .d(\PWM9/n31 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[16]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b17  (
    .clk(clk100m),
    .d(\PWM9/n31 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[17]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b18  (
    .clk(clk100m),
    .d(\PWM9/n31 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[18]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b19  (
    .clk(clk100m),
    .d(\PWM9/n31 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[19]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b2  (
    .clk(clk100m),
    .d(\PWM9/n31 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[2]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b20  (
    .clk(clk100m),
    .d(\PWM9/n31 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[20]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b21  (
    .clk(clk100m),
    .d(\PWM9/n31 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[21]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b22  (
    .clk(clk100m),
    .d(\PWM9/n31 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[22]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b23  (
    .clk(clk100m),
    .d(\PWM9/n31 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[23]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b3  (
    .clk(clk100m),
    .d(\PWM9/n31 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[3]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b4  (
    .clk(clk100m),
    .d(\PWM9/n31 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[4]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b5  (
    .clk(clk100m),
    .d(\PWM9/n31 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[5]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b6  (
    .clk(clk100m),
    .d(\PWM9/n31 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[6]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b7  (
    .clk(clk100m),
    .d(\PWM9/n31 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[7]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b8  (
    .clk(clk100m),
    .d(\PWM9/n31 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[8]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b9  (
    .clk(clk100m),
    .d(\PWM9/n31 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[9]_keep ));  // src/OnePWM.v(58)
  reg_ar_ss_w1 \PWM9/stopreq_reg  (
    .clk(clk100m),
    .d(\PWM9/n1 ),
    .en(1'b1),
    .reset(1'b0),
    .set(pwm_start_stop[9]),
    .q(\PWM9/stopreq_keep ));  // src/OnePWM.v(15)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub0/u0  (
    .a(\PWM9/FreCnt [0]),
    .b(1'b1),
    .c(\PWM9/sub0/c0 ),
    .o({\PWM9/sub0/c1 ,\PWM9/n12 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub0/u1  (
    .a(\PWM9/FreCnt [1]),
    .b(1'b0),
    .c(\PWM9/sub0/c1 ),
    .o({\PWM9/sub0/c2 ,\PWM9/n12 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub0/u10  (
    .a(\PWM9/FreCnt [10]),
    .b(1'b0),
    .c(\PWM9/sub0/c10 ),
    .o({\PWM9/sub0/c11 ,\PWM9/n12 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub0/u11  (
    .a(\PWM9/FreCnt [11]),
    .b(1'b0),
    .c(\PWM9/sub0/c11 ),
    .o({\PWM9/sub0/c12 ,\PWM9/n12 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub0/u12  (
    .a(\PWM9/FreCnt [12]),
    .b(1'b0),
    .c(\PWM9/sub0/c12 ),
    .o({\PWM9/sub0/c13 ,\PWM9/n12 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub0/u13  (
    .a(\PWM9/FreCnt [13]),
    .b(1'b0),
    .c(\PWM9/sub0/c13 ),
    .o({\PWM9/sub0/c14 ,\PWM9/n12 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub0/u14  (
    .a(\PWM9/FreCnt [14]),
    .b(1'b0),
    .c(\PWM9/sub0/c14 ),
    .o({\PWM9/sub0/c15 ,\PWM9/n12 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub0/u15  (
    .a(\PWM9/FreCnt [15]),
    .b(1'b0),
    .c(\PWM9/sub0/c15 ),
    .o({\PWM9/sub0/c16 ,\PWM9/n12 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub0/u16  (
    .a(\PWM9/FreCnt [16]),
    .b(1'b0),
    .c(\PWM9/sub0/c16 ),
    .o({\PWM9/sub0/c17 ,\PWM9/n12 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub0/u17  (
    .a(\PWM9/FreCnt [17]),
    .b(1'b0),
    .c(\PWM9/sub0/c17 ),
    .o({\PWM9/sub0/c18 ,\PWM9/n12 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub0/u18  (
    .a(\PWM9/FreCnt [18]),
    .b(1'b0),
    .c(\PWM9/sub0/c18 ),
    .o({\PWM9/sub0/c19 ,\PWM9/n12 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub0/u19  (
    .a(\PWM9/FreCnt [19]),
    .b(1'b0),
    .c(\PWM9/sub0/c19 ),
    .o({\PWM9/sub0/c20 ,\PWM9/n12 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub0/u2  (
    .a(\PWM9/FreCnt [2]),
    .b(1'b0),
    .c(\PWM9/sub0/c2 ),
    .o({\PWM9/sub0/c3 ,\PWM9/n12 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub0/u20  (
    .a(\PWM9/FreCnt [20]),
    .b(1'b0),
    .c(\PWM9/sub0/c20 ),
    .o({\PWM9/sub0/c21 ,\PWM9/n12 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub0/u21  (
    .a(\PWM9/FreCnt [21]),
    .b(1'b0),
    .c(\PWM9/sub0/c21 ),
    .o({\PWM9/sub0/c22 ,\PWM9/n12 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub0/u22  (
    .a(\PWM9/FreCnt [22]),
    .b(1'b0),
    .c(\PWM9/sub0/c22 ),
    .o({\PWM9/sub0/c23 ,\PWM9/n12 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub0/u23  (
    .a(\PWM9/FreCnt [23]),
    .b(1'b0),
    .c(\PWM9/sub0/c23 ),
    .o({\PWM9/sub0/c24 ,\PWM9/n12 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub0/u24  (
    .a(\PWM9/FreCnt [24]),
    .b(1'b0),
    .c(\PWM9/sub0/c24 ),
    .o({\PWM9/sub0/c25 ,\PWM9/n12 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub0/u25  (
    .a(\PWM9/FreCnt [25]),
    .b(1'b0),
    .c(\PWM9/sub0/c25 ),
    .o({\PWM9/sub0/c26 ,\PWM9/n12 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub0/u26  (
    .a(\PWM9/FreCnt [26]),
    .b(1'b0),
    .c(\PWM9/sub0/c26 ),
    .o({open_n72,\PWM9/n12 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub0/u3  (
    .a(\PWM9/FreCnt [3]),
    .b(1'b0),
    .c(\PWM9/sub0/c3 ),
    .o({\PWM9/sub0/c4 ,\PWM9/n12 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub0/u4  (
    .a(\PWM9/FreCnt [4]),
    .b(1'b0),
    .c(\PWM9/sub0/c4 ),
    .o({\PWM9/sub0/c5 ,\PWM9/n12 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub0/u5  (
    .a(\PWM9/FreCnt [5]),
    .b(1'b0),
    .c(\PWM9/sub0/c5 ),
    .o({\PWM9/sub0/c6 ,\PWM9/n12 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub0/u6  (
    .a(\PWM9/FreCnt [6]),
    .b(1'b0),
    .c(\PWM9/sub0/c6 ),
    .o({\PWM9/sub0/c7 ,\PWM9/n12 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub0/u7  (
    .a(\PWM9/FreCnt [7]),
    .b(1'b0),
    .c(\PWM9/sub0/c7 ),
    .o({\PWM9/sub0/c8 ,\PWM9/n12 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub0/u8  (
    .a(\PWM9/FreCnt [8]),
    .b(1'b0),
    .c(\PWM9/sub0/c8 ),
    .o({\PWM9/sub0/c9 ,\PWM9/n12 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub0/u9  (
    .a(\PWM9/FreCnt [9]),
    .b(1'b0),
    .c(\PWM9/sub0/c9 ),
    .o({\PWM9/sub0/c10 ,\PWM9/n12 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \PWM9/sub0/ucin  (
    .a(1'b0),
    .o({\PWM9/sub0/c0 ,open_n75}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub1/u0  (
    .a(pnumcnt9[0]),
    .b(1'b1),
    .c(\PWM9/sub1/c0 ),
    .o({\PWM9/sub1/c1 ,\PWM9/n26 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub1/u1  (
    .a(pnumcnt9[1]),
    .b(1'b0),
    .c(\PWM9/sub1/c1 ),
    .o({\PWM9/sub1/c2 ,\PWM9/n26 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub1/u10  (
    .a(pnumcnt9[10]),
    .b(1'b0),
    .c(\PWM9/sub1/c10 ),
    .o({\PWM9/sub1/c11 ,\PWM9/n26 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub1/u11  (
    .a(pnumcnt9[11]),
    .b(1'b0),
    .c(\PWM9/sub1/c11 ),
    .o({\PWM9/sub1/c12 ,\PWM9/n26 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub1/u12  (
    .a(pnumcnt9[12]),
    .b(1'b0),
    .c(\PWM9/sub1/c12 ),
    .o({\PWM9/sub1/c13 ,\PWM9/n26 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub1/u13  (
    .a(pnumcnt9[13]),
    .b(1'b0),
    .c(\PWM9/sub1/c13 ),
    .o({\PWM9/sub1/c14 ,\PWM9/n26 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub1/u14  (
    .a(pnumcnt9[14]),
    .b(1'b0),
    .c(\PWM9/sub1/c14 ),
    .o({\PWM9/sub1/c15 ,\PWM9/n26 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub1/u15  (
    .a(pnumcnt9[15]),
    .b(1'b0),
    .c(\PWM9/sub1/c15 ),
    .o({\PWM9/sub1/c16 ,\PWM9/n26 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub1/u16  (
    .a(pnumcnt9[16]),
    .b(1'b0),
    .c(\PWM9/sub1/c16 ),
    .o({\PWM9/sub1/c17 ,\PWM9/n26 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub1/u17  (
    .a(pnumcnt9[17]),
    .b(1'b0),
    .c(\PWM9/sub1/c17 ),
    .o({\PWM9/sub1/c18 ,\PWM9/n26 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub1/u18  (
    .a(pnumcnt9[18]),
    .b(1'b0),
    .c(\PWM9/sub1/c18 ),
    .o({\PWM9/sub1/c19 ,\PWM9/n26 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub1/u19  (
    .a(pnumcnt9[19]),
    .b(1'b0),
    .c(\PWM9/sub1/c19 ),
    .o({\PWM9/sub1/c20 ,\PWM9/n26 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub1/u2  (
    .a(pnumcnt9[2]),
    .b(1'b0),
    .c(\PWM9/sub1/c2 ),
    .o({\PWM9/sub1/c3 ,\PWM9/n26 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub1/u20  (
    .a(pnumcnt9[20]),
    .b(1'b0),
    .c(\PWM9/sub1/c20 ),
    .o({\PWM9/sub1/c21 ,\PWM9/n26 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub1/u21  (
    .a(pnumcnt9[21]),
    .b(1'b0),
    .c(\PWM9/sub1/c21 ),
    .o({\PWM9/sub1/c22 ,\PWM9/n26 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub1/u22  (
    .a(pnumcnt9[22]),
    .b(1'b0),
    .c(\PWM9/sub1/c22 ),
    .o({\PWM9/sub1/c23 ,\PWM9/n26 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub1/u23  (
    .a(pnumcnt9[23]),
    .b(1'b0),
    .c(\PWM9/sub1/c23 ),
    .o({open_n76,\PWM9/n26 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub1/u3  (
    .a(pnumcnt9[3]),
    .b(1'b0),
    .c(\PWM9/sub1/c3 ),
    .o({\PWM9/sub1/c4 ,\PWM9/n26 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub1/u4  (
    .a(pnumcnt9[4]),
    .b(1'b0),
    .c(\PWM9/sub1/c4 ),
    .o({\PWM9/sub1/c5 ,\PWM9/n26 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub1/u5  (
    .a(pnumcnt9[5]),
    .b(1'b0),
    .c(\PWM9/sub1/c5 ),
    .o({\PWM9/sub1/c6 ,\PWM9/n26 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub1/u6  (
    .a(pnumcnt9[6]),
    .b(1'b0),
    .c(\PWM9/sub1/c6 ),
    .o({\PWM9/sub1/c7 ,\PWM9/n26 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub1/u7  (
    .a(pnumcnt9[7]),
    .b(1'b0),
    .c(\PWM9/sub1/c7 ),
    .o({\PWM9/sub1/c8 ,\PWM9/n26 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub1/u8  (
    .a(pnumcnt9[8]),
    .b(1'b0),
    .c(\PWM9/sub1/c8 ),
    .o({\PWM9/sub1/c9 ,\PWM9/n26 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWM9/sub1/u9  (
    .a(pnumcnt9[9]),
    .b(1'b0),
    .c(\PWM9/sub1/c9 ),
    .o({\PWM9/sub1/c10 ,\PWM9/n26 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \PWM9/sub1/ucin  (
    .a(1'b0),
    .o({\PWM9/sub1/c0 ,open_n79}));
  reg_ar_as_w1 \PWMA/State_reg  (
    .clk(clk100m),
    .d(\PWMA/n10 ),
    .en(1'b1),
    .reset(~rstn),
    .set(1'b0),
    .q(pwm_state_read[10]));  // src/OnePWM.v(26)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[0]  (
    .i(\PWMA/RemaTxNum[0]_keep ),
    .o(pnumcntA[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[10]  (
    .i(\PWMA/RemaTxNum[10]_keep ),
    .o(pnumcntA[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[11]  (
    .i(\PWMA/RemaTxNum[11]_keep ),
    .o(pnumcntA[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[12]  (
    .i(\PWMA/RemaTxNum[12]_keep ),
    .o(pnumcntA[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[13]  (
    .i(\PWMA/RemaTxNum[13]_keep ),
    .o(pnumcntA[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[14]  (
    .i(\PWMA/RemaTxNum[14]_keep ),
    .o(pnumcntA[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[15]  (
    .i(\PWMA/RemaTxNum[15]_keep ),
    .o(pnumcntA[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[16]  (
    .i(\PWMA/RemaTxNum[16]_keep ),
    .o(pnumcntA[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[17]  (
    .i(\PWMA/RemaTxNum[17]_keep ),
    .o(pnumcntA[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[18]  (
    .i(\PWMA/RemaTxNum[18]_keep ),
    .o(pnumcntA[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[19]  (
    .i(\PWMA/RemaTxNum[19]_keep ),
    .o(pnumcntA[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[1]  (
    .i(\PWMA/RemaTxNum[1]_keep ),
    .o(pnumcntA[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[20]  (
    .i(\PWMA/RemaTxNum[20]_keep ),
    .o(pnumcntA[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[21]  (
    .i(\PWMA/RemaTxNum[21]_keep ),
    .o(pnumcntA[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[22]  (
    .i(\PWMA/RemaTxNum[22]_keep ),
    .o(pnumcntA[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[23]  (
    .i(\PWMA/RemaTxNum[23]_keep ),
    .o(pnumcntA[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[2]  (
    .i(\PWMA/RemaTxNum[2]_keep ),
    .o(pnumcntA[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[3]  (
    .i(\PWMA/RemaTxNum[3]_keep ),
    .o(pnumcntA[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[4]  (
    .i(\PWMA/RemaTxNum[4]_keep ),
    .o(pnumcntA[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[5]  (
    .i(\PWMA/RemaTxNum[5]_keep ),
    .o(pnumcntA[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[6]  (
    .i(\PWMA/RemaTxNum[6]_keep ),
    .o(pnumcntA[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[7]  (
    .i(\PWMA/RemaTxNum[7]_keep ),
    .o(pnumcntA[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[8]  (
    .i(\PWMA/RemaTxNum[8]_keep ),
    .o(pnumcntA[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[9]  (
    .i(\PWMA/RemaTxNum[9]_keep ),
    .o(pnumcntA[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_dir  (
    .i(\PWMA/dir_keep ),
    .o(dir_pad[10]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[0]  (
    .i(\PWMA/pnumr[0]_keep ),
    .o(\PWMA/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[10]  (
    .i(\PWMA/pnumr[10]_keep ),
    .o(\PWMA/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[11]  (
    .i(\PWMA/pnumr[11]_keep ),
    .o(\PWMA/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[12]  (
    .i(\PWMA/pnumr[12]_keep ),
    .o(\PWMA/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[13]  (
    .i(\PWMA/pnumr[13]_keep ),
    .o(\PWMA/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[14]  (
    .i(\PWMA/pnumr[14]_keep ),
    .o(\PWMA/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[15]  (
    .i(\PWMA/pnumr[15]_keep ),
    .o(\PWMA/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[16]  (
    .i(\PWMA/pnumr[16]_keep ),
    .o(\PWMA/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[17]  (
    .i(\PWMA/pnumr[17]_keep ),
    .o(\PWMA/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[18]  (
    .i(\PWMA/pnumr[18]_keep ),
    .o(\PWMA/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[19]  (
    .i(\PWMA/pnumr[19]_keep ),
    .o(\PWMA/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[1]  (
    .i(\PWMA/pnumr[1]_keep ),
    .o(\PWMA/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[20]  (
    .i(\PWMA/pnumr[20]_keep ),
    .o(\PWMA/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[21]  (
    .i(\PWMA/pnumr[21]_keep ),
    .o(\PWMA/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[22]  (
    .i(\PWMA/pnumr[22]_keep ),
    .o(\PWMA/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[23]  (
    .i(\PWMA/pnumr[23]_keep ),
    .o(\PWMA/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[24]  (
    .i(\PWMA/pnumr[24]_keep ),
    .o(\PWMA/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[25]  (
    .i(\PWMA/pnumr[25]_keep ),
    .o(\PWMA/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[26]  (
    .i(\PWMA/pnumr[26]_keep ),
    .o(\PWMA/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[27]  (
    .i(\PWMA/pnumr[27]_keep ),
    .o(\PWMA/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[28]  (
    .i(\PWMA/pnumr[28]_keep ),
    .o(\PWMA/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[29]  (
    .i(\PWMA/pnumr[29]_keep ),
    .o(\PWMA/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[2]  (
    .i(\PWMA/pnumr[2]_keep ),
    .o(\PWMA/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[30]  (
    .i(\PWMA/pnumr[30]_keep ),
    .o(\PWMA/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[31]  (
    .i(\PWMA/pnumr[31]_keep ),
    .o(\PWMA/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[3]  (
    .i(\PWMA/pnumr[3]_keep ),
    .o(\PWMA/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[4]  (
    .i(\PWMA/pnumr[4]_keep ),
    .o(\PWMA/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[5]  (
    .i(\PWMA/pnumr[5]_keep ),
    .o(\PWMA/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[6]  (
    .i(\PWMA/pnumr[6]_keep ),
    .o(\PWMA/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[7]  (
    .i(\PWMA/pnumr[7]_keep ),
    .o(\PWMA/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[8]  (
    .i(\PWMA/pnumr[8]_keep ),
    .o(\PWMA/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[9]  (
    .i(\PWMA/pnumr[9]_keep ),
    .o(\PWMA/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pwm  (
    .i(\PWMA/pwm_keep ),
    .o(pwm_pad[10]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_stopreq  (
    .i(\PWMA/stopreq_keep ),
    .o(\PWMA/stopreq ));  // src/OnePWM.v(14)
  reg_ar_as_w1 \PWMA/dir_reg  (
    .clk(clk100m),
    .d(\PWMA/n32 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/dir_keep ));  // src/OnePWM.v(58)
  reg_sr_as_w1 \PWMA/pwm_reg  (
    .clk(clk100m),
    .d(\pwm[10]_d ),
    .en(1'b1),
    .reset(~\PWMA/u14_sel_is_1_o ),
    .set(1'b0),
    .q(\PWMA/pwm_keep ));  // src/OnePWM.v(45)
  reg_sr_as_w1 \PWMA/reg0_b0  (
    .clk(clk100m),
    .d(\PWMA/n13 [0]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [0]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b1  (
    .clk(clk100m),
    .d(\PWMA/n13 [1]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [1]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b10  (
    .clk(clk100m),
    .d(\PWMA/n13 [10]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [10]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b11  (
    .clk(clk100m),
    .d(\PWMA/n13 [11]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [11]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b12  (
    .clk(clk100m),
    .d(\PWMA/n13 [12]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [12]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b13  (
    .clk(clk100m),
    .d(\PWMA/n13 [13]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [13]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b14  (
    .clk(clk100m),
    .d(\PWMA/n13 [14]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [14]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b15  (
    .clk(clk100m),
    .d(\PWMA/n13 [15]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [15]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b16  (
    .clk(clk100m),
    .d(\PWMA/n13 [16]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [16]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b17  (
    .clk(clk100m),
    .d(\PWMA/n13 [17]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [17]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b18  (
    .clk(clk100m),
    .d(\PWMA/n13 [18]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [18]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b19  (
    .clk(clk100m),
    .d(\PWMA/n13 [19]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [19]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b2  (
    .clk(clk100m),
    .d(\PWMA/n13 [2]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [2]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b20  (
    .clk(clk100m),
    .d(\PWMA/n13 [20]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [20]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b21  (
    .clk(clk100m),
    .d(\PWMA/n13 [21]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [21]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b22  (
    .clk(clk100m),
    .d(\PWMA/n13 [22]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [22]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b23  (
    .clk(clk100m),
    .d(\PWMA/n13 [23]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [23]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b24  (
    .clk(clk100m),
    .d(\PWMA/n13 [24]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [24]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b25  (
    .clk(clk100m),
    .d(\PWMA/n13 [25]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [25]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b26  (
    .clk(clk100m),
    .d(\PWMA/n13 [26]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [26]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b3  (
    .clk(clk100m),
    .d(\PWMA/n13 [3]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [3]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b4  (
    .clk(clk100m),
    .d(\PWMA/n13 [4]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [4]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b5  (
    .clk(clk100m),
    .d(\PWMA/n13 [5]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [5]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b6  (
    .clk(clk100m),
    .d(\PWMA/n13 [6]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [6]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b7  (
    .clk(clk100m),
    .d(\PWMA/n13 [7]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [7]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b8  (
    .clk(clk100m),
    .d(\PWMA/n13 [8]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [8]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b9  (
    .clk(clk100m),
    .d(\PWMA/n13 [9]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b0  (
    .clk(clk100m),
    .d(freqA[0]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [0]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b1  (
    .clk(clk100m),
    .d(freqA[1]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [1]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b10  (
    .clk(clk100m),
    .d(freqA[10]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [10]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b11  (
    .clk(clk100m),
    .d(freqA[11]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [11]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b12  (
    .clk(clk100m),
    .d(freqA[12]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [12]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b13  (
    .clk(clk100m),
    .d(freqA[13]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [13]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b14  (
    .clk(clk100m),
    .d(freqA[14]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [14]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b15  (
    .clk(clk100m),
    .d(freqA[15]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [15]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b16  (
    .clk(clk100m),
    .d(freqA[16]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [16]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b17  (
    .clk(clk100m),
    .d(freqA[17]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [17]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b18  (
    .clk(clk100m),
    .d(freqA[18]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [18]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b19  (
    .clk(clk100m),
    .d(freqA[19]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [19]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b2  (
    .clk(clk100m),
    .d(freqA[2]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [2]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b20  (
    .clk(clk100m),
    .d(freqA[20]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [20]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b21  (
    .clk(clk100m),
    .d(freqA[21]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [21]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b22  (
    .clk(clk100m),
    .d(freqA[22]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [22]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b23  (
    .clk(clk100m),
    .d(freqA[23]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [23]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b24  (
    .clk(clk100m),
    .d(freqA[24]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [24]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b25  (
    .clk(clk100m),
    .d(freqA[25]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [25]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b26  (
    .clk(clk100m),
    .d(freqA[26]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [26]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b3  (
    .clk(clk100m),
    .d(freqA[3]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [3]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b4  (
    .clk(clk100m),
    .d(freqA[4]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [4]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b5  (
    .clk(clk100m),
    .d(freqA[5]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [5]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b6  (
    .clk(clk100m),
    .d(freqA[6]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [6]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b7  (
    .clk(clk100m),
    .d(freqA[7]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [7]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b8  (
    .clk(clk100m),
    .d(freqA[8]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [8]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b9  (
    .clk(clk100m),
    .d(freqA[9]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg2_b0  (
    .clk(clk100m),
    .d(\PWMA/n23 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[0]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b1  (
    .clk(clk100m),
    .d(\PWMA/n23 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[1]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b10  (
    .clk(clk100m),
    .d(\PWMA/n23 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[10]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b11  (
    .clk(clk100m),
    .d(\PWMA/n23 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[11]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b12  (
    .clk(clk100m),
    .d(\PWMA/n23 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[12]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b13  (
    .clk(clk100m),
    .d(\PWMA/n23 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[13]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b14  (
    .clk(clk100m),
    .d(\PWMA/n23 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[14]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b15  (
    .clk(clk100m),
    .d(\PWMA/n23 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[15]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b16  (
    .clk(clk100m),
    .d(\PWMA/n23 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[16]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b17  (
    .clk(clk100m),
    .d(\PWMA/n23 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[17]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b18  (
    .clk(clk100m),
    .d(\PWMA/n23 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[18]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b19  (
    .clk(clk100m),
    .d(\PWMA/n23 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[19]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b2  (
    .clk(clk100m),
    .d(\PWMA/n23 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[2]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b20  (
    .clk(clk100m),
    .d(\PWMA/n23 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[20]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b21  (
    .clk(clk100m),
    .d(\PWMA/n23 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[21]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b22  (
    .clk(clk100m),
    .d(\PWMA/n23 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[22]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b23  (
    .clk(clk100m),
    .d(\PWMA/n23 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[23]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b24  (
    .clk(clk100m),
    .d(\PWMA/n23 [24]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[24]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b25  (
    .clk(clk100m),
    .d(\PWMA/n23 [25]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[25]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b26  (
    .clk(clk100m),
    .d(\PWMA/n23 [26]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[26]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b27  (
    .clk(clk100m),
    .d(\PWMA/n23 [27]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[27]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b28  (
    .clk(clk100m),
    .d(\PWMA/n23 [28]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[28]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b29  (
    .clk(clk100m),
    .d(\PWMA/n23 [29]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[29]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b3  (
    .clk(clk100m),
    .d(\PWMA/n23 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[3]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b30  (
    .clk(clk100m),
    .d(\PWMA/n23 [30]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[30]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b31  (
    .clk(clk100m),
    .d(\PWMA/n23 [31]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[31]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b4  (
    .clk(clk100m),
    .d(\PWMA/n23 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[4]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b5  (
    .clk(clk100m),
    .d(\PWMA/n23 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[5]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b6  (
    .clk(clk100m),
    .d(\PWMA/n23 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[6]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b7  (
    .clk(clk100m),
    .d(\PWMA/n23 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[7]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b8  (
    .clk(clk100m),
    .d(\PWMA/n23 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[8]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b9  (
    .clk(clk100m),
    .d(\PWMA/n23 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[9]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg3_b0  (
    .clk(clk100m),
    .d(\PWMA/n31 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[0]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b1  (
    .clk(clk100m),
    .d(\PWMA/n31 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[1]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b10  (
    .clk(clk100m),
    .d(\PWMA/n31 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[10]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b11  (
    .clk(clk100m),
    .d(\PWMA/n31 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[11]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b12  (
    .clk(clk100m),
    .d(\PWMA/n31 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[12]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b13  (
    .clk(clk100m),
    .d(\PWMA/n31 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[13]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b14  (
    .clk(clk100m),
    .d(\PWMA/n31 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[14]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b15  (
    .clk(clk100m),
    .d(\PWMA/n31 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[15]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b16  (
    .clk(clk100m),
    .d(\PWMA/n31 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[16]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b17  (
    .clk(clk100m),
    .d(\PWMA/n31 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[17]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b18  (
    .clk(clk100m),
    .d(\PWMA/n31 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[18]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b19  (
    .clk(clk100m),
    .d(\PWMA/n31 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[19]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b2  (
    .clk(clk100m),
    .d(\PWMA/n31 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[2]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b20  (
    .clk(clk100m),
    .d(\PWMA/n31 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[20]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b21  (
    .clk(clk100m),
    .d(\PWMA/n31 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[21]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b22  (
    .clk(clk100m),
    .d(\PWMA/n31 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[22]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b23  (
    .clk(clk100m),
    .d(\PWMA/n31 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[23]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b3  (
    .clk(clk100m),
    .d(\PWMA/n31 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[3]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b4  (
    .clk(clk100m),
    .d(\PWMA/n31 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[4]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b5  (
    .clk(clk100m),
    .d(\PWMA/n31 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[5]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b6  (
    .clk(clk100m),
    .d(\PWMA/n31 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[6]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b7  (
    .clk(clk100m),
    .d(\PWMA/n31 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[7]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b8  (
    .clk(clk100m),
    .d(\PWMA/n31 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[8]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b9  (
    .clk(clk100m),
    .d(\PWMA/n31 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[9]_keep ));  // src/OnePWM.v(58)
  reg_ar_ss_w1 \PWMA/stopreq_reg  (
    .clk(clk100m),
    .d(\PWMA/n1 ),
    .en(1'b1),
    .reset(1'b0),
    .set(pwm_start_stop[10]),
    .q(\PWMA/stopreq_keep ));  // src/OnePWM.v(15)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub0/u0  (
    .a(\PWMA/FreCnt [0]),
    .b(1'b1),
    .c(\PWMA/sub0/c0 ),
    .o({\PWMA/sub0/c1 ,\PWMA/n12 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub0/u1  (
    .a(\PWMA/FreCnt [1]),
    .b(1'b0),
    .c(\PWMA/sub0/c1 ),
    .o({\PWMA/sub0/c2 ,\PWMA/n12 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub0/u10  (
    .a(\PWMA/FreCnt [10]),
    .b(1'b0),
    .c(\PWMA/sub0/c10 ),
    .o({\PWMA/sub0/c11 ,\PWMA/n12 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub0/u11  (
    .a(\PWMA/FreCnt [11]),
    .b(1'b0),
    .c(\PWMA/sub0/c11 ),
    .o({\PWMA/sub0/c12 ,\PWMA/n12 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub0/u12  (
    .a(\PWMA/FreCnt [12]),
    .b(1'b0),
    .c(\PWMA/sub0/c12 ),
    .o({\PWMA/sub0/c13 ,\PWMA/n12 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub0/u13  (
    .a(\PWMA/FreCnt [13]),
    .b(1'b0),
    .c(\PWMA/sub0/c13 ),
    .o({\PWMA/sub0/c14 ,\PWMA/n12 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub0/u14  (
    .a(\PWMA/FreCnt [14]),
    .b(1'b0),
    .c(\PWMA/sub0/c14 ),
    .o({\PWMA/sub0/c15 ,\PWMA/n12 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub0/u15  (
    .a(\PWMA/FreCnt [15]),
    .b(1'b0),
    .c(\PWMA/sub0/c15 ),
    .o({\PWMA/sub0/c16 ,\PWMA/n12 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub0/u16  (
    .a(\PWMA/FreCnt [16]),
    .b(1'b0),
    .c(\PWMA/sub0/c16 ),
    .o({\PWMA/sub0/c17 ,\PWMA/n12 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub0/u17  (
    .a(\PWMA/FreCnt [17]),
    .b(1'b0),
    .c(\PWMA/sub0/c17 ),
    .o({\PWMA/sub0/c18 ,\PWMA/n12 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub0/u18  (
    .a(\PWMA/FreCnt [18]),
    .b(1'b0),
    .c(\PWMA/sub0/c18 ),
    .o({\PWMA/sub0/c19 ,\PWMA/n12 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub0/u19  (
    .a(\PWMA/FreCnt [19]),
    .b(1'b0),
    .c(\PWMA/sub0/c19 ),
    .o({\PWMA/sub0/c20 ,\PWMA/n12 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub0/u2  (
    .a(\PWMA/FreCnt [2]),
    .b(1'b0),
    .c(\PWMA/sub0/c2 ),
    .o({\PWMA/sub0/c3 ,\PWMA/n12 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub0/u20  (
    .a(\PWMA/FreCnt [20]),
    .b(1'b0),
    .c(\PWMA/sub0/c20 ),
    .o({\PWMA/sub0/c21 ,\PWMA/n12 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub0/u21  (
    .a(\PWMA/FreCnt [21]),
    .b(1'b0),
    .c(\PWMA/sub0/c21 ),
    .o({\PWMA/sub0/c22 ,\PWMA/n12 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub0/u22  (
    .a(\PWMA/FreCnt [22]),
    .b(1'b0),
    .c(\PWMA/sub0/c22 ),
    .o({\PWMA/sub0/c23 ,\PWMA/n12 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub0/u23  (
    .a(\PWMA/FreCnt [23]),
    .b(1'b0),
    .c(\PWMA/sub0/c23 ),
    .o({\PWMA/sub0/c24 ,\PWMA/n12 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub0/u24  (
    .a(\PWMA/FreCnt [24]),
    .b(1'b0),
    .c(\PWMA/sub0/c24 ),
    .o({\PWMA/sub0/c25 ,\PWMA/n12 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub0/u25  (
    .a(\PWMA/FreCnt [25]),
    .b(1'b0),
    .c(\PWMA/sub0/c25 ),
    .o({\PWMA/sub0/c26 ,\PWMA/n12 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub0/u26  (
    .a(\PWMA/FreCnt [26]),
    .b(1'b0),
    .c(\PWMA/sub0/c26 ),
    .o({open_n80,\PWMA/n12 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub0/u3  (
    .a(\PWMA/FreCnt [3]),
    .b(1'b0),
    .c(\PWMA/sub0/c3 ),
    .o({\PWMA/sub0/c4 ,\PWMA/n12 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub0/u4  (
    .a(\PWMA/FreCnt [4]),
    .b(1'b0),
    .c(\PWMA/sub0/c4 ),
    .o({\PWMA/sub0/c5 ,\PWMA/n12 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub0/u5  (
    .a(\PWMA/FreCnt [5]),
    .b(1'b0),
    .c(\PWMA/sub0/c5 ),
    .o({\PWMA/sub0/c6 ,\PWMA/n12 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub0/u6  (
    .a(\PWMA/FreCnt [6]),
    .b(1'b0),
    .c(\PWMA/sub0/c6 ),
    .o({\PWMA/sub0/c7 ,\PWMA/n12 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub0/u7  (
    .a(\PWMA/FreCnt [7]),
    .b(1'b0),
    .c(\PWMA/sub0/c7 ),
    .o({\PWMA/sub0/c8 ,\PWMA/n12 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub0/u8  (
    .a(\PWMA/FreCnt [8]),
    .b(1'b0),
    .c(\PWMA/sub0/c8 ),
    .o({\PWMA/sub0/c9 ,\PWMA/n12 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub0/u9  (
    .a(\PWMA/FreCnt [9]),
    .b(1'b0),
    .c(\PWMA/sub0/c9 ),
    .o({\PWMA/sub0/c10 ,\PWMA/n12 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \PWMA/sub0/ucin  (
    .a(1'b0),
    .o({\PWMA/sub0/c0 ,open_n83}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub1/u0  (
    .a(pnumcntA[0]),
    .b(1'b1),
    .c(\PWMA/sub1/c0 ),
    .o({\PWMA/sub1/c1 ,\PWMA/n26 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub1/u1  (
    .a(pnumcntA[1]),
    .b(1'b0),
    .c(\PWMA/sub1/c1 ),
    .o({\PWMA/sub1/c2 ,\PWMA/n26 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub1/u10  (
    .a(pnumcntA[10]),
    .b(1'b0),
    .c(\PWMA/sub1/c10 ),
    .o({\PWMA/sub1/c11 ,\PWMA/n26 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub1/u11  (
    .a(pnumcntA[11]),
    .b(1'b0),
    .c(\PWMA/sub1/c11 ),
    .o({\PWMA/sub1/c12 ,\PWMA/n26 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub1/u12  (
    .a(pnumcntA[12]),
    .b(1'b0),
    .c(\PWMA/sub1/c12 ),
    .o({\PWMA/sub1/c13 ,\PWMA/n26 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub1/u13  (
    .a(pnumcntA[13]),
    .b(1'b0),
    .c(\PWMA/sub1/c13 ),
    .o({\PWMA/sub1/c14 ,\PWMA/n26 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub1/u14  (
    .a(pnumcntA[14]),
    .b(1'b0),
    .c(\PWMA/sub1/c14 ),
    .o({\PWMA/sub1/c15 ,\PWMA/n26 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub1/u15  (
    .a(pnumcntA[15]),
    .b(1'b0),
    .c(\PWMA/sub1/c15 ),
    .o({\PWMA/sub1/c16 ,\PWMA/n26 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub1/u16  (
    .a(pnumcntA[16]),
    .b(1'b0),
    .c(\PWMA/sub1/c16 ),
    .o({\PWMA/sub1/c17 ,\PWMA/n26 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub1/u17  (
    .a(pnumcntA[17]),
    .b(1'b0),
    .c(\PWMA/sub1/c17 ),
    .o({\PWMA/sub1/c18 ,\PWMA/n26 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub1/u18  (
    .a(pnumcntA[18]),
    .b(1'b0),
    .c(\PWMA/sub1/c18 ),
    .o({\PWMA/sub1/c19 ,\PWMA/n26 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub1/u19  (
    .a(pnumcntA[19]),
    .b(1'b0),
    .c(\PWMA/sub1/c19 ),
    .o({\PWMA/sub1/c20 ,\PWMA/n26 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub1/u2  (
    .a(pnumcntA[2]),
    .b(1'b0),
    .c(\PWMA/sub1/c2 ),
    .o({\PWMA/sub1/c3 ,\PWMA/n26 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub1/u20  (
    .a(pnumcntA[20]),
    .b(1'b0),
    .c(\PWMA/sub1/c20 ),
    .o({\PWMA/sub1/c21 ,\PWMA/n26 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub1/u21  (
    .a(pnumcntA[21]),
    .b(1'b0),
    .c(\PWMA/sub1/c21 ),
    .o({\PWMA/sub1/c22 ,\PWMA/n26 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub1/u22  (
    .a(pnumcntA[22]),
    .b(1'b0),
    .c(\PWMA/sub1/c22 ),
    .o({\PWMA/sub1/c23 ,\PWMA/n26 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub1/u23  (
    .a(pnumcntA[23]),
    .b(1'b0),
    .c(\PWMA/sub1/c23 ),
    .o({open_n84,\PWMA/n26 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub1/u3  (
    .a(pnumcntA[3]),
    .b(1'b0),
    .c(\PWMA/sub1/c3 ),
    .o({\PWMA/sub1/c4 ,\PWMA/n26 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub1/u4  (
    .a(pnumcntA[4]),
    .b(1'b0),
    .c(\PWMA/sub1/c4 ),
    .o({\PWMA/sub1/c5 ,\PWMA/n26 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub1/u5  (
    .a(pnumcntA[5]),
    .b(1'b0),
    .c(\PWMA/sub1/c5 ),
    .o({\PWMA/sub1/c6 ,\PWMA/n26 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub1/u6  (
    .a(pnumcntA[6]),
    .b(1'b0),
    .c(\PWMA/sub1/c6 ),
    .o({\PWMA/sub1/c7 ,\PWMA/n26 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub1/u7  (
    .a(pnumcntA[7]),
    .b(1'b0),
    .c(\PWMA/sub1/c7 ),
    .o({\PWMA/sub1/c8 ,\PWMA/n26 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub1/u8  (
    .a(pnumcntA[8]),
    .b(1'b0),
    .c(\PWMA/sub1/c8 ),
    .o({\PWMA/sub1/c9 ,\PWMA/n26 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMA/sub1/u9  (
    .a(pnumcntA[9]),
    .b(1'b0),
    .c(\PWMA/sub1/c9 ),
    .o({\PWMA/sub1/c10 ,\PWMA/n26 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \PWMA/sub1/ucin  (
    .a(1'b0),
    .o({\PWMA/sub1/c0 ,open_n87}));
  reg_ar_as_w1 \PWMB/State_reg  (
    .clk(clk100m),
    .d(\PWMB/n10 ),
    .en(1'b1),
    .reset(~rstn),
    .set(1'b0),
    .q(pwm_state_read[11]));  // src/OnePWM.v(26)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[0]  (
    .i(\PWMB/RemaTxNum[0]_keep ),
    .o(pnumcntB[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[10]  (
    .i(\PWMB/RemaTxNum[10]_keep ),
    .o(pnumcntB[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[11]  (
    .i(\PWMB/RemaTxNum[11]_keep ),
    .o(pnumcntB[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[12]  (
    .i(\PWMB/RemaTxNum[12]_keep ),
    .o(pnumcntB[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[13]  (
    .i(\PWMB/RemaTxNum[13]_keep ),
    .o(pnumcntB[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[14]  (
    .i(\PWMB/RemaTxNum[14]_keep ),
    .o(pnumcntB[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[15]  (
    .i(\PWMB/RemaTxNum[15]_keep ),
    .o(pnumcntB[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[16]  (
    .i(\PWMB/RemaTxNum[16]_keep ),
    .o(pnumcntB[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[17]  (
    .i(\PWMB/RemaTxNum[17]_keep ),
    .o(pnumcntB[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[18]  (
    .i(\PWMB/RemaTxNum[18]_keep ),
    .o(pnumcntB[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[19]  (
    .i(\PWMB/RemaTxNum[19]_keep ),
    .o(pnumcntB[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[1]  (
    .i(\PWMB/RemaTxNum[1]_keep ),
    .o(pnumcntB[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[20]  (
    .i(\PWMB/RemaTxNum[20]_keep ),
    .o(pnumcntB[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[21]  (
    .i(\PWMB/RemaTxNum[21]_keep ),
    .o(pnumcntB[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[22]  (
    .i(\PWMB/RemaTxNum[22]_keep ),
    .o(pnumcntB[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[23]  (
    .i(\PWMB/RemaTxNum[23]_keep ),
    .o(pnumcntB[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[2]  (
    .i(\PWMB/RemaTxNum[2]_keep ),
    .o(pnumcntB[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[3]  (
    .i(\PWMB/RemaTxNum[3]_keep ),
    .o(pnumcntB[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[4]  (
    .i(\PWMB/RemaTxNum[4]_keep ),
    .o(pnumcntB[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[5]  (
    .i(\PWMB/RemaTxNum[5]_keep ),
    .o(pnumcntB[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[6]  (
    .i(\PWMB/RemaTxNum[6]_keep ),
    .o(pnumcntB[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[7]  (
    .i(\PWMB/RemaTxNum[7]_keep ),
    .o(pnumcntB[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[8]  (
    .i(\PWMB/RemaTxNum[8]_keep ),
    .o(pnumcntB[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[9]  (
    .i(\PWMB/RemaTxNum[9]_keep ),
    .o(pnumcntB[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_dir  (
    .i(\PWMB/dir_keep ),
    .o(dir_pad[11]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[0]  (
    .i(\PWMB/pnumr[0]_keep ),
    .o(\PWMB/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[10]  (
    .i(\PWMB/pnumr[10]_keep ),
    .o(\PWMB/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[11]  (
    .i(\PWMB/pnumr[11]_keep ),
    .o(\PWMB/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[12]  (
    .i(\PWMB/pnumr[12]_keep ),
    .o(\PWMB/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[13]  (
    .i(\PWMB/pnumr[13]_keep ),
    .o(\PWMB/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[14]  (
    .i(\PWMB/pnumr[14]_keep ),
    .o(\PWMB/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[15]  (
    .i(\PWMB/pnumr[15]_keep ),
    .o(\PWMB/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[16]  (
    .i(\PWMB/pnumr[16]_keep ),
    .o(\PWMB/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[17]  (
    .i(\PWMB/pnumr[17]_keep ),
    .o(\PWMB/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[18]  (
    .i(\PWMB/pnumr[18]_keep ),
    .o(\PWMB/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[19]  (
    .i(\PWMB/pnumr[19]_keep ),
    .o(\PWMB/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[1]  (
    .i(\PWMB/pnumr[1]_keep ),
    .o(\PWMB/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[20]  (
    .i(\PWMB/pnumr[20]_keep ),
    .o(\PWMB/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[21]  (
    .i(\PWMB/pnumr[21]_keep ),
    .o(\PWMB/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[22]  (
    .i(\PWMB/pnumr[22]_keep ),
    .o(\PWMB/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[23]  (
    .i(\PWMB/pnumr[23]_keep ),
    .o(\PWMB/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[24]  (
    .i(\PWMB/pnumr[24]_keep ),
    .o(\PWMB/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[25]  (
    .i(\PWMB/pnumr[25]_keep ),
    .o(\PWMB/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[26]  (
    .i(\PWMB/pnumr[26]_keep ),
    .o(\PWMB/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[27]  (
    .i(\PWMB/pnumr[27]_keep ),
    .o(\PWMB/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[28]  (
    .i(\PWMB/pnumr[28]_keep ),
    .o(\PWMB/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[29]  (
    .i(\PWMB/pnumr[29]_keep ),
    .o(\PWMB/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[2]  (
    .i(\PWMB/pnumr[2]_keep ),
    .o(\PWMB/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[30]  (
    .i(\PWMB/pnumr[30]_keep ),
    .o(\PWMB/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[31]  (
    .i(\PWMB/pnumr[31]_keep ),
    .o(\PWMB/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[3]  (
    .i(\PWMB/pnumr[3]_keep ),
    .o(\PWMB/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[4]  (
    .i(\PWMB/pnumr[4]_keep ),
    .o(\PWMB/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[5]  (
    .i(\PWMB/pnumr[5]_keep ),
    .o(\PWMB/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[6]  (
    .i(\PWMB/pnumr[6]_keep ),
    .o(\PWMB/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[7]  (
    .i(\PWMB/pnumr[7]_keep ),
    .o(\PWMB/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[8]  (
    .i(\PWMB/pnumr[8]_keep ),
    .o(\PWMB/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[9]  (
    .i(\PWMB/pnumr[9]_keep ),
    .o(\PWMB/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pwm  (
    .i(\PWMB/pwm_keep ),
    .o(pwm_pad[11]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_stopreq  (
    .i(\PWMB/stopreq_keep ),
    .o(\PWMB/stopreq ));  // src/OnePWM.v(14)
  reg_ar_as_w1 \PWMB/dir_reg  (
    .clk(clk100m),
    .d(\PWMB/n32 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/dir_keep ));  // src/OnePWM.v(58)
  reg_sr_as_w1 \PWMB/pwm_reg  (
    .clk(clk100m),
    .d(\pwm[11]_d ),
    .en(1'b1),
    .reset(~\PWMB/u14_sel_is_1_o ),
    .set(1'b0),
    .q(\PWMB/pwm_keep ));  // src/OnePWM.v(45)
  reg_sr_as_w1 \PWMB/reg0_b0  (
    .clk(clk100m),
    .d(\PWMB/n13 [0]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [0]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b1  (
    .clk(clk100m),
    .d(\PWMB/n13 [1]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [1]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b10  (
    .clk(clk100m),
    .d(\PWMB/n13 [10]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [10]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b11  (
    .clk(clk100m),
    .d(\PWMB/n13 [11]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [11]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b12  (
    .clk(clk100m),
    .d(\PWMB/n13 [12]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [12]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b13  (
    .clk(clk100m),
    .d(\PWMB/n13 [13]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [13]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b14  (
    .clk(clk100m),
    .d(\PWMB/n13 [14]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [14]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b15  (
    .clk(clk100m),
    .d(\PWMB/n13 [15]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [15]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b16  (
    .clk(clk100m),
    .d(\PWMB/n13 [16]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [16]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b17  (
    .clk(clk100m),
    .d(\PWMB/n13 [17]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [17]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b18  (
    .clk(clk100m),
    .d(\PWMB/n13 [18]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [18]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b19  (
    .clk(clk100m),
    .d(\PWMB/n13 [19]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [19]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b2  (
    .clk(clk100m),
    .d(\PWMB/n13 [2]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [2]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b20  (
    .clk(clk100m),
    .d(\PWMB/n13 [20]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [20]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b21  (
    .clk(clk100m),
    .d(\PWMB/n13 [21]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [21]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b22  (
    .clk(clk100m),
    .d(\PWMB/n13 [22]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [22]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b23  (
    .clk(clk100m),
    .d(\PWMB/n13 [23]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [23]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b24  (
    .clk(clk100m),
    .d(\PWMB/n13 [24]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [24]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b25  (
    .clk(clk100m),
    .d(\PWMB/n13 [25]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [25]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b26  (
    .clk(clk100m),
    .d(\PWMB/n13 [26]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [26]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b3  (
    .clk(clk100m),
    .d(\PWMB/n13 [3]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [3]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b4  (
    .clk(clk100m),
    .d(\PWMB/n13 [4]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [4]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b5  (
    .clk(clk100m),
    .d(\PWMB/n13 [5]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [5]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b6  (
    .clk(clk100m),
    .d(\PWMB/n13 [6]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [6]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b7  (
    .clk(clk100m),
    .d(\PWMB/n13 [7]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [7]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b8  (
    .clk(clk100m),
    .d(\PWMB/n13 [8]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [8]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b9  (
    .clk(clk100m),
    .d(\PWMB/n13 [9]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b0  (
    .clk(clk100m),
    .d(freqB[0]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [0]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b1  (
    .clk(clk100m),
    .d(freqB[1]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [1]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b10  (
    .clk(clk100m),
    .d(freqB[10]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [10]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b11  (
    .clk(clk100m),
    .d(freqB[11]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [11]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b12  (
    .clk(clk100m),
    .d(freqB[12]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [12]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b13  (
    .clk(clk100m),
    .d(freqB[13]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [13]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b14  (
    .clk(clk100m),
    .d(freqB[14]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [14]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b15  (
    .clk(clk100m),
    .d(freqB[15]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [15]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b16  (
    .clk(clk100m),
    .d(freqB[16]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [16]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b17  (
    .clk(clk100m),
    .d(freqB[17]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [17]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b18  (
    .clk(clk100m),
    .d(freqB[18]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [18]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b19  (
    .clk(clk100m),
    .d(freqB[19]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [19]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b2  (
    .clk(clk100m),
    .d(freqB[2]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [2]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b20  (
    .clk(clk100m),
    .d(freqB[20]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [20]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b21  (
    .clk(clk100m),
    .d(freqB[21]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [21]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b22  (
    .clk(clk100m),
    .d(freqB[22]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [22]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b23  (
    .clk(clk100m),
    .d(freqB[23]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [23]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b24  (
    .clk(clk100m),
    .d(freqB[24]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [24]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b25  (
    .clk(clk100m),
    .d(freqB[25]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [25]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b26  (
    .clk(clk100m),
    .d(freqB[26]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [26]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b3  (
    .clk(clk100m),
    .d(freqB[3]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [3]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b4  (
    .clk(clk100m),
    .d(freqB[4]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [4]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b5  (
    .clk(clk100m),
    .d(freqB[5]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [5]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b6  (
    .clk(clk100m),
    .d(freqB[6]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [6]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b7  (
    .clk(clk100m),
    .d(freqB[7]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [7]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b8  (
    .clk(clk100m),
    .d(freqB[8]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [8]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b9  (
    .clk(clk100m),
    .d(freqB[9]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg2_b0  (
    .clk(clk100m),
    .d(\PWMB/n23 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[0]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b1  (
    .clk(clk100m),
    .d(\PWMB/n23 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[1]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b10  (
    .clk(clk100m),
    .d(\PWMB/n23 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[10]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b11  (
    .clk(clk100m),
    .d(\PWMB/n23 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[11]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b12  (
    .clk(clk100m),
    .d(\PWMB/n23 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[12]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b13  (
    .clk(clk100m),
    .d(\PWMB/n23 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[13]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b14  (
    .clk(clk100m),
    .d(\PWMB/n23 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[14]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b15  (
    .clk(clk100m),
    .d(\PWMB/n23 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[15]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b16  (
    .clk(clk100m),
    .d(\PWMB/n23 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[16]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b17  (
    .clk(clk100m),
    .d(\PWMB/n23 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[17]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b18  (
    .clk(clk100m),
    .d(\PWMB/n23 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[18]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b19  (
    .clk(clk100m),
    .d(\PWMB/n23 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[19]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b2  (
    .clk(clk100m),
    .d(\PWMB/n23 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[2]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b20  (
    .clk(clk100m),
    .d(\PWMB/n23 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[20]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b21  (
    .clk(clk100m),
    .d(\PWMB/n23 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[21]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b22  (
    .clk(clk100m),
    .d(\PWMB/n23 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[22]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b23  (
    .clk(clk100m),
    .d(\PWMB/n23 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[23]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b24  (
    .clk(clk100m),
    .d(\PWMB/n23 [24]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[24]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b25  (
    .clk(clk100m),
    .d(\PWMB/n23 [25]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[25]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b26  (
    .clk(clk100m),
    .d(\PWMB/n23 [26]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[26]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b27  (
    .clk(clk100m),
    .d(\PWMB/n23 [27]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[27]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b28  (
    .clk(clk100m),
    .d(\PWMB/n23 [28]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[28]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b29  (
    .clk(clk100m),
    .d(\PWMB/n23 [29]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[29]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b3  (
    .clk(clk100m),
    .d(\PWMB/n23 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[3]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b30  (
    .clk(clk100m),
    .d(\PWMB/n23 [30]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[30]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b31  (
    .clk(clk100m),
    .d(\PWMB/n23 [31]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[31]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b4  (
    .clk(clk100m),
    .d(\PWMB/n23 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[4]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b5  (
    .clk(clk100m),
    .d(\PWMB/n23 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[5]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b6  (
    .clk(clk100m),
    .d(\PWMB/n23 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[6]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b7  (
    .clk(clk100m),
    .d(\PWMB/n23 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[7]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b8  (
    .clk(clk100m),
    .d(\PWMB/n23 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[8]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b9  (
    .clk(clk100m),
    .d(\PWMB/n23 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[9]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg3_b0  (
    .clk(clk100m),
    .d(\PWMB/n31 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[0]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b1  (
    .clk(clk100m),
    .d(\PWMB/n31 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[1]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b10  (
    .clk(clk100m),
    .d(\PWMB/n31 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[10]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b11  (
    .clk(clk100m),
    .d(\PWMB/n31 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[11]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b12  (
    .clk(clk100m),
    .d(\PWMB/n31 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[12]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b13  (
    .clk(clk100m),
    .d(\PWMB/n31 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[13]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b14  (
    .clk(clk100m),
    .d(\PWMB/n31 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[14]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b15  (
    .clk(clk100m),
    .d(\PWMB/n31 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[15]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b16  (
    .clk(clk100m),
    .d(\PWMB/n31 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[16]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b17  (
    .clk(clk100m),
    .d(\PWMB/n31 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[17]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b18  (
    .clk(clk100m),
    .d(\PWMB/n31 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[18]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b19  (
    .clk(clk100m),
    .d(\PWMB/n31 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[19]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b2  (
    .clk(clk100m),
    .d(\PWMB/n31 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[2]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b20  (
    .clk(clk100m),
    .d(\PWMB/n31 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[20]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b21  (
    .clk(clk100m),
    .d(\PWMB/n31 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[21]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b22  (
    .clk(clk100m),
    .d(\PWMB/n31 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[22]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b23  (
    .clk(clk100m),
    .d(\PWMB/n31 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[23]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b3  (
    .clk(clk100m),
    .d(\PWMB/n31 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[3]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b4  (
    .clk(clk100m),
    .d(\PWMB/n31 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[4]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b5  (
    .clk(clk100m),
    .d(\PWMB/n31 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[5]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b6  (
    .clk(clk100m),
    .d(\PWMB/n31 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[6]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b7  (
    .clk(clk100m),
    .d(\PWMB/n31 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[7]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b8  (
    .clk(clk100m),
    .d(\PWMB/n31 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[8]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b9  (
    .clk(clk100m),
    .d(\PWMB/n31 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[9]_keep ));  // src/OnePWM.v(58)
  reg_ar_ss_w1 \PWMB/stopreq_reg  (
    .clk(clk100m),
    .d(\PWMB/n1 ),
    .en(1'b1),
    .reset(1'b0),
    .set(pwm_start_stop[11]),
    .q(\PWMB/stopreq_keep ));  // src/OnePWM.v(15)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub0/u0  (
    .a(\PWMB/FreCnt [0]),
    .b(1'b1),
    .c(\PWMB/sub0/c0 ),
    .o({\PWMB/sub0/c1 ,\PWMB/n12 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub0/u1  (
    .a(\PWMB/FreCnt [1]),
    .b(1'b0),
    .c(\PWMB/sub0/c1 ),
    .o({\PWMB/sub0/c2 ,\PWMB/n12 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub0/u10  (
    .a(\PWMB/FreCnt [10]),
    .b(1'b0),
    .c(\PWMB/sub0/c10 ),
    .o({\PWMB/sub0/c11 ,\PWMB/n12 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub0/u11  (
    .a(\PWMB/FreCnt [11]),
    .b(1'b0),
    .c(\PWMB/sub0/c11 ),
    .o({\PWMB/sub0/c12 ,\PWMB/n12 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub0/u12  (
    .a(\PWMB/FreCnt [12]),
    .b(1'b0),
    .c(\PWMB/sub0/c12 ),
    .o({\PWMB/sub0/c13 ,\PWMB/n12 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub0/u13  (
    .a(\PWMB/FreCnt [13]),
    .b(1'b0),
    .c(\PWMB/sub0/c13 ),
    .o({\PWMB/sub0/c14 ,\PWMB/n12 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub0/u14  (
    .a(\PWMB/FreCnt [14]),
    .b(1'b0),
    .c(\PWMB/sub0/c14 ),
    .o({\PWMB/sub0/c15 ,\PWMB/n12 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub0/u15  (
    .a(\PWMB/FreCnt [15]),
    .b(1'b0),
    .c(\PWMB/sub0/c15 ),
    .o({\PWMB/sub0/c16 ,\PWMB/n12 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub0/u16  (
    .a(\PWMB/FreCnt [16]),
    .b(1'b0),
    .c(\PWMB/sub0/c16 ),
    .o({\PWMB/sub0/c17 ,\PWMB/n12 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub0/u17  (
    .a(\PWMB/FreCnt [17]),
    .b(1'b0),
    .c(\PWMB/sub0/c17 ),
    .o({\PWMB/sub0/c18 ,\PWMB/n12 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub0/u18  (
    .a(\PWMB/FreCnt [18]),
    .b(1'b0),
    .c(\PWMB/sub0/c18 ),
    .o({\PWMB/sub0/c19 ,\PWMB/n12 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub0/u19  (
    .a(\PWMB/FreCnt [19]),
    .b(1'b0),
    .c(\PWMB/sub0/c19 ),
    .o({\PWMB/sub0/c20 ,\PWMB/n12 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub0/u2  (
    .a(\PWMB/FreCnt [2]),
    .b(1'b0),
    .c(\PWMB/sub0/c2 ),
    .o({\PWMB/sub0/c3 ,\PWMB/n12 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub0/u20  (
    .a(\PWMB/FreCnt [20]),
    .b(1'b0),
    .c(\PWMB/sub0/c20 ),
    .o({\PWMB/sub0/c21 ,\PWMB/n12 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub0/u21  (
    .a(\PWMB/FreCnt [21]),
    .b(1'b0),
    .c(\PWMB/sub0/c21 ),
    .o({\PWMB/sub0/c22 ,\PWMB/n12 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub0/u22  (
    .a(\PWMB/FreCnt [22]),
    .b(1'b0),
    .c(\PWMB/sub0/c22 ),
    .o({\PWMB/sub0/c23 ,\PWMB/n12 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub0/u23  (
    .a(\PWMB/FreCnt [23]),
    .b(1'b0),
    .c(\PWMB/sub0/c23 ),
    .o({\PWMB/sub0/c24 ,\PWMB/n12 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub0/u24  (
    .a(\PWMB/FreCnt [24]),
    .b(1'b0),
    .c(\PWMB/sub0/c24 ),
    .o({\PWMB/sub0/c25 ,\PWMB/n12 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub0/u25  (
    .a(\PWMB/FreCnt [25]),
    .b(1'b0),
    .c(\PWMB/sub0/c25 ),
    .o({\PWMB/sub0/c26 ,\PWMB/n12 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub0/u26  (
    .a(\PWMB/FreCnt [26]),
    .b(1'b0),
    .c(\PWMB/sub0/c26 ),
    .o({open_n88,\PWMB/n12 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub0/u3  (
    .a(\PWMB/FreCnt [3]),
    .b(1'b0),
    .c(\PWMB/sub0/c3 ),
    .o({\PWMB/sub0/c4 ,\PWMB/n12 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub0/u4  (
    .a(\PWMB/FreCnt [4]),
    .b(1'b0),
    .c(\PWMB/sub0/c4 ),
    .o({\PWMB/sub0/c5 ,\PWMB/n12 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub0/u5  (
    .a(\PWMB/FreCnt [5]),
    .b(1'b0),
    .c(\PWMB/sub0/c5 ),
    .o({\PWMB/sub0/c6 ,\PWMB/n12 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub0/u6  (
    .a(\PWMB/FreCnt [6]),
    .b(1'b0),
    .c(\PWMB/sub0/c6 ),
    .o({\PWMB/sub0/c7 ,\PWMB/n12 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub0/u7  (
    .a(\PWMB/FreCnt [7]),
    .b(1'b0),
    .c(\PWMB/sub0/c7 ),
    .o({\PWMB/sub0/c8 ,\PWMB/n12 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub0/u8  (
    .a(\PWMB/FreCnt [8]),
    .b(1'b0),
    .c(\PWMB/sub0/c8 ),
    .o({\PWMB/sub0/c9 ,\PWMB/n12 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub0/u9  (
    .a(\PWMB/FreCnt [9]),
    .b(1'b0),
    .c(\PWMB/sub0/c9 ),
    .o({\PWMB/sub0/c10 ,\PWMB/n12 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \PWMB/sub0/ucin  (
    .a(1'b0),
    .o({\PWMB/sub0/c0 ,open_n91}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub1/u0  (
    .a(pnumcntB[0]),
    .b(1'b1),
    .c(\PWMB/sub1/c0 ),
    .o({\PWMB/sub1/c1 ,\PWMB/n26 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub1/u1  (
    .a(pnumcntB[1]),
    .b(1'b0),
    .c(\PWMB/sub1/c1 ),
    .o({\PWMB/sub1/c2 ,\PWMB/n26 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub1/u10  (
    .a(pnumcntB[10]),
    .b(1'b0),
    .c(\PWMB/sub1/c10 ),
    .o({\PWMB/sub1/c11 ,\PWMB/n26 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub1/u11  (
    .a(pnumcntB[11]),
    .b(1'b0),
    .c(\PWMB/sub1/c11 ),
    .o({\PWMB/sub1/c12 ,\PWMB/n26 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub1/u12  (
    .a(pnumcntB[12]),
    .b(1'b0),
    .c(\PWMB/sub1/c12 ),
    .o({\PWMB/sub1/c13 ,\PWMB/n26 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub1/u13  (
    .a(pnumcntB[13]),
    .b(1'b0),
    .c(\PWMB/sub1/c13 ),
    .o({\PWMB/sub1/c14 ,\PWMB/n26 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub1/u14  (
    .a(pnumcntB[14]),
    .b(1'b0),
    .c(\PWMB/sub1/c14 ),
    .o({\PWMB/sub1/c15 ,\PWMB/n26 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub1/u15  (
    .a(pnumcntB[15]),
    .b(1'b0),
    .c(\PWMB/sub1/c15 ),
    .o({\PWMB/sub1/c16 ,\PWMB/n26 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub1/u16  (
    .a(pnumcntB[16]),
    .b(1'b0),
    .c(\PWMB/sub1/c16 ),
    .o({\PWMB/sub1/c17 ,\PWMB/n26 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub1/u17  (
    .a(pnumcntB[17]),
    .b(1'b0),
    .c(\PWMB/sub1/c17 ),
    .o({\PWMB/sub1/c18 ,\PWMB/n26 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub1/u18  (
    .a(pnumcntB[18]),
    .b(1'b0),
    .c(\PWMB/sub1/c18 ),
    .o({\PWMB/sub1/c19 ,\PWMB/n26 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub1/u19  (
    .a(pnumcntB[19]),
    .b(1'b0),
    .c(\PWMB/sub1/c19 ),
    .o({\PWMB/sub1/c20 ,\PWMB/n26 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub1/u2  (
    .a(pnumcntB[2]),
    .b(1'b0),
    .c(\PWMB/sub1/c2 ),
    .o({\PWMB/sub1/c3 ,\PWMB/n26 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub1/u20  (
    .a(pnumcntB[20]),
    .b(1'b0),
    .c(\PWMB/sub1/c20 ),
    .o({\PWMB/sub1/c21 ,\PWMB/n26 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub1/u21  (
    .a(pnumcntB[21]),
    .b(1'b0),
    .c(\PWMB/sub1/c21 ),
    .o({\PWMB/sub1/c22 ,\PWMB/n26 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub1/u22  (
    .a(pnumcntB[22]),
    .b(1'b0),
    .c(\PWMB/sub1/c22 ),
    .o({\PWMB/sub1/c23 ,\PWMB/n26 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub1/u23  (
    .a(pnumcntB[23]),
    .b(1'b0),
    .c(\PWMB/sub1/c23 ),
    .o({open_n92,\PWMB/n26 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub1/u3  (
    .a(pnumcntB[3]),
    .b(1'b0),
    .c(\PWMB/sub1/c3 ),
    .o({\PWMB/sub1/c4 ,\PWMB/n26 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub1/u4  (
    .a(pnumcntB[4]),
    .b(1'b0),
    .c(\PWMB/sub1/c4 ),
    .o({\PWMB/sub1/c5 ,\PWMB/n26 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub1/u5  (
    .a(pnumcntB[5]),
    .b(1'b0),
    .c(\PWMB/sub1/c5 ),
    .o({\PWMB/sub1/c6 ,\PWMB/n26 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub1/u6  (
    .a(pnumcntB[6]),
    .b(1'b0),
    .c(\PWMB/sub1/c6 ),
    .o({\PWMB/sub1/c7 ,\PWMB/n26 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub1/u7  (
    .a(pnumcntB[7]),
    .b(1'b0),
    .c(\PWMB/sub1/c7 ),
    .o({\PWMB/sub1/c8 ,\PWMB/n26 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub1/u8  (
    .a(pnumcntB[8]),
    .b(1'b0),
    .c(\PWMB/sub1/c8 ),
    .o({\PWMB/sub1/c9 ,\PWMB/n26 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMB/sub1/u9  (
    .a(pnumcntB[9]),
    .b(1'b0),
    .c(\PWMB/sub1/c9 ),
    .o({\PWMB/sub1/c10 ,\PWMB/n26 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \PWMB/sub1/ucin  (
    .a(1'b0),
    .o({\PWMB/sub1/c0 ,open_n95}));
  reg_ar_as_w1 \PWMC/State_reg  (
    .clk(clk100m),
    .d(\PWMC/n10 ),
    .en(1'b1),
    .reset(~rstn),
    .set(1'b0),
    .q(pwm_state_read[12]));  // src/OnePWM.v(26)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[0]  (
    .i(\PWMC/RemaTxNum[0]_keep ),
    .o(pnumcntC[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[10]  (
    .i(\PWMC/RemaTxNum[10]_keep ),
    .o(pnumcntC[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[11]  (
    .i(\PWMC/RemaTxNum[11]_keep ),
    .o(pnumcntC[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[12]  (
    .i(\PWMC/RemaTxNum[12]_keep ),
    .o(pnumcntC[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[13]  (
    .i(\PWMC/RemaTxNum[13]_keep ),
    .o(pnumcntC[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[14]  (
    .i(\PWMC/RemaTxNum[14]_keep ),
    .o(pnumcntC[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[15]  (
    .i(\PWMC/RemaTxNum[15]_keep ),
    .o(pnumcntC[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[16]  (
    .i(\PWMC/RemaTxNum[16]_keep ),
    .o(pnumcntC[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[17]  (
    .i(\PWMC/RemaTxNum[17]_keep ),
    .o(pnumcntC[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[18]  (
    .i(\PWMC/RemaTxNum[18]_keep ),
    .o(pnumcntC[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[19]  (
    .i(\PWMC/RemaTxNum[19]_keep ),
    .o(pnumcntC[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[1]  (
    .i(\PWMC/RemaTxNum[1]_keep ),
    .o(pnumcntC[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[20]  (
    .i(\PWMC/RemaTxNum[20]_keep ),
    .o(pnumcntC[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[21]  (
    .i(\PWMC/RemaTxNum[21]_keep ),
    .o(pnumcntC[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[22]  (
    .i(\PWMC/RemaTxNum[22]_keep ),
    .o(pnumcntC[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[23]  (
    .i(\PWMC/RemaTxNum[23]_keep ),
    .o(pnumcntC[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[2]  (
    .i(\PWMC/RemaTxNum[2]_keep ),
    .o(pnumcntC[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[3]  (
    .i(\PWMC/RemaTxNum[3]_keep ),
    .o(pnumcntC[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[4]  (
    .i(\PWMC/RemaTxNum[4]_keep ),
    .o(pnumcntC[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[5]  (
    .i(\PWMC/RemaTxNum[5]_keep ),
    .o(pnumcntC[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[6]  (
    .i(\PWMC/RemaTxNum[6]_keep ),
    .o(pnumcntC[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[7]  (
    .i(\PWMC/RemaTxNum[7]_keep ),
    .o(pnumcntC[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[8]  (
    .i(\PWMC/RemaTxNum[8]_keep ),
    .o(pnumcntC[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[9]  (
    .i(\PWMC/RemaTxNum[9]_keep ),
    .o(pnumcntC[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_dir  (
    .i(\PWMC/dir_keep ),
    .o(dir_pad[12]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[0]  (
    .i(\PWMC/pnumr[0]_keep ),
    .o(\PWMC/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[10]  (
    .i(\PWMC/pnumr[10]_keep ),
    .o(\PWMC/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[11]  (
    .i(\PWMC/pnumr[11]_keep ),
    .o(\PWMC/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[12]  (
    .i(\PWMC/pnumr[12]_keep ),
    .o(\PWMC/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[13]  (
    .i(\PWMC/pnumr[13]_keep ),
    .o(\PWMC/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[14]  (
    .i(\PWMC/pnumr[14]_keep ),
    .o(\PWMC/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[15]  (
    .i(\PWMC/pnumr[15]_keep ),
    .o(\PWMC/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[16]  (
    .i(\PWMC/pnumr[16]_keep ),
    .o(\PWMC/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[17]  (
    .i(\PWMC/pnumr[17]_keep ),
    .o(\PWMC/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[18]  (
    .i(\PWMC/pnumr[18]_keep ),
    .o(\PWMC/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[19]  (
    .i(\PWMC/pnumr[19]_keep ),
    .o(\PWMC/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[1]  (
    .i(\PWMC/pnumr[1]_keep ),
    .o(\PWMC/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[20]  (
    .i(\PWMC/pnumr[20]_keep ),
    .o(\PWMC/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[21]  (
    .i(\PWMC/pnumr[21]_keep ),
    .o(\PWMC/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[22]  (
    .i(\PWMC/pnumr[22]_keep ),
    .o(\PWMC/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[23]  (
    .i(\PWMC/pnumr[23]_keep ),
    .o(\PWMC/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[24]  (
    .i(\PWMC/pnumr[24]_keep ),
    .o(\PWMC/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[25]  (
    .i(\PWMC/pnumr[25]_keep ),
    .o(\PWMC/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[26]  (
    .i(\PWMC/pnumr[26]_keep ),
    .o(\PWMC/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[27]  (
    .i(\PWMC/pnumr[27]_keep ),
    .o(\PWMC/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[28]  (
    .i(\PWMC/pnumr[28]_keep ),
    .o(\PWMC/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[29]  (
    .i(\PWMC/pnumr[29]_keep ),
    .o(\PWMC/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[2]  (
    .i(\PWMC/pnumr[2]_keep ),
    .o(\PWMC/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[30]  (
    .i(\PWMC/pnumr[30]_keep ),
    .o(\PWMC/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[31]  (
    .i(\PWMC/pnumr[31]_keep ),
    .o(\PWMC/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[3]  (
    .i(\PWMC/pnumr[3]_keep ),
    .o(\PWMC/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[4]  (
    .i(\PWMC/pnumr[4]_keep ),
    .o(\PWMC/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[5]  (
    .i(\PWMC/pnumr[5]_keep ),
    .o(\PWMC/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[6]  (
    .i(\PWMC/pnumr[6]_keep ),
    .o(\PWMC/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[7]  (
    .i(\PWMC/pnumr[7]_keep ),
    .o(\PWMC/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[8]  (
    .i(\PWMC/pnumr[8]_keep ),
    .o(\PWMC/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[9]  (
    .i(\PWMC/pnumr[9]_keep ),
    .o(\PWMC/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pwm  (
    .i(\PWMC/pwm_keep ),
    .o(pwm_pad[12]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_stopreq  (
    .i(\PWMC/stopreq_keep ),
    .o(\PWMC/stopreq ));  // src/OnePWM.v(14)
  reg_ar_as_w1 \PWMC/dir_reg  (
    .clk(clk100m),
    .d(\PWMC/n32 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/dir_keep ));  // src/OnePWM.v(58)
  reg_sr_as_w1 \PWMC/pwm_reg  (
    .clk(clk100m),
    .d(\pwm[12]_d ),
    .en(1'b1),
    .reset(~\PWMC/u14_sel_is_1_o ),
    .set(1'b0),
    .q(\PWMC/pwm_keep ));  // src/OnePWM.v(45)
  reg_sr_as_w1 \PWMC/reg0_b0  (
    .clk(clk100m),
    .d(\PWMC/n13 [0]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [0]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b1  (
    .clk(clk100m),
    .d(\PWMC/n13 [1]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [1]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b10  (
    .clk(clk100m),
    .d(\PWMC/n13 [10]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [10]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b11  (
    .clk(clk100m),
    .d(\PWMC/n13 [11]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [11]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b12  (
    .clk(clk100m),
    .d(\PWMC/n13 [12]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [12]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b13  (
    .clk(clk100m),
    .d(\PWMC/n13 [13]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [13]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b14  (
    .clk(clk100m),
    .d(\PWMC/n13 [14]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [14]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b15  (
    .clk(clk100m),
    .d(\PWMC/n13 [15]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [15]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b16  (
    .clk(clk100m),
    .d(\PWMC/n13 [16]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [16]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b17  (
    .clk(clk100m),
    .d(\PWMC/n13 [17]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [17]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b18  (
    .clk(clk100m),
    .d(\PWMC/n13 [18]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [18]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b19  (
    .clk(clk100m),
    .d(\PWMC/n13 [19]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [19]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b2  (
    .clk(clk100m),
    .d(\PWMC/n13 [2]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [2]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b20  (
    .clk(clk100m),
    .d(\PWMC/n13 [20]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [20]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b21  (
    .clk(clk100m),
    .d(\PWMC/n13 [21]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [21]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b22  (
    .clk(clk100m),
    .d(\PWMC/n13 [22]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [22]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b23  (
    .clk(clk100m),
    .d(\PWMC/n13 [23]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [23]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b24  (
    .clk(clk100m),
    .d(\PWMC/n13 [24]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [24]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b25  (
    .clk(clk100m),
    .d(\PWMC/n13 [25]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [25]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b26  (
    .clk(clk100m),
    .d(\PWMC/n13 [26]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [26]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b3  (
    .clk(clk100m),
    .d(\PWMC/n13 [3]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [3]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b4  (
    .clk(clk100m),
    .d(\PWMC/n13 [4]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [4]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b5  (
    .clk(clk100m),
    .d(\PWMC/n13 [5]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [5]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b6  (
    .clk(clk100m),
    .d(\PWMC/n13 [6]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [6]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b7  (
    .clk(clk100m),
    .d(\PWMC/n13 [7]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [7]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b8  (
    .clk(clk100m),
    .d(\PWMC/n13 [8]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [8]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b9  (
    .clk(clk100m),
    .d(\PWMC/n13 [9]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b0  (
    .clk(clk100m),
    .d(freqC[0]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [0]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b1  (
    .clk(clk100m),
    .d(freqC[1]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [1]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b10  (
    .clk(clk100m),
    .d(freqC[10]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [10]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b11  (
    .clk(clk100m),
    .d(freqC[11]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [11]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b12  (
    .clk(clk100m),
    .d(freqC[12]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [12]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b13  (
    .clk(clk100m),
    .d(freqC[13]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [13]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b14  (
    .clk(clk100m),
    .d(freqC[14]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [14]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b15  (
    .clk(clk100m),
    .d(freqC[15]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [15]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b16  (
    .clk(clk100m),
    .d(freqC[16]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [16]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b17  (
    .clk(clk100m),
    .d(freqC[17]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [17]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b18  (
    .clk(clk100m),
    .d(freqC[18]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [18]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b19  (
    .clk(clk100m),
    .d(freqC[19]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [19]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b2  (
    .clk(clk100m),
    .d(freqC[2]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [2]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b20  (
    .clk(clk100m),
    .d(freqC[20]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [20]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b21  (
    .clk(clk100m),
    .d(freqC[21]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [21]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b22  (
    .clk(clk100m),
    .d(freqC[22]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [22]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b23  (
    .clk(clk100m),
    .d(freqC[23]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [23]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b24  (
    .clk(clk100m),
    .d(freqC[24]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [24]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b25  (
    .clk(clk100m),
    .d(freqC[25]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [25]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b26  (
    .clk(clk100m),
    .d(freqC[26]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [26]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b3  (
    .clk(clk100m),
    .d(freqC[3]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [3]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b4  (
    .clk(clk100m),
    .d(freqC[4]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [4]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b5  (
    .clk(clk100m),
    .d(freqC[5]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [5]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b6  (
    .clk(clk100m),
    .d(freqC[6]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [6]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b7  (
    .clk(clk100m),
    .d(freqC[7]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [7]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b8  (
    .clk(clk100m),
    .d(freqC[8]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [8]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b9  (
    .clk(clk100m),
    .d(freqC[9]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg2_b0  (
    .clk(clk100m),
    .d(\PWMC/n23 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[0]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b1  (
    .clk(clk100m),
    .d(\PWMC/n23 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[1]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b10  (
    .clk(clk100m),
    .d(\PWMC/n23 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[10]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b11  (
    .clk(clk100m),
    .d(\PWMC/n23 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[11]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b12  (
    .clk(clk100m),
    .d(\PWMC/n23 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[12]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b13  (
    .clk(clk100m),
    .d(\PWMC/n23 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[13]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b14  (
    .clk(clk100m),
    .d(\PWMC/n23 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[14]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b15  (
    .clk(clk100m),
    .d(\PWMC/n23 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[15]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b16  (
    .clk(clk100m),
    .d(\PWMC/n23 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[16]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b17  (
    .clk(clk100m),
    .d(\PWMC/n23 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[17]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b18  (
    .clk(clk100m),
    .d(\PWMC/n23 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[18]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b19  (
    .clk(clk100m),
    .d(\PWMC/n23 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[19]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b2  (
    .clk(clk100m),
    .d(\PWMC/n23 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[2]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b20  (
    .clk(clk100m),
    .d(\PWMC/n23 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[20]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b21  (
    .clk(clk100m),
    .d(\PWMC/n23 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[21]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b22  (
    .clk(clk100m),
    .d(\PWMC/n23 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[22]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b23  (
    .clk(clk100m),
    .d(\PWMC/n23 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[23]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b24  (
    .clk(clk100m),
    .d(\PWMC/n23 [24]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[24]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b25  (
    .clk(clk100m),
    .d(\PWMC/n23 [25]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[25]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b26  (
    .clk(clk100m),
    .d(\PWMC/n23 [26]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[26]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b27  (
    .clk(clk100m),
    .d(\PWMC/n23 [27]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[27]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b28  (
    .clk(clk100m),
    .d(\PWMC/n23 [28]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[28]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b29  (
    .clk(clk100m),
    .d(\PWMC/n23 [29]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[29]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b3  (
    .clk(clk100m),
    .d(\PWMC/n23 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[3]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b30  (
    .clk(clk100m),
    .d(\PWMC/n23 [30]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[30]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b31  (
    .clk(clk100m),
    .d(\PWMC/n23 [31]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[31]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b4  (
    .clk(clk100m),
    .d(\PWMC/n23 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[4]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b5  (
    .clk(clk100m),
    .d(\PWMC/n23 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[5]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b6  (
    .clk(clk100m),
    .d(\PWMC/n23 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[6]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b7  (
    .clk(clk100m),
    .d(\PWMC/n23 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[7]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b8  (
    .clk(clk100m),
    .d(\PWMC/n23 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[8]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b9  (
    .clk(clk100m),
    .d(\PWMC/n23 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[9]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg3_b0  (
    .clk(clk100m),
    .d(\PWMC/n31 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[0]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b1  (
    .clk(clk100m),
    .d(\PWMC/n31 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[1]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b10  (
    .clk(clk100m),
    .d(\PWMC/n31 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[10]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b11  (
    .clk(clk100m),
    .d(\PWMC/n31 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[11]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b12  (
    .clk(clk100m),
    .d(\PWMC/n31 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[12]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b13  (
    .clk(clk100m),
    .d(\PWMC/n31 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[13]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b14  (
    .clk(clk100m),
    .d(\PWMC/n31 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[14]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b15  (
    .clk(clk100m),
    .d(\PWMC/n31 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[15]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b16  (
    .clk(clk100m),
    .d(\PWMC/n31 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[16]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b17  (
    .clk(clk100m),
    .d(\PWMC/n31 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[17]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b18  (
    .clk(clk100m),
    .d(\PWMC/n31 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[18]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b19  (
    .clk(clk100m),
    .d(\PWMC/n31 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[19]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b2  (
    .clk(clk100m),
    .d(\PWMC/n31 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[2]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b20  (
    .clk(clk100m),
    .d(\PWMC/n31 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[20]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b21  (
    .clk(clk100m),
    .d(\PWMC/n31 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[21]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b22  (
    .clk(clk100m),
    .d(\PWMC/n31 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[22]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b23  (
    .clk(clk100m),
    .d(\PWMC/n31 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[23]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b3  (
    .clk(clk100m),
    .d(\PWMC/n31 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[3]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b4  (
    .clk(clk100m),
    .d(\PWMC/n31 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[4]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b5  (
    .clk(clk100m),
    .d(\PWMC/n31 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[5]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b6  (
    .clk(clk100m),
    .d(\PWMC/n31 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[6]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b7  (
    .clk(clk100m),
    .d(\PWMC/n31 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[7]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b8  (
    .clk(clk100m),
    .d(\PWMC/n31 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[8]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b9  (
    .clk(clk100m),
    .d(\PWMC/n31 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[9]_keep ));  // src/OnePWM.v(58)
  reg_ar_ss_w1 \PWMC/stopreq_reg  (
    .clk(clk100m),
    .d(\PWMC/n1 ),
    .en(1'b1),
    .reset(1'b0),
    .set(pwm_start_stop[12]),
    .q(\PWMC/stopreq_keep ));  // src/OnePWM.v(15)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub0/u0  (
    .a(\PWMC/FreCnt [0]),
    .b(1'b1),
    .c(\PWMC/sub0/c0 ),
    .o({\PWMC/sub0/c1 ,\PWMC/n12 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub0/u1  (
    .a(\PWMC/FreCnt [1]),
    .b(1'b0),
    .c(\PWMC/sub0/c1 ),
    .o({\PWMC/sub0/c2 ,\PWMC/n12 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub0/u10  (
    .a(\PWMC/FreCnt [10]),
    .b(1'b0),
    .c(\PWMC/sub0/c10 ),
    .o({\PWMC/sub0/c11 ,\PWMC/n12 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub0/u11  (
    .a(\PWMC/FreCnt [11]),
    .b(1'b0),
    .c(\PWMC/sub0/c11 ),
    .o({\PWMC/sub0/c12 ,\PWMC/n12 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub0/u12  (
    .a(\PWMC/FreCnt [12]),
    .b(1'b0),
    .c(\PWMC/sub0/c12 ),
    .o({\PWMC/sub0/c13 ,\PWMC/n12 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub0/u13  (
    .a(\PWMC/FreCnt [13]),
    .b(1'b0),
    .c(\PWMC/sub0/c13 ),
    .o({\PWMC/sub0/c14 ,\PWMC/n12 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub0/u14  (
    .a(\PWMC/FreCnt [14]),
    .b(1'b0),
    .c(\PWMC/sub0/c14 ),
    .o({\PWMC/sub0/c15 ,\PWMC/n12 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub0/u15  (
    .a(\PWMC/FreCnt [15]),
    .b(1'b0),
    .c(\PWMC/sub0/c15 ),
    .o({\PWMC/sub0/c16 ,\PWMC/n12 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub0/u16  (
    .a(\PWMC/FreCnt [16]),
    .b(1'b0),
    .c(\PWMC/sub0/c16 ),
    .o({\PWMC/sub0/c17 ,\PWMC/n12 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub0/u17  (
    .a(\PWMC/FreCnt [17]),
    .b(1'b0),
    .c(\PWMC/sub0/c17 ),
    .o({\PWMC/sub0/c18 ,\PWMC/n12 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub0/u18  (
    .a(\PWMC/FreCnt [18]),
    .b(1'b0),
    .c(\PWMC/sub0/c18 ),
    .o({\PWMC/sub0/c19 ,\PWMC/n12 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub0/u19  (
    .a(\PWMC/FreCnt [19]),
    .b(1'b0),
    .c(\PWMC/sub0/c19 ),
    .o({\PWMC/sub0/c20 ,\PWMC/n12 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub0/u2  (
    .a(\PWMC/FreCnt [2]),
    .b(1'b0),
    .c(\PWMC/sub0/c2 ),
    .o({\PWMC/sub0/c3 ,\PWMC/n12 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub0/u20  (
    .a(\PWMC/FreCnt [20]),
    .b(1'b0),
    .c(\PWMC/sub0/c20 ),
    .o({\PWMC/sub0/c21 ,\PWMC/n12 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub0/u21  (
    .a(\PWMC/FreCnt [21]),
    .b(1'b0),
    .c(\PWMC/sub0/c21 ),
    .o({\PWMC/sub0/c22 ,\PWMC/n12 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub0/u22  (
    .a(\PWMC/FreCnt [22]),
    .b(1'b0),
    .c(\PWMC/sub0/c22 ),
    .o({\PWMC/sub0/c23 ,\PWMC/n12 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub0/u23  (
    .a(\PWMC/FreCnt [23]),
    .b(1'b0),
    .c(\PWMC/sub0/c23 ),
    .o({\PWMC/sub0/c24 ,\PWMC/n12 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub0/u24  (
    .a(\PWMC/FreCnt [24]),
    .b(1'b0),
    .c(\PWMC/sub0/c24 ),
    .o({\PWMC/sub0/c25 ,\PWMC/n12 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub0/u25  (
    .a(\PWMC/FreCnt [25]),
    .b(1'b0),
    .c(\PWMC/sub0/c25 ),
    .o({\PWMC/sub0/c26 ,\PWMC/n12 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub0/u26  (
    .a(\PWMC/FreCnt [26]),
    .b(1'b0),
    .c(\PWMC/sub0/c26 ),
    .o({open_n96,\PWMC/n12 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub0/u3  (
    .a(\PWMC/FreCnt [3]),
    .b(1'b0),
    .c(\PWMC/sub0/c3 ),
    .o({\PWMC/sub0/c4 ,\PWMC/n12 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub0/u4  (
    .a(\PWMC/FreCnt [4]),
    .b(1'b0),
    .c(\PWMC/sub0/c4 ),
    .o({\PWMC/sub0/c5 ,\PWMC/n12 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub0/u5  (
    .a(\PWMC/FreCnt [5]),
    .b(1'b0),
    .c(\PWMC/sub0/c5 ),
    .o({\PWMC/sub0/c6 ,\PWMC/n12 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub0/u6  (
    .a(\PWMC/FreCnt [6]),
    .b(1'b0),
    .c(\PWMC/sub0/c6 ),
    .o({\PWMC/sub0/c7 ,\PWMC/n12 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub0/u7  (
    .a(\PWMC/FreCnt [7]),
    .b(1'b0),
    .c(\PWMC/sub0/c7 ),
    .o({\PWMC/sub0/c8 ,\PWMC/n12 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub0/u8  (
    .a(\PWMC/FreCnt [8]),
    .b(1'b0),
    .c(\PWMC/sub0/c8 ),
    .o({\PWMC/sub0/c9 ,\PWMC/n12 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub0/u9  (
    .a(\PWMC/FreCnt [9]),
    .b(1'b0),
    .c(\PWMC/sub0/c9 ),
    .o({\PWMC/sub0/c10 ,\PWMC/n12 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \PWMC/sub0/ucin  (
    .a(1'b0),
    .o({\PWMC/sub0/c0 ,open_n99}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub1/u0  (
    .a(pnumcntC[0]),
    .b(1'b1),
    .c(\PWMC/sub1/c0 ),
    .o({\PWMC/sub1/c1 ,\PWMC/n26 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub1/u1  (
    .a(pnumcntC[1]),
    .b(1'b0),
    .c(\PWMC/sub1/c1 ),
    .o({\PWMC/sub1/c2 ,\PWMC/n26 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub1/u10  (
    .a(pnumcntC[10]),
    .b(1'b0),
    .c(\PWMC/sub1/c10 ),
    .o({\PWMC/sub1/c11 ,\PWMC/n26 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub1/u11  (
    .a(pnumcntC[11]),
    .b(1'b0),
    .c(\PWMC/sub1/c11 ),
    .o({\PWMC/sub1/c12 ,\PWMC/n26 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub1/u12  (
    .a(pnumcntC[12]),
    .b(1'b0),
    .c(\PWMC/sub1/c12 ),
    .o({\PWMC/sub1/c13 ,\PWMC/n26 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub1/u13  (
    .a(pnumcntC[13]),
    .b(1'b0),
    .c(\PWMC/sub1/c13 ),
    .o({\PWMC/sub1/c14 ,\PWMC/n26 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub1/u14  (
    .a(pnumcntC[14]),
    .b(1'b0),
    .c(\PWMC/sub1/c14 ),
    .o({\PWMC/sub1/c15 ,\PWMC/n26 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub1/u15  (
    .a(pnumcntC[15]),
    .b(1'b0),
    .c(\PWMC/sub1/c15 ),
    .o({\PWMC/sub1/c16 ,\PWMC/n26 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub1/u16  (
    .a(pnumcntC[16]),
    .b(1'b0),
    .c(\PWMC/sub1/c16 ),
    .o({\PWMC/sub1/c17 ,\PWMC/n26 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub1/u17  (
    .a(pnumcntC[17]),
    .b(1'b0),
    .c(\PWMC/sub1/c17 ),
    .o({\PWMC/sub1/c18 ,\PWMC/n26 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub1/u18  (
    .a(pnumcntC[18]),
    .b(1'b0),
    .c(\PWMC/sub1/c18 ),
    .o({\PWMC/sub1/c19 ,\PWMC/n26 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub1/u19  (
    .a(pnumcntC[19]),
    .b(1'b0),
    .c(\PWMC/sub1/c19 ),
    .o({\PWMC/sub1/c20 ,\PWMC/n26 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub1/u2  (
    .a(pnumcntC[2]),
    .b(1'b0),
    .c(\PWMC/sub1/c2 ),
    .o({\PWMC/sub1/c3 ,\PWMC/n26 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub1/u20  (
    .a(pnumcntC[20]),
    .b(1'b0),
    .c(\PWMC/sub1/c20 ),
    .o({\PWMC/sub1/c21 ,\PWMC/n26 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub1/u21  (
    .a(pnumcntC[21]),
    .b(1'b0),
    .c(\PWMC/sub1/c21 ),
    .o({\PWMC/sub1/c22 ,\PWMC/n26 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub1/u22  (
    .a(pnumcntC[22]),
    .b(1'b0),
    .c(\PWMC/sub1/c22 ),
    .o({\PWMC/sub1/c23 ,\PWMC/n26 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub1/u23  (
    .a(pnumcntC[23]),
    .b(1'b0),
    .c(\PWMC/sub1/c23 ),
    .o({open_n100,\PWMC/n26 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub1/u3  (
    .a(pnumcntC[3]),
    .b(1'b0),
    .c(\PWMC/sub1/c3 ),
    .o({\PWMC/sub1/c4 ,\PWMC/n26 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub1/u4  (
    .a(pnumcntC[4]),
    .b(1'b0),
    .c(\PWMC/sub1/c4 ),
    .o({\PWMC/sub1/c5 ,\PWMC/n26 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub1/u5  (
    .a(pnumcntC[5]),
    .b(1'b0),
    .c(\PWMC/sub1/c5 ),
    .o({\PWMC/sub1/c6 ,\PWMC/n26 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub1/u6  (
    .a(pnumcntC[6]),
    .b(1'b0),
    .c(\PWMC/sub1/c6 ),
    .o({\PWMC/sub1/c7 ,\PWMC/n26 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub1/u7  (
    .a(pnumcntC[7]),
    .b(1'b0),
    .c(\PWMC/sub1/c7 ),
    .o({\PWMC/sub1/c8 ,\PWMC/n26 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub1/u8  (
    .a(pnumcntC[8]),
    .b(1'b0),
    .c(\PWMC/sub1/c8 ),
    .o({\PWMC/sub1/c9 ,\PWMC/n26 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMC/sub1/u9  (
    .a(pnumcntC[9]),
    .b(1'b0),
    .c(\PWMC/sub1/c9 ),
    .o({\PWMC/sub1/c10 ,\PWMC/n26 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \PWMC/sub1/ucin  (
    .a(1'b0),
    .o({\PWMC/sub1/c0 ,open_n103}));
  reg_ar_as_w1 \PWMD/State_reg  (
    .clk(clk100m),
    .d(\PWMD/n10 ),
    .en(1'b1),
    .reset(~rstn),
    .set(1'b0),
    .q(pwm_state_read[13]));  // src/OnePWM.v(26)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[0]  (
    .i(\PWMD/RemaTxNum[0]_keep ),
    .o(pnumcntD[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[10]  (
    .i(\PWMD/RemaTxNum[10]_keep ),
    .o(pnumcntD[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[11]  (
    .i(\PWMD/RemaTxNum[11]_keep ),
    .o(pnumcntD[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[12]  (
    .i(\PWMD/RemaTxNum[12]_keep ),
    .o(pnumcntD[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[13]  (
    .i(\PWMD/RemaTxNum[13]_keep ),
    .o(pnumcntD[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[14]  (
    .i(\PWMD/RemaTxNum[14]_keep ),
    .o(pnumcntD[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[15]  (
    .i(\PWMD/RemaTxNum[15]_keep ),
    .o(pnumcntD[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[16]  (
    .i(\PWMD/RemaTxNum[16]_keep ),
    .o(pnumcntD[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[17]  (
    .i(\PWMD/RemaTxNum[17]_keep ),
    .o(pnumcntD[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[18]  (
    .i(\PWMD/RemaTxNum[18]_keep ),
    .o(pnumcntD[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[19]  (
    .i(\PWMD/RemaTxNum[19]_keep ),
    .o(pnumcntD[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[1]  (
    .i(\PWMD/RemaTxNum[1]_keep ),
    .o(pnumcntD[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[20]  (
    .i(\PWMD/RemaTxNum[20]_keep ),
    .o(pnumcntD[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[21]  (
    .i(\PWMD/RemaTxNum[21]_keep ),
    .o(pnumcntD[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[22]  (
    .i(\PWMD/RemaTxNum[22]_keep ),
    .o(pnumcntD[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[23]  (
    .i(\PWMD/RemaTxNum[23]_keep ),
    .o(pnumcntD[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[2]  (
    .i(\PWMD/RemaTxNum[2]_keep ),
    .o(pnumcntD[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[3]  (
    .i(\PWMD/RemaTxNum[3]_keep ),
    .o(pnumcntD[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[4]  (
    .i(\PWMD/RemaTxNum[4]_keep ),
    .o(pnumcntD[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[5]  (
    .i(\PWMD/RemaTxNum[5]_keep ),
    .o(pnumcntD[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[6]  (
    .i(\PWMD/RemaTxNum[6]_keep ),
    .o(pnumcntD[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[7]  (
    .i(\PWMD/RemaTxNum[7]_keep ),
    .o(pnumcntD[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[8]  (
    .i(\PWMD/RemaTxNum[8]_keep ),
    .o(pnumcntD[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[9]  (
    .i(\PWMD/RemaTxNum[9]_keep ),
    .o(pnumcntD[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_dir  (
    .i(\PWMD/dir_keep ),
    .o(dir_pad[13]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[0]  (
    .i(\PWMD/pnumr[0]_keep ),
    .o(\PWMD/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[10]  (
    .i(\PWMD/pnumr[10]_keep ),
    .o(\PWMD/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[11]  (
    .i(\PWMD/pnumr[11]_keep ),
    .o(\PWMD/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[12]  (
    .i(\PWMD/pnumr[12]_keep ),
    .o(\PWMD/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[13]  (
    .i(\PWMD/pnumr[13]_keep ),
    .o(\PWMD/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[14]  (
    .i(\PWMD/pnumr[14]_keep ),
    .o(\PWMD/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[15]  (
    .i(\PWMD/pnumr[15]_keep ),
    .o(\PWMD/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[16]  (
    .i(\PWMD/pnumr[16]_keep ),
    .o(\PWMD/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[17]  (
    .i(\PWMD/pnumr[17]_keep ),
    .o(\PWMD/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[18]  (
    .i(\PWMD/pnumr[18]_keep ),
    .o(\PWMD/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[19]  (
    .i(\PWMD/pnumr[19]_keep ),
    .o(\PWMD/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[1]  (
    .i(\PWMD/pnumr[1]_keep ),
    .o(\PWMD/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[20]  (
    .i(\PWMD/pnumr[20]_keep ),
    .o(\PWMD/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[21]  (
    .i(\PWMD/pnumr[21]_keep ),
    .o(\PWMD/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[22]  (
    .i(\PWMD/pnumr[22]_keep ),
    .o(\PWMD/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[23]  (
    .i(\PWMD/pnumr[23]_keep ),
    .o(\PWMD/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[24]  (
    .i(\PWMD/pnumr[24]_keep ),
    .o(\PWMD/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[25]  (
    .i(\PWMD/pnumr[25]_keep ),
    .o(\PWMD/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[26]  (
    .i(\PWMD/pnumr[26]_keep ),
    .o(\PWMD/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[27]  (
    .i(\PWMD/pnumr[27]_keep ),
    .o(\PWMD/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[28]  (
    .i(\PWMD/pnumr[28]_keep ),
    .o(\PWMD/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[29]  (
    .i(\PWMD/pnumr[29]_keep ),
    .o(\PWMD/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[2]  (
    .i(\PWMD/pnumr[2]_keep ),
    .o(\PWMD/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[30]  (
    .i(\PWMD/pnumr[30]_keep ),
    .o(\PWMD/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[31]  (
    .i(\PWMD/pnumr[31]_keep ),
    .o(\PWMD/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[3]  (
    .i(\PWMD/pnumr[3]_keep ),
    .o(\PWMD/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[4]  (
    .i(\PWMD/pnumr[4]_keep ),
    .o(\PWMD/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[5]  (
    .i(\PWMD/pnumr[5]_keep ),
    .o(\PWMD/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[6]  (
    .i(\PWMD/pnumr[6]_keep ),
    .o(\PWMD/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[7]  (
    .i(\PWMD/pnumr[7]_keep ),
    .o(\PWMD/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[8]  (
    .i(\PWMD/pnumr[8]_keep ),
    .o(\PWMD/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[9]  (
    .i(\PWMD/pnumr[9]_keep ),
    .o(\PWMD/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pwm  (
    .i(\PWMD/pwm_keep ),
    .o(pwm_pad[13]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_stopreq  (
    .i(\PWMD/stopreq_keep ),
    .o(\PWMD/stopreq ));  // src/OnePWM.v(14)
  reg_ar_as_w1 \PWMD/dir_reg  (
    .clk(clk100m),
    .d(\PWMD/n32 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/dir_keep ));  // src/OnePWM.v(58)
  reg_sr_as_w1 \PWMD/pwm_reg  (
    .clk(clk100m),
    .d(\pwm[13]_d ),
    .en(1'b1),
    .reset(~\PWMD/u14_sel_is_1_o ),
    .set(1'b0),
    .q(\PWMD/pwm_keep ));  // src/OnePWM.v(45)
  reg_sr_as_w1 \PWMD/reg0_b0  (
    .clk(clk100m),
    .d(\PWMD/n13 [0]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [0]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b1  (
    .clk(clk100m),
    .d(\PWMD/n13 [1]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [1]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b10  (
    .clk(clk100m),
    .d(\PWMD/n13 [10]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [10]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b11  (
    .clk(clk100m),
    .d(\PWMD/n13 [11]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [11]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b12  (
    .clk(clk100m),
    .d(\PWMD/n13 [12]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [12]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b13  (
    .clk(clk100m),
    .d(\PWMD/n13 [13]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [13]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b14  (
    .clk(clk100m),
    .d(\PWMD/n13 [14]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [14]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b15  (
    .clk(clk100m),
    .d(\PWMD/n13 [15]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [15]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b16  (
    .clk(clk100m),
    .d(\PWMD/n13 [16]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [16]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b17  (
    .clk(clk100m),
    .d(\PWMD/n13 [17]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [17]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b18  (
    .clk(clk100m),
    .d(\PWMD/n13 [18]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [18]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b19  (
    .clk(clk100m),
    .d(\PWMD/n13 [19]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [19]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b2  (
    .clk(clk100m),
    .d(\PWMD/n13 [2]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [2]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b20  (
    .clk(clk100m),
    .d(\PWMD/n13 [20]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [20]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b21  (
    .clk(clk100m),
    .d(\PWMD/n13 [21]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [21]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b22  (
    .clk(clk100m),
    .d(\PWMD/n13 [22]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [22]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b23  (
    .clk(clk100m),
    .d(\PWMD/n13 [23]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [23]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b24  (
    .clk(clk100m),
    .d(\PWMD/n13 [24]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [24]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b25  (
    .clk(clk100m),
    .d(\PWMD/n13 [25]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [25]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b26  (
    .clk(clk100m),
    .d(\PWMD/n13 [26]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [26]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b3  (
    .clk(clk100m),
    .d(\PWMD/n13 [3]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [3]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b4  (
    .clk(clk100m),
    .d(\PWMD/n13 [4]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [4]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b5  (
    .clk(clk100m),
    .d(\PWMD/n13 [5]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [5]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b6  (
    .clk(clk100m),
    .d(\PWMD/n13 [6]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [6]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b7  (
    .clk(clk100m),
    .d(\PWMD/n13 [7]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [7]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b8  (
    .clk(clk100m),
    .d(\PWMD/n13 [8]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [8]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b9  (
    .clk(clk100m),
    .d(\PWMD/n13 [9]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b0  (
    .clk(clk100m),
    .d(freqD[0]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [0]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b1  (
    .clk(clk100m),
    .d(freqD[1]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [1]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b10  (
    .clk(clk100m),
    .d(freqD[10]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [10]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b11  (
    .clk(clk100m),
    .d(freqD[11]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [11]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b12  (
    .clk(clk100m),
    .d(freqD[12]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [12]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b13  (
    .clk(clk100m),
    .d(freqD[13]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [13]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b14  (
    .clk(clk100m),
    .d(freqD[14]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [14]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b15  (
    .clk(clk100m),
    .d(freqD[15]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [15]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b16  (
    .clk(clk100m),
    .d(freqD[16]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [16]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b17  (
    .clk(clk100m),
    .d(freqD[17]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [17]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b18  (
    .clk(clk100m),
    .d(freqD[18]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [18]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b19  (
    .clk(clk100m),
    .d(freqD[19]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [19]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b2  (
    .clk(clk100m),
    .d(freqD[2]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [2]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b20  (
    .clk(clk100m),
    .d(freqD[20]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [20]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b21  (
    .clk(clk100m),
    .d(freqD[21]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [21]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b22  (
    .clk(clk100m),
    .d(freqD[22]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [22]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b23  (
    .clk(clk100m),
    .d(freqD[23]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [23]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b24  (
    .clk(clk100m),
    .d(freqD[24]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [24]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b25  (
    .clk(clk100m),
    .d(freqD[25]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [25]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b26  (
    .clk(clk100m),
    .d(freqD[26]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [26]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b3  (
    .clk(clk100m),
    .d(freqD[3]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [3]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b4  (
    .clk(clk100m),
    .d(freqD[4]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [4]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b5  (
    .clk(clk100m),
    .d(freqD[5]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [5]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b6  (
    .clk(clk100m),
    .d(freqD[6]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [6]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b7  (
    .clk(clk100m),
    .d(freqD[7]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [7]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b8  (
    .clk(clk100m),
    .d(freqD[8]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [8]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b9  (
    .clk(clk100m),
    .d(freqD[9]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg2_b0  (
    .clk(clk100m),
    .d(\PWMD/n23 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[0]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b1  (
    .clk(clk100m),
    .d(\PWMD/n23 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[1]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b10  (
    .clk(clk100m),
    .d(\PWMD/n23 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[10]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b11  (
    .clk(clk100m),
    .d(\PWMD/n23 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[11]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b12  (
    .clk(clk100m),
    .d(\PWMD/n23 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[12]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b13  (
    .clk(clk100m),
    .d(\PWMD/n23 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[13]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b14  (
    .clk(clk100m),
    .d(\PWMD/n23 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[14]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b15  (
    .clk(clk100m),
    .d(\PWMD/n23 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[15]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b16  (
    .clk(clk100m),
    .d(\PWMD/n23 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[16]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b17  (
    .clk(clk100m),
    .d(\PWMD/n23 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[17]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b18  (
    .clk(clk100m),
    .d(\PWMD/n23 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[18]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b19  (
    .clk(clk100m),
    .d(\PWMD/n23 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[19]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b2  (
    .clk(clk100m),
    .d(\PWMD/n23 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[2]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b20  (
    .clk(clk100m),
    .d(\PWMD/n23 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[20]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b21  (
    .clk(clk100m),
    .d(\PWMD/n23 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[21]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b22  (
    .clk(clk100m),
    .d(\PWMD/n23 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[22]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b23  (
    .clk(clk100m),
    .d(\PWMD/n23 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[23]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b24  (
    .clk(clk100m),
    .d(\PWMD/n23 [24]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[24]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b25  (
    .clk(clk100m),
    .d(\PWMD/n23 [25]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[25]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b26  (
    .clk(clk100m),
    .d(\PWMD/n23 [26]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[26]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b27  (
    .clk(clk100m),
    .d(\PWMD/n23 [27]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[27]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b28  (
    .clk(clk100m),
    .d(\PWMD/n23 [28]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[28]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b29  (
    .clk(clk100m),
    .d(\PWMD/n23 [29]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[29]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b3  (
    .clk(clk100m),
    .d(\PWMD/n23 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[3]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b30  (
    .clk(clk100m),
    .d(\PWMD/n23 [30]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[30]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b31  (
    .clk(clk100m),
    .d(\PWMD/n23 [31]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[31]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b4  (
    .clk(clk100m),
    .d(\PWMD/n23 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[4]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b5  (
    .clk(clk100m),
    .d(\PWMD/n23 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[5]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b6  (
    .clk(clk100m),
    .d(\PWMD/n23 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[6]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b7  (
    .clk(clk100m),
    .d(\PWMD/n23 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[7]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b8  (
    .clk(clk100m),
    .d(\PWMD/n23 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[8]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b9  (
    .clk(clk100m),
    .d(\PWMD/n23 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[9]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg3_b0  (
    .clk(clk100m),
    .d(\PWMD/n31 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[0]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b1  (
    .clk(clk100m),
    .d(\PWMD/n31 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[1]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b10  (
    .clk(clk100m),
    .d(\PWMD/n31 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[10]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b11  (
    .clk(clk100m),
    .d(\PWMD/n31 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[11]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b12  (
    .clk(clk100m),
    .d(\PWMD/n31 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[12]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b13  (
    .clk(clk100m),
    .d(\PWMD/n31 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[13]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b14  (
    .clk(clk100m),
    .d(\PWMD/n31 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[14]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b15  (
    .clk(clk100m),
    .d(\PWMD/n31 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[15]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b16  (
    .clk(clk100m),
    .d(\PWMD/n31 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[16]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b17  (
    .clk(clk100m),
    .d(\PWMD/n31 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[17]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b18  (
    .clk(clk100m),
    .d(\PWMD/n31 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[18]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b19  (
    .clk(clk100m),
    .d(\PWMD/n31 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[19]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b2  (
    .clk(clk100m),
    .d(\PWMD/n31 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[2]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b20  (
    .clk(clk100m),
    .d(\PWMD/n31 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[20]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b21  (
    .clk(clk100m),
    .d(\PWMD/n31 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[21]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b22  (
    .clk(clk100m),
    .d(\PWMD/n31 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[22]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b23  (
    .clk(clk100m),
    .d(\PWMD/n31 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[23]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b3  (
    .clk(clk100m),
    .d(\PWMD/n31 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[3]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b4  (
    .clk(clk100m),
    .d(\PWMD/n31 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[4]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b5  (
    .clk(clk100m),
    .d(\PWMD/n31 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[5]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b6  (
    .clk(clk100m),
    .d(\PWMD/n31 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[6]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b7  (
    .clk(clk100m),
    .d(\PWMD/n31 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[7]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b8  (
    .clk(clk100m),
    .d(\PWMD/n31 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[8]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b9  (
    .clk(clk100m),
    .d(\PWMD/n31 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[9]_keep ));  // src/OnePWM.v(58)
  reg_ar_ss_w1 \PWMD/stopreq_reg  (
    .clk(clk100m),
    .d(\PWMD/n1 ),
    .en(1'b1),
    .reset(1'b0),
    .set(pwm_start_stop[13]),
    .q(\PWMD/stopreq_keep ));  // src/OnePWM.v(15)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub0/u0  (
    .a(\PWMD/FreCnt [0]),
    .b(1'b1),
    .c(\PWMD/sub0/c0 ),
    .o({\PWMD/sub0/c1 ,\PWMD/n12 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub0/u1  (
    .a(\PWMD/FreCnt [1]),
    .b(1'b0),
    .c(\PWMD/sub0/c1 ),
    .o({\PWMD/sub0/c2 ,\PWMD/n12 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub0/u10  (
    .a(\PWMD/FreCnt [10]),
    .b(1'b0),
    .c(\PWMD/sub0/c10 ),
    .o({\PWMD/sub0/c11 ,\PWMD/n12 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub0/u11  (
    .a(\PWMD/FreCnt [11]),
    .b(1'b0),
    .c(\PWMD/sub0/c11 ),
    .o({\PWMD/sub0/c12 ,\PWMD/n12 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub0/u12  (
    .a(\PWMD/FreCnt [12]),
    .b(1'b0),
    .c(\PWMD/sub0/c12 ),
    .o({\PWMD/sub0/c13 ,\PWMD/n12 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub0/u13  (
    .a(\PWMD/FreCnt [13]),
    .b(1'b0),
    .c(\PWMD/sub0/c13 ),
    .o({\PWMD/sub0/c14 ,\PWMD/n12 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub0/u14  (
    .a(\PWMD/FreCnt [14]),
    .b(1'b0),
    .c(\PWMD/sub0/c14 ),
    .o({\PWMD/sub0/c15 ,\PWMD/n12 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub0/u15  (
    .a(\PWMD/FreCnt [15]),
    .b(1'b0),
    .c(\PWMD/sub0/c15 ),
    .o({\PWMD/sub0/c16 ,\PWMD/n12 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub0/u16  (
    .a(\PWMD/FreCnt [16]),
    .b(1'b0),
    .c(\PWMD/sub0/c16 ),
    .o({\PWMD/sub0/c17 ,\PWMD/n12 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub0/u17  (
    .a(\PWMD/FreCnt [17]),
    .b(1'b0),
    .c(\PWMD/sub0/c17 ),
    .o({\PWMD/sub0/c18 ,\PWMD/n12 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub0/u18  (
    .a(\PWMD/FreCnt [18]),
    .b(1'b0),
    .c(\PWMD/sub0/c18 ),
    .o({\PWMD/sub0/c19 ,\PWMD/n12 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub0/u19  (
    .a(\PWMD/FreCnt [19]),
    .b(1'b0),
    .c(\PWMD/sub0/c19 ),
    .o({\PWMD/sub0/c20 ,\PWMD/n12 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub0/u2  (
    .a(\PWMD/FreCnt [2]),
    .b(1'b0),
    .c(\PWMD/sub0/c2 ),
    .o({\PWMD/sub0/c3 ,\PWMD/n12 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub0/u20  (
    .a(\PWMD/FreCnt [20]),
    .b(1'b0),
    .c(\PWMD/sub0/c20 ),
    .o({\PWMD/sub0/c21 ,\PWMD/n12 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub0/u21  (
    .a(\PWMD/FreCnt [21]),
    .b(1'b0),
    .c(\PWMD/sub0/c21 ),
    .o({\PWMD/sub0/c22 ,\PWMD/n12 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub0/u22  (
    .a(\PWMD/FreCnt [22]),
    .b(1'b0),
    .c(\PWMD/sub0/c22 ),
    .o({\PWMD/sub0/c23 ,\PWMD/n12 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub0/u23  (
    .a(\PWMD/FreCnt [23]),
    .b(1'b0),
    .c(\PWMD/sub0/c23 ),
    .o({\PWMD/sub0/c24 ,\PWMD/n12 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub0/u24  (
    .a(\PWMD/FreCnt [24]),
    .b(1'b0),
    .c(\PWMD/sub0/c24 ),
    .o({\PWMD/sub0/c25 ,\PWMD/n12 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub0/u25  (
    .a(\PWMD/FreCnt [25]),
    .b(1'b0),
    .c(\PWMD/sub0/c25 ),
    .o({\PWMD/sub0/c26 ,\PWMD/n12 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub0/u26  (
    .a(\PWMD/FreCnt [26]),
    .b(1'b0),
    .c(\PWMD/sub0/c26 ),
    .o({open_n104,\PWMD/n12 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub0/u3  (
    .a(\PWMD/FreCnt [3]),
    .b(1'b0),
    .c(\PWMD/sub0/c3 ),
    .o({\PWMD/sub0/c4 ,\PWMD/n12 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub0/u4  (
    .a(\PWMD/FreCnt [4]),
    .b(1'b0),
    .c(\PWMD/sub0/c4 ),
    .o({\PWMD/sub0/c5 ,\PWMD/n12 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub0/u5  (
    .a(\PWMD/FreCnt [5]),
    .b(1'b0),
    .c(\PWMD/sub0/c5 ),
    .o({\PWMD/sub0/c6 ,\PWMD/n12 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub0/u6  (
    .a(\PWMD/FreCnt [6]),
    .b(1'b0),
    .c(\PWMD/sub0/c6 ),
    .o({\PWMD/sub0/c7 ,\PWMD/n12 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub0/u7  (
    .a(\PWMD/FreCnt [7]),
    .b(1'b0),
    .c(\PWMD/sub0/c7 ),
    .o({\PWMD/sub0/c8 ,\PWMD/n12 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub0/u8  (
    .a(\PWMD/FreCnt [8]),
    .b(1'b0),
    .c(\PWMD/sub0/c8 ),
    .o({\PWMD/sub0/c9 ,\PWMD/n12 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub0/u9  (
    .a(\PWMD/FreCnt [9]),
    .b(1'b0),
    .c(\PWMD/sub0/c9 ),
    .o({\PWMD/sub0/c10 ,\PWMD/n12 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \PWMD/sub0/ucin  (
    .a(1'b0),
    .o({\PWMD/sub0/c0 ,open_n107}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub1/u0  (
    .a(pnumcntD[0]),
    .b(1'b1),
    .c(\PWMD/sub1/c0 ),
    .o({\PWMD/sub1/c1 ,\PWMD/n26 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub1/u1  (
    .a(pnumcntD[1]),
    .b(1'b0),
    .c(\PWMD/sub1/c1 ),
    .o({\PWMD/sub1/c2 ,\PWMD/n26 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub1/u10  (
    .a(pnumcntD[10]),
    .b(1'b0),
    .c(\PWMD/sub1/c10 ),
    .o({\PWMD/sub1/c11 ,\PWMD/n26 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub1/u11  (
    .a(pnumcntD[11]),
    .b(1'b0),
    .c(\PWMD/sub1/c11 ),
    .o({\PWMD/sub1/c12 ,\PWMD/n26 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub1/u12  (
    .a(pnumcntD[12]),
    .b(1'b0),
    .c(\PWMD/sub1/c12 ),
    .o({\PWMD/sub1/c13 ,\PWMD/n26 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub1/u13  (
    .a(pnumcntD[13]),
    .b(1'b0),
    .c(\PWMD/sub1/c13 ),
    .o({\PWMD/sub1/c14 ,\PWMD/n26 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub1/u14  (
    .a(pnumcntD[14]),
    .b(1'b0),
    .c(\PWMD/sub1/c14 ),
    .o({\PWMD/sub1/c15 ,\PWMD/n26 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub1/u15  (
    .a(pnumcntD[15]),
    .b(1'b0),
    .c(\PWMD/sub1/c15 ),
    .o({\PWMD/sub1/c16 ,\PWMD/n26 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub1/u16  (
    .a(pnumcntD[16]),
    .b(1'b0),
    .c(\PWMD/sub1/c16 ),
    .o({\PWMD/sub1/c17 ,\PWMD/n26 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub1/u17  (
    .a(pnumcntD[17]),
    .b(1'b0),
    .c(\PWMD/sub1/c17 ),
    .o({\PWMD/sub1/c18 ,\PWMD/n26 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub1/u18  (
    .a(pnumcntD[18]),
    .b(1'b0),
    .c(\PWMD/sub1/c18 ),
    .o({\PWMD/sub1/c19 ,\PWMD/n26 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub1/u19  (
    .a(pnumcntD[19]),
    .b(1'b0),
    .c(\PWMD/sub1/c19 ),
    .o({\PWMD/sub1/c20 ,\PWMD/n26 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub1/u2  (
    .a(pnumcntD[2]),
    .b(1'b0),
    .c(\PWMD/sub1/c2 ),
    .o({\PWMD/sub1/c3 ,\PWMD/n26 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub1/u20  (
    .a(pnumcntD[20]),
    .b(1'b0),
    .c(\PWMD/sub1/c20 ),
    .o({\PWMD/sub1/c21 ,\PWMD/n26 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub1/u21  (
    .a(pnumcntD[21]),
    .b(1'b0),
    .c(\PWMD/sub1/c21 ),
    .o({\PWMD/sub1/c22 ,\PWMD/n26 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub1/u22  (
    .a(pnumcntD[22]),
    .b(1'b0),
    .c(\PWMD/sub1/c22 ),
    .o({\PWMD/sub1/c23 ,\PWMD/n26 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub1/u23  (
    .a(pnumcntD[23]),
    .b(1'b0),
    .c(\PWMD/sub1/c23 ),
    .o({open_n108,\PWMD/n26 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub1/u3  (
    .a(pnumcntD[3]),
    .b(1'b0),
    .c(\PWMD/sub1/c3 ),
    .o({\PWMD/sub1/c4 ,\PWMD/n26 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub1/u4  (
    .a(pnumcntD[4]),
    .b(1'b0),
    .c(\PWMD/sub1/c4 ),
    .o({\PWMD/sub1/c5 ,\PWMD/n26 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub1/u5  (
    .a(pnumcntD[5]),
    .b(1'b0),
    .c(\PWMD/sub1/c5 ),
    .o({\PWMD/sub1/c6 ,\PWMD/n26 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub1/u6  (
    .a(pnumcntD[6]),
    .b(1'b0),
    .c(\PWMD/sub1/c6 ),
    .o({\PWMD/sub1/c7 ,\PWMD/n26 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub1/u7  (
    .a(pnumcntD[7]),
    .b(1'b0),
    .c(\PWMD/sub1/c7 ),
    .o({\PWMD/sub1/c8 ,\PWMD/n26 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub1/u8  (
    .a(pnumcntD[8]),
    .b(1'b0),
    .c(\PWMD/sub1/c8 ),
    .o({\PWMD/sub1/c9 ,\PWMD/n26 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMD/sub1/u9  (
    .a(pnumcntD[9]),
    .b(1'b0),
    .c(\PWMD/sub1/c9 ),
    .o({\PWMD/sub1/c10 ,\PWMD/n26 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \PWMD/sub1/ucin  (
    .a(1'b0),
    .o({\PWMD/sub1/c0 ,open_n111}));
  reg_ar_as_w1 \PWME/State_reg  (
    .clk(clk100m),
    .d(\PWME/n10 ),
    .en(1'b1),
    .reset(~rstn),
    .set(1'b0),
    .q(pwm_state_read[14]));  // src/OnePWM.v(26)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[0]  (
    .i(\PWME/RemaTxNum[0]_keep ),
    .o(pnumcntE[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[10]  (
    .i(\PWME/RemaTxNum[10]_keep ),
    .o(pnumcntE[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[11]  (
    .i(\PWME/RemaTxNum[11]_keep ),
    .o(pnumcntE[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[12]  (
    .i(\PWME/RemaTxNum[12]_keep ),
    .o(pnumcntE[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[13]  (
    .i(\PWME/RemaTxNum[13]_keep ),
    .o(pnumcntE[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[14]  (
    .i(\PWME/RemaTxNum[14]_keep ),
    .o(pnumcntE[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[15]  (
    .i(\PWME/RemaTxNum[15]_keep ),
    .o(pnumcntE[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[16]  (
    .i(\PWME/RemaTxNum[16]_keep ),
    .o(pnumcntE[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[17]  (
    .i(\PWME/RemaTxNum[17]_keep ),
    .o(pnumcntE[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[18]  (
    .i(\PWME/RemaTxNum[18]_keep ),
    .o(pnumcntE[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[19]  (
    .i(\PWME/RemaTxNum[19]_keep ),
    .o(pnumcntE[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[1]  (
    .i(\PWME/RemaTxNum[1]_keep ),
    .o(pnumcntE[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[20]  (
    .i(\PWME/RemaTxNum[20]_keep ),
    .o(pnumcntE[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[21]  (
    .i(\PWME/RemaTxNum[21]_keep ),
    .o(pnumcntE[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[22]  (
    .i(\PWME/RemaTxNum[22]_keep ),
    .o(pnumcntE[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[23]  (
    .i(\PWME/RemaTxNum[23]_keep ),
    .o(pnumcntE[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[2]  (
    .i(\PWME/RemaTxNum[2]_keep ),
    .o(pnumcntE[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[3]  (
    .i(\PWME/RemaTxNum[3]_keep ),
    .o(pnumcntE[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[4]  (
    .i(\PWME/RemaTxNum[4]_keep ),
    .o(pnumcntE[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[5]  (
    .i(\PWME/RemaTxNum[5]_keep ),
    .o(pnumcntE[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[6]  (
    .i(\PWME/RemaTxNum[6]_keep ),
    .o(pnumcntE[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[7]  (
    .i(\PWME/RemaTxNum[7]_keep ),
    .o(pnumcntE[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[8]  (
    .i(\PWME/RemaTxNum[8]_keep ),
    .o(pnumcntE[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[9]  (
    .i(\PWME/RemaTxNum[9]_keep ),
    .o(pnumcntE[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_dir  (
    .i(\PWME/dir_keep ),
    .o(dir_pad[14]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[0]  (
    .i(\PWME/pnumr[0]_keep ),
    .o(\PWME/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[10]  (
    .i(\PWME/pnumr[10]_keep ),
    .o(\PWME/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[11]  (
    .i(\PWME/pnumr[11]_keep ),
    .o(\PWME/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[12]  (
    .i(\PWME/pnumr[12]_keep ),
    .o(\PWME/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[13]  (
    .i(\PWME/pnumr[13]_keep ),
    .o(\PWME/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[14]  (
    .i(\PWME/pnumr[14]_keep ),
    .o(\PWME/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[15]  (
    .i(\PWME/pnumr[15]_keep ),
    .o(\PWME/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[16]  (
    .i(\PWME/pnumr[16]_keep ),
    .o(\PWME/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[17]  (
    .i(\PWME/pnumr[17]_keep ),
    .o(\PWME/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[18]  (
    .i(\PWME/pnumr[18]_keep ),
    .o(\PWME/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[19]  (
    .i(\PWME/pnumr[19]_keep ),
    .o(\PWME/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[1]  (
    .i(\PWME/pnumr[1]_keep ),
    .o(\PWME/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[20]  (
    .i(\PWME/pnumr[20]_keep ),
    .o(\PWME/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[21]  (
    .i(\PWME/pnumr[21]_keep ),
    .o(\PWME/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[22]  (
    .i(\PWME/pnumr[22]_keep ),
    .o(\PWME/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[23]  (
    .i(\PWME/pnumr[23]_keep ),
    .o(\PWME/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[24]  (
    .i(\PWME/pnumr[24]_keep ),
    .o(\PWME/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[25]  (
    .i(\PWME/pnumr[25]_keep ),
    .o(\PWME/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[26]  (
    .i(\PWME/pnumr[26]_keep ),
    .o(\PWME/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[27]  (
    .i(\PWME/pnumr[27]_keep ),
    .o(\PWME/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[28]  (
    .i(\PWME/pnumr[28]_keep ),
    .o(\PWME/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[29]  (
    .i(\PWME/pnumr[29]_keep ),
    .o(\PWME/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[2]  (
    .i(\PWME/pnumr[2]_keep ),
    .o(\PWME/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[30]  (
    .i(\PWME/pnumr[30]_keep ),
    .o(\PWME/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[31]  (
    .i(\PWME/pnumr[31]_keep ),
    .o(\PWME/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[3]  (
    .i(\PWME/pnumr[3]_keep ),
    .o(\PWME/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[4]  (
    .i(\PWME/pnumr[4]_keep ),
    .o(\PWME/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[5]  (
    .i(\PWME/pnumr[5]_keep ),
    .o(\PWME/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[6]  (
    .i(\PWME/pnumr[6]_keep ),
    .o(\PWME/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[7]  (
    .i(\PWME/pnumr[7]_keep ),
    .o(\PWME/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[8]  (
    .i(\PWME/pnumr[8]_keep ),
    .o(\PWME/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[9]  (
    .i(\PWME/pnumr[9]_keep ),
    .o(\PWME/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pwm  (
    .i(\PWME/pwm_keep ),
    .o(pwm_pad[14]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_stopreq  (
    .i(\PWME/stopreq_keep ),
    .o(\PWME/stopreq ));  // src/OnePWM.v(14)
  reg_ar_as_w1 \PWME/dir_reg  (
    .clk(clk100m),
    .d(\PWME/n32 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/dir_keep ));  // src/OnePWM.v(58)
  reg_sr_as_w1 \PWME/pwm_reg  (
    .clk(clk100m),
    .d(\pwm[14]_d ),
    .en(1'b1),
    .reset(~\PWME/u14_sel_is_1_o ),
    .set(1'b0),
    .q(\PWME/pwm_keep ));  // src/OnePWM.v(45)
  reg_sr_as_w1 \PWME/reg0_b0  (
    .clk(clk100m),
    .d(\PWME/n13 [0]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [0]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b1  (
    .clk(clk100m),
    .d(\PWME/n13 [1]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [1]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b10  (
    .clk(clk100m),
    .d(\PWME/n13 [10]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [10]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b11  (
    .clk(clk100m),
    .d(\PWME/n13 [11]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [11]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b12  (
    .clk(clk100m),
    .d(\PWME/n13 [12]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [12]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b13  (
    .clk(clk100m),
    .d(\PWME/n13 [13]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [13]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b14  (
    .clk(clk100m),
    .d(\PWME/n13 [14]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [14]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b15  (
    .clk(clk100m),
    .d(\PWME/n13 [15]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [15]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b16  (
    .clk(clk100m),
    .d(\PWME/n13 [16]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [16]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b17  (
    .clk(clk100m),
    .d(\PWME/n13 [17]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [17]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b18  (
    .clk(clk100m),
    .d(\PWME/n13 [18]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [18]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b19  (
    .clk(clk100m),
    .d(\PWME/n13 [19]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [19]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b2  (
    .clk(clk100m),
    .d(\PWME/n13 [2]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [2]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b20  (
    .clk(clk100m),
    .d(\PWME/n13 [20]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [20]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b21  (
    .clk(clk100m),
    .d(\PWME/n13 [21]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [21]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b22  (
    .clk(clk100m),
    .d(\PWME/n13 [22]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [22]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b23  (
    .clk(clk100m),
    .d(\PWME/n13 [23]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [23]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b24  (
    .clk(clk100m),
    .d(\PWME/n13 [24]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [24]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b25  (
    .clk(clk100m),
    .d(\PWME/n13 [25]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [25]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b26  (
    .clk(clk100m),
    .d(\PWME/n13 [26]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [26]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b3  (
    .clk(clk100m),
    .d(\PWME/n13 [3]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [3]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b4  (
    .clk(clk100m),
    .d(\PWME/n13 [4]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [4]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b5  (
    .clk(clk100m),
    .d(\PWME/n13 [5]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [5]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b6  (
    .clk(clk100m),
    .d(\PWME/n13 [6]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [6]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b7  (
    .clk(clk100m),
    .d(\PWME/n13 [7]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [7]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b8  (
    .clk(clk100m),
    .d(\PWME/n13 [8]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [8]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b9  (
    .clk(clk100m),
    .d(\PWME/n13 [9]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b0  (
    .clk(clk100m),
    .d(freqE[0]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [0]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b1  (
    .clk(clk100m),
    .d(freqE[1]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [1]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b10  (
    .clk(clk100m),
    .d(freqE[10]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [10]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b11  (
    .clk(clk100m),
    .d(freqE[11]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [11]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b12  (
    .clk(clk100m),
    .d(freqE[12]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [12]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b13  (
    .clk(clk100m),
    .d(freqE[13]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [13]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b14  (
    .clk(clk100m),
    .d(freqE[14]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [14]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b15  (
    .clk(clk100m),
    .d(freqE[15]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [15]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b16  (
    .clk(clk100m),
    .d(freqE[16]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [16]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b17  (
    .clk(clk100m),
    .d(freqE[17]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [17]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b18  (
    .clk(clk100m),
    .d(freqE[18]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [18]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b19  (
    .clk(clk100m),
    .d(freqE[19]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [19]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b2  (
    .clk(clk100m),
    .d(freqE[2]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [2]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b20  (
    .clk(clk100m),
    .d(freqE[20]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [20]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b21  (
    .clk(clk100m),
    .d(freqE[21]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [21]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b22  (
    .clk(clk100m),
    .d(freqE[22]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [22]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b23  (
    .clk(clk100m),
    .d(freqE[23]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [23]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b24  (
    .clk(clk100m),
    .d(freqE[24]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [24]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b25  (
    .clk(clk100m),
    .d(freqE[25]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [25]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b26  (
    .clk(clk100m),
    .d(freqE[26]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [26]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b3  (
    .clk(clk100m),
    .d(freqE[3]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [3]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b4  (
    .clk(clk100m),
    .d(freqE[4]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [4]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b5  (
    .clk(clk100m),
    .d(freqE[5]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [5]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b6  (
    .clk(clk100m),
    .d(freqE[6]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [6]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b7  (
    .clk(clk100m),
    .d(freqE[7]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [7]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b8  (
    .clk(clk100m),
    .d(freqE[8]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [8]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b9  (
    .clk(clk100m),
    .d(freqE[9]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg2_b0  (
    .clk(clk100m),
    .d(\PWME/n23 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[0]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b1  (
    .clk(clk100m),
    .d(\PWME/n23 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[1]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b10  (
    .clk(clk100m),
    .d(\PWME/n23 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[10]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b11  (
    .clk(clk100m),
    .d(\PWME/n23 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[11]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b12  (
    .clk(clk100m),
    .d(\PWME/n23 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[12]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b13  (
    .clk(clk100m),
    .d(\PWME/n23 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[13]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b14  (
    .clk(clk100m),
    .d(\PWME/n23 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[14]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b15  (
    .clk(clk100m),
    .d(\PWME/n23 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[15]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b16  (
    .clk(clk100m),
    .d(\PWME/n23 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[16]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b17  (
    .clk(clk100m),
    .d(\PWME/n23 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[17]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b18  (
    .clk(clk100m),
    .d(\PWME/n23 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[18]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b19  (
    .clk(clk100m),
    .d(\PWME/n23 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[19]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b2  (
    .clk(clk100m),
    .d(\PWME/n23 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[2]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b20  (
    .clk(clk100m),
    .d(\PWME/n23 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[20]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b21  (
    .clk(clk100m),
    .d(\PWME/n23 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[21]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b22  (
    .clk(clk100m),
    .d(\PWME/n23 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[22]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b23  (
    .clk(clk100m),
    .d(\PWME/n23 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[23]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b24  (
    .clk(clk100m),
    .d(\PWME/n23 [24]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[24]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b25  (
    .clk(clk100m),
    .d(\PWME/n23 [25]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[25]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b26  (
    .clk(clk100m),
    .d(\PWME/n23 [26]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[26]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b27  (
    .clk(clk100m),
    .d(\PWME/n23 [27]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[27]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b28  (
    .clk(clk100m),
    .d(\PWME/n23 [28]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[28]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b29  (
    .clk(clk100m),
    .d(\PWME/n23 [29]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[29]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b3  (
    .clk(clk100m),
    .d(\PWME/n23 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[3]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b30  (
    .clk(clk100m),
    .d(\PWME/n23 [30]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[30]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b31  (
    .clk(clk100m),
    .d(\PWME/n23 [31]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[31]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b4  (
    .clk(clk100m),
    .d(\PWME/n23 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[4]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b5  (
    .clk(clk100m),
    .d(\PWME/n23 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[5]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b6  (
    .clk(clk100m),
    .d(\PWME/n23 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[6]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b7  (
    .clk(clk100m),
    .d(\PWME/n23 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[7]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b8  (
    .clk(clk100m),
    .d(\PWME/n23 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[8]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b9  (
    .clk(clk100m),
    .d(\PWME/n23 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[9]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg3_b0  (
    .clk(clk100m),
    .d(\PWME/n31 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[0]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b1  (
    .clk(clk100m),
    .d(\PWME/n31 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[1]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b10  (
    .clk(clk100m),
    .d(\PWME/n31 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[10]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b11  (
    .clk(clk100m),
    .d(\PWME/n31 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[11]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b12  (
    .clk(clk100m),
    .d(\PWME/n31 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[12]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b13  (
    .clk(clk100m),
    .d(\PWME/n31 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[13]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b14  (
    .clk(clk100m),
    .d(\PWME/n31 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[14]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b15  (
    .clk(clk100m),
    .d(\PWME/n31 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[15]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b16  (
    .clk(clk100m),
    .d(\PWME/n31 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[16]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b17  (
    .clk(clk100m),
    .d(\PWME/n31 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[17]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b18  (
    .clk(clk100m),
    .d(\PWME/n31 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[18]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b19  (
    .clk(clk100m),
    .d(\PWME/n31 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[19]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b2  (
    .clk(clk100m),
    .d(\PWME/n31 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[2]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b20  (
    .clk(clk100m),
    .d(\PWME/n31 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[20]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b21  (
    .clk(clk100m),
    .d(\PWME/n31 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[21]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b22  (
    .clk(clk100m),
    .d(\PWME/n31 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[22]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b23  (
    .clk(clk100m),
    .d(\PWME/n31 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[23]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b3  (
    .clk(clk100m),
    .d(\PWME/n31 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[3]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b4  (
    .clk(clk100m),
    .d(\PWME/n31 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[4]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b5  (
    .clk(clk100m),
    .d(\PWME/n31 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[5]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b6  (
    .clk(clk100m),
    .d(\PWME/n31 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[6]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b7  (
    .clk(clk100m),
    .d(\PWME/n31 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[7]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b8  (
    .clk(clk100m),
    .d(\PWME/n31 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[8]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b9  (
    .clk(clk100m),
    .d(\PWME/n31 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[9]_keep ));  // src/OnePWM.v(58)
  reg_ar_ss_w1 \PWME/stopreq_reg  (
    .clk(clk100m),
    .d(\PWME/n1 ),
    .en(1'b1),
    .reset(1'b0),
    .set(pwm_start_stop[14]),
    .q(\PWME/stopreq_keep ));  // src/OnePWM.v(15)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub0/u0  (
    .a(\PWME/FreCnt [0]),
    .b(1'b1),
    .c(\PWME/sub0/c0 ),
    .o({\PWME/sub0/c1 ,\PWME/n12 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub0/u1  (
    .a(\PWME/FreCnt [1]),
    .b(1'b0),
    .c(\PWME/sub0/c1 ),
    .o({\PWME/sub0/c2 ,\PWME/n12 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub0/u10  (
    .a(\PWME/FreCnt [10]),
    .b(1'b0),
    .c(\PWME/sub0/c10 ),
    .o({\PWME/sub0/c11 ,\PWME/n12 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub0/u11  (
    .a(\PWME/FreCnt [11]),
    .b(1'b0),
    .c(\PWME/sub0/c11 ),
    .o({\PWME/sub0/c12 ,\PWME/n12 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub0/u12  (
    .a(\PWME/FreCnt [12]),
    .b(1'b0),
    .c(\PWME/sub0/c12 ),
    .o({\PWME/sub0/c13 ,\PWME/n12 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub0/u13  (
    .a(\PWME/FreCnt [13]),
    .b(1'b0),
    .c(\PWME/sub0/c13 ),
    .o({\PWME/sub0/c14 ,\PWME/n12 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub0/u14  (
    .a(\PWME/FreCnt [14]),
    .b(1'b0),
    .c(\PWME/sub0/c14 ),
    .o({\PWME/sub0/c15 ,\PWME/n12 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub0/u15  (
    .a(\PWME/FreCnt [15]),
    .b(1'b0),
    .c(\PWME/sub0/c15 ),
    .o({\PWME/sub0/c16 ,\PWME/n12 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub0/u16  (
    .a(\PWME/FreCnt [16]),
    .b(1'b0),
    .c(\PWME/sub0/c16 ),
    .o({\PWME/sub0/c17 ,\PWME/n12 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub0/u17  (
    .a(\PWME/FreCnt [17]),
    .b(1'b0),
    .c(\PWME/sub0/c17 ),
    .o({\PWME/sub0/c18 ,\PWME/n12 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub0/u18  (
    .a(\PWME/FreCnt [18]),
    .b(1'b0),
    .c(\PWME/sub0/c18 ),
    .o({\PWME/sub0/c19 ,\PWME/n12 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub0/u19  (
    .a(\PWME/FreCnt [19]),
    .b(1'b0),
    .c(\PWME/sub0/c19 ),
    .o({\PWME/sub0/c20 ,\PWME/n12 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub0/u2  (
    .a(\PWME/FreCnt [2]),
    .b(1'b0),
    .c(\PWME/sub0/c2 ),
    .o({\PWME/sub0/c3 ,\PWME/n12 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub0/u20  (
    .a(\PWME/FreCnt [20]),
    .b(1'b0),
    .c(\PWME/sub0/c20 ),
    .o({\PWME/sub0/c21 ,\PWME/n12 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub0/u21  (
    .a(\PWME/FreCnt [21]),
    .b(1'b0),
    .c(\PWME/sub0/c21 ),
    .o({\PWME/sub0/c22 ,\PWME/n12 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub0/u22  (
    .a(\PWME/FreCnt [22]),
    .b(1'b0),
    .c(\PWME/sub0/c22 ),
    .o({\PWME/sub0/c23 ,\PWME/n12 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub0/u23  (
    .a(\PWME/FreCnt [23]),
    .b(1'b0),
    .c(\PWME/sub0/c23 ),
    .o({\PWME/sub0/c24 ,\PWME/n12 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub0/u24  (
    .a(\PWME/FreCnt [24]),
    .b(1'b0),
    .c(\PWME/sub0/c24 ),
    .o({\PWME/sub0/c25 ,\PWME/n12 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub0/u25  (
    .a(\PWME/FreCnt [25]),
    .b(1'b0),
    .c(\PWME/sub0/c25 ),
    .o({\PWME/sub0/c26 ,\PWME/n12 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub0/u26  (
    .a(\PWME/FreCnt [26]),
    .b(1'b0),
    .c(\PWME/sub0/c26 ),
    .o({open_n112,\PWME/n12 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub0/u3  (
    .a(\PWME/FreCnt [3]),
    .b(1'b0),
    .c(\PWME/sub0/c3 ),
    .o({\PWME/sub0/c4 ,\PWME/n12 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub0/u4  (
    .a(\PWME/FreCnt [4]),
    .b(1'b0),
    .c(\PWME/sub0/c4 ),
    .o({\PWME/sub0/c5 ,\PWME/n12 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub0/u5  (
    .a(\PWME/FreCnt [5]),
    .b(1'b0),
    .c(\PWME/sub0/c5 ),
    .o({\PWME/sub0/c6 ,\PWME/n12 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub0/u6  (
    .a(\PWME/FreCnt [6]),
    .b(1'b0),
    .c(\PWME/sub0/c6 ),
    .o({\PWME/sub0/c7 ,\PWME/n12 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub0/u7  (
    .a(\PWME/FreCnt [7]),
    .b(1'b0),
    .c(\PWME/sub0/c7 ),
    .o({\PWME/sub0/c8 ,\PWME/n12 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub0/u8  (
    .a(\PWME/FreCnt [8]),
    .b(1'b0),
    .c(\PWME/sub0/c8 ),
    .o({\PWME/sub0/c9 ,\PWME/n12 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub0/u9  (
    .a(\PWME/FreCnt [9]),
    .b(1'b0),
    .c(\PWME/sub0/c9 ),
    .o({\PWME/sub0/c10 ,\PWME/n12 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \PWME/sub0/ucin  (
    .a(1'b0),
    .o({\PWME/sub0/c0 ,open_n115}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub1/u0  (
    .a(pnumcntE[0]),
    .b(1'b1),
    .c(\PWME/sub1/c0 ),
    .o({\PWME/sub1/c1 ,\PWME/n26 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub1/u1  (
    .a(pnumcntE[1]),
    .b(1'b0),
    .c(\PWME/sub1/c1 ),
    .o({\PWME/sub1/c2 ,\PWME/n26 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub1/u10  (
    .a(pnumcntE[10]),
    .b(1'b0),
    .c(\PWME/sub1/c10 ),
    .o({\PWME/sub1/c11 ,\PWME/n26 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub1/u11  (
    .a(pnumcntE[11]),
    .b(1'b0),
    .c(\PWME/sub1/c11 ),
    .o({\PWME/sub1/c12 ,\PWME/n26 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub1/u12  (
    .a(pnumcntE[12]),
    .b(1'b0),
    .c(\PWME/sub1/c12 ),
    .o({\PWME/sub1/c13 ,\PWME/n26 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub1/u13  (
    .a(pnumcntE[13]),
    .b(1'b0),
    .c(\PWME/sub1/c13 ),
    .o({\PWME/sub1/c14 ,\PWME/n26 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub1/u14  (
    .a(pnumcntE[14]),
    .b(1'b0),
    .c(\PWME/sub1/c14 ),
    .o({\PWME/sub1/c15 ,\PWME/n26 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub1/u15  (
    .a(pnumcntE[15]),
    .b(1'b0),
    .c(\PWME/sub1/c15 ),
    .o({\PWME/sub1/c16 ,\PWME/n26 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub1/u16  (
    .a(pnumcntE[16]),
    .b(1'b0),
    .c(\PWME/sub1/c16 ),
    .o({\PWME/sub1/c17 ,\PWME/n26 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub1/u17  (
    .a(pnumcntE[17]),
    .b(1'b0),
    .c(\PWME/sub1/c17 ),
    .o({\PWME/sub1/c18 ,\PWME/n26 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub1/u18  (
    .a(pnumcntE[18]),
    .b(1'b0),
    .c(\PWME/sub1/c18 ),
    .o({\PWME/sub1/c19 ,\PWME/n26 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub1/u19  (
    .a(pnumcntE[19]),
    .b(1'b0),
    .c(\PWME/sub1/c19 ),
    .o({\PWME/sub1/c20 ,\PWME/n26 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub1/u2  (
    .a(pnumcntE[2]),
    .b(1'b0),
    .c(\PWME/sub1/c2 ),
    .o({\PWME/sub1/c3 ,\PWME/n26 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub1/u20  (
    .a(pnumcntE[20]),
    .b(1'b0),
    .c(\PWME/sub1/c20 ),
    .o({\PWME/sub1/c21 ,\PWME/n26 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub1/u21  (
    .a(pnumcntE[21]),
    .b(1'b0),
    .c(\PWME/sub1/c21 ),
    .o({\PWME/sub1/c22 ,\PWME/n26 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub1/u22  (
    .a(pnumcntE[22]),
    .b(1'b0),
    .c(\PWME/sub1/c22 ),
    .o({\PWME/sub1/c23 ,\PWME/n26 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub1/u23  (
    .a(pnumcntE[23]),
    .b(1'b0),
    .c(\PWME/sub1/c23 ),
    .o({open_n116,\PWME/n26 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub1/u3  (
    .a(pnumcntE[3]),
    .b(1'b0),
    .c(\PWME/sub1/c3 ),
    .o({\PWME/sub1/c4 ,\PWME/n26 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub1/u4  (
    .a(pnumcntE[4]),
    .b(1'b0),
    .c(\PWME/sub1/c4 ),
    .o({\PWME/sub1/c5 ,\PWME/n26 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub1/u5  (
    .a(pnumcntE[5]),
    .b(1'b0),
    .c(\PWME/sub1/c5 ),
    .o({\PWME/sub1/c6 ,\PWME/n26 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub1/u6  (
    .a(pnumcntE[6]),
    .b(1'b0),
    .c(\PWME/sub1/c6 ),
    .o({\PWME/sub1/c7 ,\PWME/n26 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub1/u7  (
    .a(pnumcntE[7]),
    .b(1'b0),
    .c(\PWME/sub1/c7 ),
    .o({\PWME/sub1/c8 ,\PWME/n26 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub1/u8  (
    .a(pnumcntE[8]),
    .b(1'b0),
    .c(\PWME/sub1/c8 ),
    .o({\PWME/sub1/c9 ,\PWME/n26 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWME/sub1/u9  (
    .a(pnumcntE[9]),
    .b(1'b0),
    .c(\PWME/sub1/c9 ),
    .o({\PWME/sub1/c10 ,\PWME/n26 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \PWME/sub1/ucin  (
    .a(1'b0),
    .o({\PWME/sub1/c0 ,open_n119}));
  reg_ar_as_w1 \PWMF/State_reg  (
    .clk(clk100m),
    .d(\PWMF/n10 ),
    .en(1'b1),
    .reset(~rstn),
    .set(1'b0),
    .q(pwm_state_read[15]));  // src/OnePWM.v(26)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[0]  (
    .i(\PWMF/RemaTxNum[0]_keep ),
    .o(pnumcntF[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[10]  (
    .i(\PWMF/RemaTxNum[10]_keep ),
    .o(pnumcntF[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[11]  (
    .i(\PWMF/RemaTxNum[11]_keep ),
    .o(pnumcntF[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[12]  (
    .i(\PWMF/RemaTxNum[12]_keep ),
    .o(pnumcntF[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[13]  (
    .i(\PWMF/RemaTxNum[13]_keep ),
    .o(pnumcntF[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[14]  (
    .i(\PWMF/RemaTxNum[14]_keep ),
    .o(pnumcntF[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[15]  (
    .i(\PWMF/RemaTxNum[15]_keep ),
    .o(pnumcntF[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[16]  (
    .i(\PWMF/RemaTxNum[16]_keep ),
    .o(pnumcntF[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[17]  (
    .i(\PWMF/RemaTxNum[17]_keep ),
    .o(pnumcntF[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[18]  (
    .i(\PWMF/RemaTxNum[18]_keep ),
    .o(pnumcntF[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[19]  (
    .i(\PWMF/RemaTxNum[19]_keep ),
    .o(pnumcntF[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[1]  (
    .i(\PWMF/RemaTxNum[1]_keep ),
    .o(pnumcntF[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[20]  (
    .i(\PWMF/RemaTxNum[20]_keep ),
    .o(pnumcntF[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[21]  (
    .i(\PWMF/RemaTxNum[21]_keep ),
    .o(pnumcntF[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[22]  (
    .i(\PWMF/RemaTxNum[22]_keep ),
    .o(pnumcntF[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[23]  (
    .i(\PWMF/RemaTxNum[23]_keep ),
    .o(pnumcntF[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[2]  (
    .i(\PWMF/RemaTxNum[2]_keep ),
    .o(pnumcntF[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[3]  (
    .i(\PWMF/RemaTxNum[3]_keep ),
    .o(pnumcntF[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[4]  (
    .i(\PWMF/RemaTxNum[4]_keep ),
    .o(pnumcntF[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[5]  (
    .i(\PWMF/RemaTxNum[5]_keep ),
    .o(pnumcntF[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[6]  (
    .i(\PWMF/RemaTxNum[6]_keep ),
    .o(pnumcntF[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[7]  (
    .i(\PWMF/RemaTxNum[7]_keep ),
    .o(pnumcntF[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[8]  (
    .i(\PWMF/RemaTxNum[8]_keep ),
    .o(pnumcntF[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[9]  (
    .i(\PWMF/RemaTxNum[9]_keep ),
    .o(pnumcntF[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_dir  (
    .i(\PWMF/dir_keep ),
    .o(dir_pad[15]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[0]  (
    .i(\PWMF/pnumr[0]_keep ),
    .o(\PWMF/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[10]  (
    .i(\PWMF/pnumr[10]_keep ),
    .o(\PWMF/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[11]  (
    .i(\PWMF/pnumr[11]_keep ),
    .o(\PWMF/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[12]  (
    .i(\PWMF/pnumr[12]_keep ),
    .o(\PWMF/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[13]  (
    .i(\PWMF/pnumr[13]_keep ),
    .o(\PWMF/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[14]  (
    .i(\PWMF/pnumr[14]_keep ),
    .o(\PWMF/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[15]  (
    .i(\PWMF/pnumr[15]_keep ),
    .o(\PWMF/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[16]  (
    .i(\PWMF/pnumr[16]_keep ),
    .o(\PWMF/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[17]  (
    .i(\PWMF/pnumr[17]_keep ),
    .o(\PWMF/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[18]  (
    .i(\PWMF/pnumr[18]_keep ),
    .o(\PWMF/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[19]  (
    .i(\PWMF/pnumr[19]_keep ),
    .o(\PWMF/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[1]  (
    .i(\PWMF/pnumr[1]_keep ),
    .o(\PWMF/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[20]  (
    .i(\PWMF/pnumr[20]_keep ),
    .o(\PWMF/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[21]  (
    .i(\PWMF/pnumr[21]_keep ),
    .o(\PWMF/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[22]  (
    .i(\PWMF/pnumr[22]_keep ),
    .o(\PWMF/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[23]  (
    .i(\PWMF/pnumr[23]_keep ),
    .o(\PWMF/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[24]  (
    .i(\PWMF/pnumr[24]_keep ),
    .o(\PWMF/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[25]  (
    .i(\PWMF/pnumr[25]_keep ),
    .o(\PWMF/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[26]  (
    .i(\PWMF/pnumr[26]_keep ),
    .o(\PWMF/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[27]  (
    .i(\PWMF/pnumr[27]_keep ),
    .o(\PWMF/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[28]  (
    .i(\PWMF/pnumr[28]_keep ),
    .o(\PWMF/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[29]  (
    .i(\PWMF/pnumr[29]_keep ),
    .o(\PWMF/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[2]  (
    .i(\PWMF/pnumr[2]_keep ),
    .o(\PWMF/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[30]  (
    .i(\PWMF/pnumr[30]_keep ),
    .o(\PWMF/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[31]  (
    .i(\PWMF/pnumr[31]_keep ),
    .o(\PWMF/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[3]  (
    .i(\PWMF/pnumr[3]_keep ),
    .o(\PWMF/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[4]  (
    .i(\PWMF/pnumr[4]_keep ),
    .o(\PWMF/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[5]  (
    .i(\PWMF/pnumr[5]_keep ),
    .o(\PWMF/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[6]  (
    .i(\PWMF/pnumr[6]_keep ),
    .o(\PWMF/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[7]  (
    .i(\PWMF/pnumr[7]_keep ),
    .o(\PWMF/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[8]  (
    .i(\PWMF/pnumr[8]_keep ),
    .o(\PWMF/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[9]  (
    .i(\PWMF/pnumr[9]_keep ),
    .o(\PWMF/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pwm  (
    .i(\PWMF/pwm_keep ),
    .o(pwm_pad[15]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_stopreq  (
    .i(\PWMF/stopreq_keep ),
    .o(\PWMF/stopreq ));  // src/OnePWM.v(14)
  reg_ar_as_w1 \PWMF/dir_reg  (
    .clk(clk100m),
    .d(\PWMF/n32 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/dir_keep ));  // src/OnePWM.v(58)
  reg_sr_as_w1 \PWMF/pwm_reg  (
    .clk(clk100m),
    .d(\pwm[15]_d ),
    .en(1'b1),
    .reset(~\PWMF/u14_sel_is_1_o ),
    .set(1'b0),
    .q(\PWMF/pwm_keep ));  // src/OnePWM.v(45)
  reg_sr_as_w1 \PWMF/reg0_b0  (
    .clk(clk100m),
    .d(\PWMF/n13 [0]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [0]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b1  (
    .clk(clk100m),
    .d(\PWMF/n13 [1]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [1]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b10  (
    .clk(clk100m),
    .d(\PWMF/n13 [10]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [10]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b11  (
    .clk(clk100m),
    .d(\PWMF/n13 [11]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [11]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b12  (
    .clk(clk100m),
    .d(\PWMF/n13 [12]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [12]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b13  (
    .clk(clk100m),
    .d(\PWMF/n13 [13]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [13]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b14  (
    .clk(clk100m),
    .d(\PWMF/n13 [14]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [14]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b15  (
    .clk(clk100m),
    .d(\PWMF/n13 [15]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [15]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b16  (
    .clk(clk100m),
    .d(\PWMF/n13 [16]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [16]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b17  (
    .clk(clk100m),
    .d(\PWMF/n13 [17]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [17]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b18  (
    .clk(clk100m),
    .d(\PWMF/n13 [18]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [18]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b19  (
    .clk(clk100m),
    .d(\PWMF/n13 [19]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [19]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b2  (
    .clk(clk100m),
    .d(\PWMF/n13 [2]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [2]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b20  (
    .clk(clk100m),
    .d(\PWMF/n13 [20]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [20]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b21  (
    .clk(clk100m),
    .d(\PWMF/n13 [21]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [21]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b22  (
    .clk(clk100m),
    .d(\PWMF/n13 [22]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [22]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b23  (
    .clk(clk100m),
    .d(\PWMF/n13 [23]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [23]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b24  (
    .clk(clk100m),
    .d(\PWMF/n13 [24]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [24]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b25  (
    .clk(clk100m),
    .d(\PWMF/n13 [25]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [25]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b26  (
    .clk(clk100m),
    .d(\PWMF/n13 [26]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [26]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b3  (
    .clk(clk100m),
    .d(\PWMF/n13 [3]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [3]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b4  (
    .clk(clk100m),
    .d(\PWMF/n13 [4]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [4]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b5  (
    .clk(clk100m),
    .d(\PWMF/n13 [5]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [5]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b6  (
    .clk(clk100m),
    .d(\PWMF/n13 [6]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [6]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b7  (
    .clk(clk100m),
    .d(\PWMF/n13 [7]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [7]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b8  (
    .clk(clk100m),
    .d(\PWMF/n13 [8]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [8]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b9  (
    .clk(clk100m),
    .d(\PWMF/n13 [9]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b0  (
    .clk(clk100m),
    .d(freqF[0]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [0]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b1  (
    .clk(clk100m),
    .d(freqF[1]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [1]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b10  (
    .clk(clk100m),
    .d(freqF[10]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [10]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b11  (
    .clk(clk100m),
    .d(freqF[11]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [11]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b12  (
    .clk(clk100m),
    .d(freqF[12]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [12]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b13  (
    .clk(clk100m),
    .d(freqF[13]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [13]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b14  (
    .clk(clk100m),
    .d(freqF[14]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [14]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b15  (
    .clk(clk100m),
    .d(freqF[15]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [15]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b16  (
    .clk(clk100m),
    .d(freqF[16]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [16]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b17  (
    .clk(clk100m),
    .d(freqF[17]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [17]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b18  (
    .clk(clk100m),
    .d(freqF[18]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [18]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b19  (
    .clk(clk100m),
    .d(freqF[19]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [19]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b2  (
    .clk(clk100m),
    .d(freqF[2]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [2]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b20  (
    .clk(clk100m),
    .d(freqF[20]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [20]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b21  (
    .clk(clk100m),
    .d(freqF[21]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [21]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b22  (
    .clk(clk100m),
    .d(freqF[22]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [22]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b23  (
    .clk(clk100m),
    .d(freqF[23]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [23]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b24  (
    .clk(clk100m),
    .d(freqF[24]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [24]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b25  (
    .clk(clk100m),
    .d(freqF[25]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [25]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b26  (
    .clk(clk100m),
    .d(freqF[26]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [26]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b3  (
    .clk(clk100m),
    .d(freqF[3]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [3]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b4  (
    .clk(clk100m),
    .d(freqF[4]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [4]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b5  (
    .clk(clk100m),
    .d(freqF[5]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [5]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b6  (
    .clk(clk100m),
    .d(freqF[6]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [6]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b7  (
    .clk(clk100m),
    .d(freqF[7]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [7]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b8  (
    .clk(clk100m),
    .d(freqF[8]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [8]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b9  (
    .clk(clk100m),
    .d(freqF[9]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg2_b0  (
    .clk(clk100m),
    .d(\PWMF/n23 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[0]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b1  (
    .clk(clk100m),
    .d(\PWMF/n23 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[1]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b10  (
    .clk(clk100m),
    .d(\PWMF/n23 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[10]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b11  (
    .clk(clk100m),
    .d(\PWMF/n23 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[11]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b12  (
    .clk(clk100m),
    .d(\PWMF/n23 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[12]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b13  (
    .clk(clk100m),
    .d(\PWMF/n23 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[13]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b14  (
    .clk(clk100m),
    .d(\PWMF/n23 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[14]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b15  (
    .clk(clk100m),
    .d(\PWMF/n23 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[15]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b16  (
    .clk(clk100m),
    .d(\PWMF/n23 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[16]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b17  (
    .clk(clk100m),
    .d(\PWMF/n23 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[17]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b18  (
    .clk(clk100m),
    .d(\PWMF/n23 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[18]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b19  (
    .clk(clk100m),
    .d(\PWMF/n23 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[19]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b2  (
    .clk(clk100m),
    .d(\PWMF/n23 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[2]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b20  (
    .clk(clk100m),
    .d(\PWMF/n23 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[20]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b21  (
    .clk(clk100m),
    .d(\PWMF/n23 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[21]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b22  (
    .clk(clk100m),
    .d(\PWMF/n23 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[22]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b23  (
    .clk(clk100m),
    .d(\PWMF/n23 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[23]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b24  (
    .clk(clk100m),
    .d(\PWMF/n23 [24]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[24]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b25  (
    .clk(clk100m),
    .d(\PWMF/n23 [25]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[25]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b26  (
    .clk(clk100m),
    .d(\PWMF/n23 [26]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[26]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b27  (
    .clk(clk100m),
    .d(\PWMF/n23 [27]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[27]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b28  (
    .clk(clk100m),
    .d(\PWMF/n23 [28]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[28]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b29  (
    .clk(clk100m),
    .d(\PWMF/n23 [29]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[29]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b3  (
    .clk(clk100m),
    .d(\PWMF/n23 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[3]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b30  (
    .clk(clk100m),
    .d(\PWMF/n23 [30]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[30]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b31  (
    .clk(clk100m),
    .d(\PWMF/n23 [31]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[31]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b4  (
    .clk(clk100m),
    .d(\PWMF/n23 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[4]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b5  (
    .clk(clk100m),
    .d(\PWMF/n23 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[5]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b6  (
    .clk(clk100m),
    .d(\PWMF/n23 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[6]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b7  (
    .clk(clk100m),
    .d(\PWMF/n23 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[7]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b8  (
    .clk(clk100m),
    .d(\PWMF/n23 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[8]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b9  (
    .clk(clk100m),
    .d(\PWMF/n23 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[9]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg3_b0  (
    .clk(clk100m),
    .d(\PWMF/n31 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[0]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b1  (
    .clk(clk100m),
    .d(\PWMF/n31 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[1]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b10  (
    .clk(clk100m),
    .d(\PWMF/n31 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[10]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b11  (
    .clk(clk100m),
    .d(\PWMF/n31 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[11]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b12  (
    .clk(clk100m),
    .d(\PWMF/n31 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[12]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b13  (
    .clk(clk100m),
    .d(\PWMF/n31 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[13]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b14  (
    .clk(clk100m),
    .d(\PWMF/n31 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[14]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b15  (
    .clk(clk100m),
    .d(\PWMF/n31 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[15]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b16  (
    .clk(clk100m),
    .d(\PWMF/n31 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[16]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b17  (
    .clk(clk100m),
    .d(\PWMF/n31 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[17]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b18  (
    .clk(clk100m),
    .d(\PWMF/n31 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[18]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b19  (
    .clk(clk100m),
    .d(\PWMF/n31 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[19]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b2  (
    .clk(clk100m),
    .d(\PWMF/n31 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[2]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b20  (
    .clk(clk100m),
    .d(\PWMF/n31 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[20]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b21  (
    .clk(clk100m),
    .d(\PWMF/n31 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[21]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b22  (
    .clk(clk100m),
    .d(\PWMF/n31 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[22]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b23  (
    .clk(clk100m),
    .d(\PWMF/n31 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[23]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b3  (
    .clk(clk100m),
    .d(\PWMF/n31 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[3]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b4  (
    .clk(clk100m),
    .d(\PWMF/n31 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[4]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b5  (
    .clk(clk100m),
    .d(\PWMF/n31 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[5]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b6  (
    .clk(clk100m),
    .d(\PWMF/n31 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[6]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b7  (
    .clk(clk100m),
    .d(\PWMF/n31 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[7]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b8  (
    .clk(clk100m),
    .d(\PWMF/n31 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[8]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b9  (
    .clk(clk100m),
    .d(\PWMF/n31 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[9]_keep ));  // src/OnePWM.v(58)
  reg_ar_ss_w1 \PWMF/stopreq_reg  (
    .clk(clk100m),
    .d(\PWMF/n1 ),
    .en(1'b1),
    .reset(1'b0),
    .set(pwm_start_stop[15]),
    .q(\PWMF/stopreq_keep ));  // src/OnePWM.v(15)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub0/u0  (
    .a(\PWMF/FreCnt [0]),
    .b(1'b1),
    .c(\PWMF/sub0/c0 ),
    .o({\PWMF/sub0/c1 ,\PWMF/n12 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub0/u1  (
    .a(\PWMF/FreCnt [1]),
    .b(1'b0),
    .c(\PWMF/sub0/c1 ),
    .o({\PWMF/sub0/c2 ,\PWMF/n12 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub0/u10  (
    .a(\PWMF/FreCnt [10]),
    .b(1'b0),
    .c(\PWMF/sub0/c10 ),
    .o({\PWMF/sub0/c11 ,\PWMF/n12 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub0/u11  (
    .a(\PWMF/FreCnt [11]),
    .b(1'b0),
    .c(\PWMF/sub0/c11 ),
    .o({\PWMF/sub0/c12 ,\PWMF/n12 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub0/u12  (
    .a(\PWMF/FreCnt [12]),
    .b(1'b0),
    .c(\PWMF/sub0/c12 ),
    .o({\PWMF/sub0/c13 ,\PWMF/n12 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub0/u13  (
    .a(\PWMF/FreCnt [13]),
    .b(1'b0),
    .c(\PWMF/sub0/c13 ),
    .o({\PWMF/sub0/c14 ,\PWMF/n12 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub0/u14  (
    .a(\PWMF/FreCnt [14]),
    .b(1'b0),
    .c(\PWMF/sub0/c14 ),
    .o({\PWMF/sub0/c15 ,\PWMF/n12 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub0/u15  (
    .a(\PWMF/FreCnt [15]),
    .b(1'b0),
    .c(\PWMF/sub0/c15 ),
    .o({\PWMF/sub0/c16 ,\PWMF/n12 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub0/u16  (
    .a(\PWMF/FreCnt [16]),
    .b(1'b0),
    .c(\PWMF/sub0/c16 ),
    .o({\PWMF/sub0/c17 ,\PWMF/n12 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub0/u17  (
    .a(\PWMF/FreCnt [17]),
    .b(1'b0),
    .c(\PWMF/sub0/c17 ),
    .o({\PWMF/sub0/c18 ,\PWMF/n12 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub0/u18  (
    .a(\PWMF/FreCnt [18]),
    .b(1'b0),
    .c(\PWMF/sub0/c18 ),
    .o({\PWMF/sub0/c19 ,\PWMF/n12 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub0/u19  (
    .a(\PWMF/FreCnt [19]),
    .b(1'b0),
    .c(\PWMF/sub0/c19 ),
    .o({\PWMF/sub0/c20 ,\PWMF/n12 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub0/u2  (
    .a(\PWMF/FreCnt [2]),
    .b(1'b0),
    .c(\PWMF/sub0/c2 ),
    .o({\PWMF/sub0/c3 ,\PWMF/n12 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub0/u20  (
    .a(\PWMF/FreCnt [20]),
    .b(1'b0),
    .c(\PWMF/sub0/c20 ),
    .o({\PWMF/sub0/c21 ,\PWMF/n12 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub0/u21  (
    .a(\PWMF/FreCnt [21]),
    .b(1'b0),
    .c(\PWMF/sub0/c21 ),
    .o({\PWMF/sub0/c22 ,\PWMF/n12 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub0/u22  (
    .a(\PWMF/FreCnt [22]),
    .b(1'b0),
    .c(\PWMF/sub0/c22 ),
    .o({\PWMF/sub0/c23 ,\PWMF/n12 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub0/u23  (
    .a(\PWMF/FreCnt [23]),
    .b(1'b0),
    .c(\PWMF/sub0/c23 ),
    .o({\PWMF/sub0/c24 ,\PWMF/n12 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub0/u24  (
    .a(\PWMF/FreCnt [24]),
    .b(1'b0),
    .c(\PWMF/sub0/c24 ),
    .o({\PWMF/sub0/c25 ,\PWMF/n12 [24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub0/u25  (
    .a(\PWMF/FreCnt [25]),
    .b(1'b0),
    .c(\PWMF/sub0/c25 ),
    .o({\PWMF/sub0/c26 ,\PWMF/n12 [25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub0/u26  (
    .a(\PWMF/FreCnt [26]),
    .b(1'b0),
    .c(\PWMF/sub0/c26 ),
    .o({open_n120,\PWMF/n12 [26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub0/u3  (
    .a(\PWMF/FreCnt [3]),
    .b(1'b0),
    .c(\PWMF/sub0/c3 ),
    .o({\PWMF/sub0/c4 ,\PWMF/n12 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub0/u4  (
    .a(\PWMF/FreCnt [4]),
    .b(1'b0),
    .c(\PWMF/sub0/c4 ),
    .o({\PWMF/sub0/c5 ,\PWMF/n12 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub0/u5  (
    .a(\PWMF/FreCnt [5]),
    .b(1'b0),
    .c(\PWMF/sub0/c5 ),
    .o({\PWMF/sub0/c6 ,\PWMF/n12 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub0/u6  (
    .a(\PWMF/FreCnt [6]),
    .b(1'b0),
    .c(\PWMF/sub0/c6 ),
    .o({\PWMF/sub0/c7 ,\PWMF/n12 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub0/u7  (
    .a(\PWMF/FreCnt [7]),
    .b(1'b0),
    .c(\PWMF/sub0/c7 ),
    .o({\PWMF/sub0/c8 ,\PWMF/n12 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub0/u8  (
    .a(\PWMF/FreCnt [8]),
    .b(1'b0),
    .c(\PWMF/sub0/c8 ),
    .o({\PWMF/sub0/c9 ,\PWMF/n12 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub0/u9  (
    .a(\PWMF/FreCnt [9]),
    .b(1'b0),
    .c(\PWMF/sub0/c9 ),
    .o({\PWMF/sub0/c10 ,\PWMF/n12 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \PWMF/sub0/ucin  (
    .a(1'b0),
    .o({\PWMF/sub0/c0 ,open_n123}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub1/u0  (
    .a(pnumcntF[0]),
    .b(1'b1),
    .c(\PWMF/sub1/c0 ),
    .o({\PWMF/sub1/c1 ,\PWMF/n26 [0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub1/u1  (
    .a(pnumcntF[1]),
    .b(1'b0),
    .c(\PWMF/sub1/c1 ),
    .o({\PWMF/sub1/c2 ,\PWMF/n26 [1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub1/u10  (
    .a(pnumcntF[10]),
    .b(1'b0),
    .c(\PWMF/sub1/c10 ),
    .o({\PWMF/sub1/c11 ,\PWMF/n26 [10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub1/u11  (
    .a(pnumcntF[11]),
    .b(1'b0),
    .c(\PWMF/sub1/c11 ),
    .o({\PWMF/sub1/c12 ,\PWMF/n26 [11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub1/u12  (
    .a(pnumcntF[12]),
    .b(1'b0),
    .c(\PWMF/sub1/c12 ),
    .o({\PWMF/sub1/c13 ,\PWMF/n26 [12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub1/u13  (
    .a(pnumcntF[13]),
    .b(1'b0),
    .c(\PWMF/sub1/c13 ),
    .o({\PWMF/sub1/c14 ,\PWMF/n26 [13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub1/u14  (
    .a(pnumcntF[14]),
    .b(1'b0),
    .c(\PWMF/sub1/c14 ),
    .o({\PWMF/sub1/c15 ,\PWMF/n26 [14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub1/u15  (
    .a(pnumcntF[15]),
    .b(1'b0),
    .c(\PWMF/sub1/c15 ),
    .o({\PWMF/sub1/c16 ,\PWMF/n26 [15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub1/u16  (
    .a(pnumcntF[16]),
    .b(1'b0),
    .c(\PWMF/sub1/c16 ),
    .o({\PWMF/sub1/c17 ,\PWMF/n26 [16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub1/u17  (
    .a(pnumcntF[17]),
    .b(1'b0),
    .c(\PWMF/sub1/c17 ),
    .o({\PWMF/sub1/c18 ,\PWMF/n26 [17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub1/u18  (
    .a(pnumcntF[18]),
    .b(1'b0),
    .c(\PWMF/sub1/c18 ),
    .o({\PWMF/sub1/c19 ,\PWMF/n26 [18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub1/u19  (
    .a(pnumcntF[19]),
    .b(1'b0),
    .c(\PWMF/sub1/c19 ),
    .o({\PWMF/sub1/c20 ,\PWMF/n26 [19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub1/u2  (
    .a(pnumcntF[2]),
    .b(1'b0),
    .c(\PWMF/sub1/c2 ),
    .o({\PWMF/sub1/c3 ,\PWMF/n26 [2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub1/u20  (
    .a(pnumcntF[20]),
    .b(1'b0),
    .c(\PWMF/sub1/c20 ),
    .o({\PWMF/sub1/c21 ,\PWMF/n26 [20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub1/u21  (
    .a(pnumcntF[21]),
    .b(1'b0),
    .c(\PWMF/sub1/c21 ),
    .o({\PWMF/sub1/c22 ,\PWMF/n26 [21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub1/u22  (
    .a(pnumcntF[22]),
    .b(1'b0),
    .c(\PWMF/sub1/c22 ),
    .o({\PWMF/sub1/c23 ,\PWMF/n26 [22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub1/u23  (
    .a(pnumcntF[23]),
    .b(1'b0),
    .c(\PWMF/sub1/c23 ),
    .o({open_n124,\PWMF/n26 [23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub1/u3  (
    .a(pnumcntF[3]),
    .b(1'b0),
    .c(\PWMF/sub1/c3 ),
    .o({\PWMF/sub1/c4 ,\PWMF/n26 [3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub1/u4  (
    .a(pnumcntF[4]),
    .b(1'b0),
    .c(\PWMF/sub1/c4 ),
    .o({\PWMF/sub1/c5 ,\PWMF/n26 [4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub1/u5  (
    .a(pnumcntF[5]),
    .b(1'b0),
    .c(\PWMF/sub1/c5 ),
    .o({\PWMF/sub1/c6 ,\PWMF/n26 [5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub1/u6  (
    .a(pnumcntF[6]),
    .b(1'b0),
    .c(\PWMF/sub1/c6 ),
    .o({\PWMF/sub1/c7 ,\PWMF/n26 [6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub1/u7  (
    .a(pnumcntF[7]),
    .b(1'b0),
    .c(\PWMF/sub1/c7 ),
    .o({\PWMF/sub1/c8 ,\PWMF/n26 [7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub1/u8  (
    .a(pnumcntF[8]),
    .b(1'b0),
    .c(\PWMF/sub1/c8 ),
    .o({\PWMF/sub1/c9 ,\PWMF/n26 [8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \PWMF/sub1/u9  (
    .a(pnumcntF[9]),
    .b(1'b0),
    .c(\PWMF/sub1/c9 ),
    .o({\PWMF/sub1/c10 ,\PWMF/n26 [9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \PWMF/sub1/ucin  (
    .a(1'b0),
    .o({\PWMF/sub1/c0 ,open_n127}));
  EF2_PHY_MCU #(
    .GPIO_L0("ENABLE"),
    .GPIO_L1("ENABLE"),
    .GPIO_L10("DISABLE"),
    .GPIO_L11("DISABLE"),
    .GPIO_L12("DISABLE"),
    .GPIO_L13("DISABLE"),
    .GPIO_L14("DISABLE"),
    .GPIO_L15("DISABLE"),
    .GPIO_L2("DISABLE"),
    .GPIO_L3("DISABLE"),
    .GPIO_L4("DISABLE"),
    .GPIO_L5("DISABLE"),
    .GPIO_L6("DISABLE"),
    .GPIO_L7("DISABLE"),
    .GPIO_L8("ENABLE"),
    .GPIO_L9("ENABLE"))
    \U_AHB/M3WithAHB/mcu_inst  (
    .gpio_h_in(16'b0000000000000000),
    .h2h_hrdata(\U_AHB/h2h_hrdata ),
    .h2h_hreadyout(1'b1),
    .h2h_hresp(2'b00),
    .h2h_mclk(clk100m),
    .h2h_rstn(rstn),
    .ppm_clk(clk25m),
    .h2h_haddr({open_n171,open_n172,open_n173,open_n174,open_n175,open_n176,open_n177,open_n178,open_n179,open_n180,open_n181,open_n182,open_n183,open_n184,open_n185,open_n186,open_n187,\U_AHB/h2h_haddrw [14:2],open_n188,open_n189}),
    .h2h_hwdata(\U_AHB/h2h_hwdata ),
    .h2h_hwrite(\U_AHB/h2h_hwritew ));  // al_ip/M3WithAHB.v(46)
  reg_ar_as_w1 \U_AHB/h2h_hwrite_reg  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwritew ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hwrite ));  // src/AHB.v(24)
  reg_ar_as_w1 \U_AHB/reg0_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_haddrw [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_haddr [2]));  // src/AHB.v(25)
  reg_ar_as_w1 \U_AHB/reg0_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_haddrw [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_haddr [3]));  // src/AHB.v(25)
  reg_ar_as_w1 \U_AHB/reg0_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_haddrw [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_haddr [12]));  // src/AHB.v(25)
  reg_ar_as_w1 \U_AHB/reg0_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_haddrw [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_haddr [13]));  // src/AHB.v(25)
  reg_ar_as_w1 \U_AHB/reg0_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_haddrw [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_haddr [14]));  // src/AHB.v(25)
  reg_ar_as_w1 \U_AHB/reg0_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_haddrw [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_haddr [4]));  // src/AHB.v(25)
  reg_ar_as_w1 \U_AHB/reg0_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_haddrw [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_haddr [5]));  // src/AHB.v(25)
  reg_ar_as_w1 \U_AHB/reg0_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_haddrw [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_haddr [6]));  // src/AHB.v(25)
  reg_ar_as_w1 \U_AHB/reg0_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_haddrw [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_haddr [7]));  // src/AHB.v(25)
  reg_ar_as_w1 \U_AHB/reg0_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_haddrw [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_haddr [8]));  // src/AHB.v(25)
  reg_ar_as_w1 \U_AHB/reg0_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_haddrw [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_haddr [9]));  // src/AHB.v(25)
  reg_ar_as_w1 \U_AHB/reg0_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_haddrw [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_haddr [10]));  // src/AHB.v(25)
  reg_ar_as_w1 \U_AHB/reg0_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_haddrw [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_haddr [11]));  // src/AHB.v(25)
  reg_ar_as_w1 \U_AHB/reg10_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[0]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[1]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[10]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[11]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[12]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[13]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[14]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[15]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[16]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[17]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[18]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[19]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[2]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[20]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[21]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[22]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[23]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[24]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[25]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[26]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[3]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[4]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[5]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[6]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[7]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[8]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[9]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg11_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[0]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[1]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[10]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[11]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[12]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[13]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[14]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[15]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[16]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[17]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[18]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[19]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[2]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[20]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[21]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[22]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[23]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[24]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[25]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[26]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[3]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[4]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[5]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[6]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[7]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[8]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[9]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg12_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[0]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[1]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[10]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[11]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[12]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[13]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[14]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[15]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[16]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[17]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[18]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[19]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[2]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[20]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[21]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[22]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[23]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[24]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[25]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[26]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[3]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[4]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[5]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[6]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[7]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[8]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[9]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg13_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[0]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[1]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[10]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[11]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[12]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[13]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[14]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[15]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[16]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[17]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[18]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[19]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[2]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[20]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[21]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[22]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[23]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[24]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[25]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[26]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[3]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[4]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[5]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[6]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[7]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[8]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[9]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg14_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[0]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[1]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[10]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[11]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[12]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[13]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[14]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[15]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[16]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[17]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[18]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[19]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[2]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[20]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[21]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[22]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[23]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[24]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[25]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[26]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[3]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[4]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[5]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[6]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[7]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[8]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[9]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg15_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[0]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[1]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[10]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[11]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[12]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[13]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[14]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[15]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[16]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[17]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[18]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[19]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[2]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[20]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[21]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[22]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[23]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[24]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[25]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[26]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[3]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[4]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[5]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[6]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[7]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[8]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[9]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg16_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[0]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[1]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[10]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[11]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[12]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[13]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[14]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[15]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[16]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[17]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[18]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[19]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[2]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[20]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[21]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[22]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[23]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[24]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[25]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[26]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[3]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[4]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[5]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[6]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[7]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[8]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[9]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg17_b0  (
    .clk(clk100m),
    .d(\U_AHB/n42 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out_pad[0]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b1  (
    .clk(clk100m),
    .d(\U_AHB/n42 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out_pad[1]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b10  (
    .clk(clk100m),
    .d(\U_AHB/n42 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out_pad[10]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b11  (
    .clk(clk100m),
    .d(\U_AHB/n42 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out_pad[11]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b12  (
    .clk(clk100m),
    .d(\U_AHB/n42 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out_pad[12]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b13  (
    .clk(clk100m),
    .d(\U_AHB/n42 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out_pad[13]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b14  (
    .clk(clk100m),
    .d(\U_AHB/n42 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out_pad[14]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b15  (
    .clk(clk100m),
    .d(\U_AHB/n42 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out_pad[15]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b16  (
    .clk(clk100m),
    .d(\U_AHB/n42 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out_pad[16]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b17  (
    .clk(clk100m),
    .d(\U_AHB/n42 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out_pad[17]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b18  (
    .clk(clk100m),
    .d(\U_AHB/n42 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out_pad[18]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b19  (
    .clk(clk100m),
    .d(\U_AHB/n42 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out_pad[19]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b2  (
    .clk(clk100m),
    .d(\U_AHB/n42 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out_pad[2]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b20  (
    .clk(clk100m),
    .d(\U_AHB/n42 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out_pad[20]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b21  (
    .clk(clk100m),
    .d(\U_AHB/n42 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out_pad[21]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b22  (
    .clk(clk100m),
    .d(\U_AHB/n42 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out_pad[22]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b23  (
    .clk(clk100m),
    .d(\U_AHB/n42 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out_pad[23]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b24  (
    .clk(clk100m),
    .d(\U_AHB/n42 [24]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out_pad[24]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b25  (
    .clk(clk100m),
    .d(\U_AHB/n42 [25]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out_pad[25]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b26  (
    .clk(clk100m),
    .d(\U_AHB/n42 [26]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out_pad[26]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b27  (
    .clk(clk100m),
    .d(\U_AHB/n42 [27]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out_pad[27]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b28  (
    .clk(clk100m),
    .d(\U_AHB/n42 [28]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out_pad[28]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b29  (
    .clk(clk100m),
    .d(\U_AHB/n42 [29]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out_pad[29]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b3  (
    .clk(clk100m),
    .d(\U_AHB/n42 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out_pad[3]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b30  (
    .clk(clk100m),
    .d(\U_AHB/n42 [30]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out_pad[30]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b31  (
    .clk(clk100m),
    .d(\U_AHB/n42 [31]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out_pad[31]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b4  (
    .clk(clk100m),
    .d(\U_AHB/n42 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out_pad[4]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b5  (
    .clk(clk100m),
    .d(\U_AHB/n42 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out_pad[5]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b6  (
    .clk(clk100m),
    .d(\U_AHB/n42 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out_pad[6]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b7  (
    .clk(clk100m),
    .d(\U_AHB/n42 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out_pad[7]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b8  (
    .clk(clk100m),
    .d(\U_AHB/n42 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out_pad[8]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b9  (
    .clk(clk100m),
    .d(\U_AHB/n42 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out_pad[9]));  // src/AHB.v(64)
  reg_sr_as_w1 \U_AHB/reg18_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[0]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[1]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[10]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[11]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[12]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[13]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[14]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[15]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[16]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[17]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[18]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[19]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[2]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[20]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[21]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[22]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[23]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[24]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[25]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[26]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b27  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [27]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[27]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b28  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [28]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[28]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b29  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [29]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[29]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[3]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b30  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [30]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[30]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b31  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [31]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[31]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b32  (
    .clk(clk100m),
    .d(1'b1),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[32]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[4]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[5]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[6]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[7]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[8]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[9]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg19_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[0]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[1]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[10]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[11]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[12]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[13]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[14]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[15]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[16]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[17]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[18]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[19]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[2]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[20]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[21]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[22]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[23]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[24]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[25]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[26]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b27  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [27]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[27]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b28  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [28]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[28]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b29  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [29]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[29]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[3]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b30  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [30]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[30]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b31  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [31]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[31]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b32  (
    .clk(clk100m),
    .d(1'b1),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[32]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[4]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[5]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[6]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[7]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[8]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[9]));  // src/AHB.v(68)
  reg_ar_as_w1 \U_AHB/reg1_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[0]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[1]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[10]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[11]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[12]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[13]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[14]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[15]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[16]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[17]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[18]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[19]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[2]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[20]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[21]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[22]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[23]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[24]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[25]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[26]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[3]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[4]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[5]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[6]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[7]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[8]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[9]));  // src/AHB.v(46)
  reg_sr_as_w1 \U_AHB/reg20_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[0]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[1]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[10]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[11]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[12]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[13]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[14]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[15]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[16]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[17]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[18]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[19]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[2]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[20]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[21]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[22]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[23]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[24]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[25]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[26]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b27  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [27]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[27]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b28  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [28]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[28]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b29  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [29]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[29]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[3]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b30  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [30]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[30]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b31  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [31]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[31]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b32  (
    .clk(clk100m),
    .d(1'b1),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[32]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[4]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[5]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[6]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[7]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[8]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[9]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg21_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[0]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[1]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[10]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[11]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[12]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[13]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[14]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[15]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[16]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[17]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[18]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[19]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[2]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[20]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[21]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[22]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[23]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[24]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[25]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[26]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b27  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [27]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[27]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b28  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [28]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[28]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b29  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [29]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[29]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[3]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b30  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [30]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[30]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b31  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [31]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[31]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b32  (
    .clk(clk100m),
    .d(1'b1),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[32]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[4]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[5]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[6]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[7]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[8]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[9]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg22_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[0]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[1]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[10]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[11]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[12]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[13]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[14]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[15]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[16]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[17]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[18]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[19]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[2]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[20]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[21]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[22]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[23]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[24]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[25]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[26]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b27  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [27]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[27]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b28  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [28]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[28]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b29  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [29]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[29]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[3]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b30  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [30]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[30]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b31  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [31]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[31]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b32  (
    .clk(clk100m),
    .d(1'b1),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[32]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[4]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[5]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[6]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[7]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[8]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[9]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg23_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[0]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[1]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[10]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[11]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[12]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[13]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[14]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[15]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[16]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[17]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[18]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[19]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[2]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[20]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[21]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[22]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[23]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[24]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[25]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[26]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b27  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [27]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[27]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b28  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [28]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[28]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b29  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [29]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[29]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[3]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b30  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [30]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[30]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b31  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [31]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[31]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b32  (
    .clk(clk100m),
    .d(1'b1),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[32]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[4]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[5]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[6]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[7]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[8]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[9]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg24_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[0]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[1]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[10]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[11]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[12]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[13]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[14]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[15]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[16]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[17]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[18]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[19]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[2]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[20]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[21]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[22]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[23]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[24]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[25]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[26]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b27  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [27]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[27]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b28  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [28]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[28]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b29  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [29]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[29]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[3]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b30  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [30]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[30]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b31  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [31]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[31]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b32  (
    .clk(clk100m),
    .d(1'b1),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[32]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[4]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[5]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[6]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[7]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[8]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[9]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg25_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[0]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[1]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[10]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[11]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[12]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[13]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[14]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[15]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[16]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[17]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[18]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[19]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[2]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[20]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[21]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[22]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[23]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[24]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[25]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[26]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b27  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [27]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[27]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b28  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [28]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[28]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b29  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [29]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[29]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[3]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b30  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [30]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[30]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b31  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [31]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[31]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b32  (
    .clk(clk100m),
    .d(1'b1),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[32]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[4]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[5]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[6]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[7]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[8]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[9]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg26_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[0]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[1]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[10]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[11]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[12]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[13]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[14]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[15]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[16]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[17]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[18]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[19]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[2]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[20]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[21]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[22]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[23]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[24]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[25]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[26]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b27  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [27]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[27]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b28  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [28]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[28]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b29  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [29]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[29]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[3]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b30  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [30]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[30]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b31  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [31]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[31]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b32  (
    .clk(clk100m),
    .d(1'b1),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[32]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[4]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[5]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[6]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[7]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[8]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[9]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg27_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[0]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[1]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[10]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[11]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[12]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[13]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[14]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[15]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[16]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[17]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[18]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[19]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[2]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[20]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[21]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[22]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[23]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[24]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[25]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[26]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b27  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [27]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[27]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b28  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [28]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[28]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b29  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [29]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[29]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[3]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b30  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [30]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[30]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b31  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [31]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[31]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b32  (
    .clk(clk100m),
    .d(1'b1),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[32]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[4]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[5]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[6]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[7]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[8]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[9]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg28_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[0]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[1]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[10]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[11]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[12]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[13]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[14]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[15]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[16]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[17]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[18]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[19]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[2]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[20]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[21]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[22]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[23]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[24]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[25]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[26]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b27  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [27]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[27]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b28  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [28]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[28]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b29  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [29]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[29]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[3]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b30  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [30]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[30]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b31  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [31]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[31]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b32  (
    .clk(clk100m),
    .d(1'b1),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[32]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[4]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[5]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[6]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[7]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[8]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[9]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg29_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[0]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[1]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[10]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[11]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[12]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[13]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[14]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[15]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[16]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[17]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[18]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[19]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[2]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[20]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[21]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[22]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[23]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[24]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[25]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[26]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b27  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [27]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[27]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b28  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [28]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[28]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b29  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [29]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[29]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[3]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b30  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [30]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[30]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b31  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [31]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[31]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b32  (
    .clk(clk100m),
    .d(1'b1),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[32]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[4]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[5]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[6]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[7]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[8]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[9]));  // src/AHB.v(78)
  reg_ar_as_w1 \U_AHB/reg2_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[0]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[1]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[10]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[11]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[12]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[13]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[14]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[15]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[16]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[17]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[18]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[19]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[2]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[20]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[21]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[22]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[23]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[24]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[25]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[26]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[3]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[4]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[5]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[6]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[7]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[8]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[9]));  // src/AHB.v(47)
  reg_sr_as_w1 \U_AHB/reg30_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[0]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[1]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[10]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[11]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[12]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[13]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[14]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[15]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[16]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[17]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[18]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[19]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[2]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[20]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[21]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[22]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[23]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[24]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[25]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[26]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b27  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [27]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[27]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b28  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [28]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[28]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b29  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [29]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[29]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[3]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b30  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [30]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[30]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b31  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [31]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[31]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b32  (
    .clk(clk100m),
    .d(1'b1),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[32]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[4]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[5]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[6]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[7]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[8]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[9]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg31_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[0]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[1]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[10]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[11]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[12]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[13]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[14]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[15]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[16]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[17]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[18]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[19]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[2]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[20]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[21]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[22]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[23]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[24]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[25]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[26]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b27  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [27]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[27]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b28  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [28]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[28]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b29  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [29]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[29]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[3]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b30  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [30]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[30]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b31  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [31]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[31]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b32  (
    .clk(clk100m),
    .d(1'b1),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[32]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[4]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[5]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[6]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[7]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[8]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[9]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg32_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[0]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[1]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[10]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[11]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[12]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[13]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[14]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[15]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[16]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[17]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[18]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[19]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[2]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[20]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[21]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[22]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[23]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[24]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[25]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[26]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b27  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [27]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[27]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b28  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [28]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[28]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b29  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [29]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[29]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[3]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b30  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [30]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[30]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b31  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [31]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[31]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b32  (
    .clk(clk100m),
    .d(1'b1),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[32]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[4]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[5]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[6]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[7]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[8]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[9]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg33_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[0]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[1]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[10]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[11]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[12]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[13]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[14]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[15]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[16]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[17]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[18]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[19]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[2]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[20]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[21]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[22]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[23]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[24]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[25]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[26]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b27  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [27]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[27]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b28  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [28]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[28]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b29  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [29]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[29]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[3]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b30  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [30]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[30]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b31  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [31]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[31]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b32  (
    .clk(clk100m),
    .d(1'b1),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[32]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[4]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[5]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[6]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[7]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[8]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[9]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg34_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[0]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[1]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[10]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[11]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[12]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[13]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[14]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[15]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[16]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[17]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[18]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[19]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[2]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[20]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[21]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[22]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[23]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[24]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[25]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[26]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b27  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [27]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[27]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b28  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [28]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[28]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b29  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [29]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[29]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[3]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b30  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [30]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[30]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b31  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [31]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[31]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[4]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[5]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[6]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[7]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[8]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[9]));  // src/AHB.v(84)
  reg_ar_as_w1 \U_AHB/reg35_b0  (
    .clk(clk100m),
    .d(\U_AHB/n118 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [0]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b1  (
    .clk(clk100m),
    .d(\U_AHB/n118 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [1]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b10  (
    .clk(clk100m),
    .d(\U_AHB/n118 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [10]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b11  (
    .clk(clk100m),
    .d(\U_AHB/n118 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [11]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b12  (
    .clk(clk100m),
    .d(\U_AHB/n118 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [12]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b13  (
    .clk(clk100m),
    .d(\U_AHB/n118 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [13]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b14  (
    .clk(clk100m),
    .d(\U_AHB/n118 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [14]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b15  (
    .clk(clk100m),
    .d(\U_AHB/n118 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [15]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b16  (
    .clk(clk100m),
    .d(\U_AHB/n118 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [16]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b17  (
    .clk(clk100m),
    .d(\U_AHB/n118 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [17]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b18  (
    .clk(clk100m),
    .d(\U_AHB/n118 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [18]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b19  (
    .clk(clk100m),
    .d(\U_AHB/n118 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [19]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b2  (
    .clk(clk100m),
    .d(\U_AHB/n118 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [2]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b20  (
    .clk(clk100m),
    .d(\U_AHB/n118 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [20]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b21  (
    .clk(clk100m),
    .d(\U_AHB/n118 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [21]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b22  (
    .clk(clk100m),
    .d(\U_AHB/n118 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [22]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b23  (
    .clk(clk100m),
    .d(\U_AHB/n118 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [23]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b24  (
    .clk(clk100m),
    .d(\U_AHB/n118 [24]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [24]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b25  (
    .clk(clk100m),
    .d(\U_AHB/n118 [25]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [25]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b26  (
    .clk(clk100m),
    .d(\U_AHB/n118 [26]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [26]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b27  (
    .clk(clk100m),
    .d(\U_AHB/n118 [27]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [27]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b28  (
    .clk(clk100m),
    .d(\U_AHB/n118 [28]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [28]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b29  (
    .clk(clk100m),
    .d(\U_AHB/n118 [29]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [29]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b3  (
    .clk(clk100m),
    .d(\U_AHB/n118 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [3]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b30  (
    .clk(clk100m),
    .d(\U_AHB/n118 [30]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [30]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b31  (
    .clk(clk100m),
    .d(\U_AHB/n118 [31]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [31]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b4  (
    .clk(clk100m),
    .d(\U_AHB/n118 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [4]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b5  (
    .clk(clk100m),
    .d(\U_AHB/n118 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [5]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b6  (
    .clk(clk100m),
    .d(\U_AHB/n118 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [6]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b7  (
    .clk(clk100m),
    .d(\U_AHB/n118 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [7]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b8  (
    .clk(clk100m),
    .d(\U_AHB/n118 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [8]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b9  (
    .clk(clk100m),
    .d(\U_AHB/n118 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [9]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg3_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[0]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[1]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[10]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[11]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[12]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[13]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[14]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[15]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[16]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[17]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[18]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[19]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[2]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[20]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[21]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[22]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[23]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[24]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[25]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[26]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[3]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[4]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[5]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[6]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[7]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[8]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[9]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg4_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[0]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[1]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[10]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[11]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[12]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[13]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[14]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[15]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[16]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[17]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[18]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[19]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[2]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[20]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[21]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[22]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[23]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[24]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[25]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[26]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[3]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[4]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[5]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[6]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[7]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[8]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[9]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg5_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[0]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[1]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[10]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[11]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[12]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[13]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[14]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[15]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[16]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[17]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[18]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[19]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[2]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[20]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[21]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[22]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[23]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[24]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[25]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[26]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[3]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[4]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[5]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[6]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[7]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[8]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[9]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg6_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[0]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[1]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[10]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[11]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[12]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[13]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[14]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[15]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[16]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[17]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[18]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[19]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[2]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[20]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[21]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[22]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[23]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[24]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[25]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[26]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[3]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[4]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[5]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[6]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[7]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[8]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[9]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg7_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[0]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[1]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[10]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[11]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[12]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[13]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[14]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[15]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[16]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[17]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[18]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[19]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[2]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[20]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[21]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[22]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[23]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[24]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[25]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[26]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[3]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[4]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[5]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[6]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[7]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[8]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[9]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg8_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[0]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[1]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[10]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[11]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[12]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[13]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[14]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[15]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[16]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[17]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[18]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[19]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[2]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[20]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[21]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[22]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[23]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[24]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[25]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[26]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[3]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[4]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[5]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[6]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[7]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[8]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[9]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg9_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[0]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[1]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[10]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[11]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[12]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[13]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[14]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[15]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[16]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[17]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[18]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[19]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[2]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[20]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[21]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[22]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[23]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[24]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[25]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[26]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[3]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[4]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[5]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[6]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[7]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[8]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[9]));  // src/AHB.v(54)
  EF2_PHY_PLL #(
    .CLKC0_CPHASE(4),
    .CLKC0_DIV(5),
    .CLKC0_DIV2_ENABLE("DISABLE"),
    .CLKC0_DUTY(0.500000),
    .CLKC0_DUTY50("ENABLE"),
    .CLKC0_DUTY_INT(3),
    .CLKC0_ENABLE("ENABLE"),
    .CLKC0_FPHASE(0),
    .CLKC1_CPHASE(9),
    .CLKC1_DIV(10),
    .CLKC1_DIV2_ENABLE("DISABLE"),
    .CLKC1_DUTY(0.500000),
    .CLKC1_DUTY50("ENABLE"),
    .CLKC1_DUTY_INT(5),
    .CLKC1_ENABLE("ENABLE"),
    .CLKC1_FPHASE(0),
    .CLKC2_CPHASE(39),
    .CLKC2_DIV(40),
    .CLKC2_DIV2_ENABLE("DISABLE"),
    .CLKC2_ENABLE("ENABLE"),
    .CLKC2_FPHASE(0),
    .CLKC3_CPHASE(124),
    .CLKC3_DIV(125),
    .CLKC3_DIV2_ENABLE("DISABLE"),
    .CLKC3_ENABLE("ENABLE"),
    .CLKC3_FPHASE(0),
    .CLKC4_CPHASE(1),
    .CLKC4_DIV(1),
    .CLKC4_DIV2_ENABLE("DISABLE"),
    .CLKC4_ENABLE("DISABLE"),
    .CLKC4_FPHASE(0),
    .CLKC5_CPHASE(1),
    .CLKC5_DIV(1),
    .CLKC5_DIV2_ENABLE("DISABLE"),
    .CLKC5_ENABLE("DISABLE"),
    .CLKC6_CPHASE(1),
    .CLKC6_DIV(1),
    .CLKC6_DIV2_ENABLE("DISABLE"),
    .CLKC6_ENABLE("DISABLE"),
    .DERIVE_PLL_CLOCKS("DISABLE"),
    .DPHASE_SOURCE("DISABLE"),
    .DYNCFG("DISABLE"),
    .FBCLK_DIV(40),
    .FEEDBK_MODE("NOCOMP"),
    .FEEDBK_PATH("VCO_PHASE_0"),
    .FIN("25.000"),
    .FREQ_LOCK_ACCURACY(2),
    .FREQ_OFFSET("0.000000"),
    .FREQ_OFFSET_INT("0"),
    .GEN_BASIC_CLOCK("DISABLE"),
    .GMC_GAIN(6),
    .GMC_TEST(14),
    .HIGH_SPEED_EN("ENABLE"),
    .ICP_CURRENT(3),
    .IF_ESCLKSTSW("DISABLE"),
    .INTFB_WAKE("DISABLE"),
    .INTPI(3),
    .KVCO(6),
    .LPF_CAPACITOR(3),
    .LPF_RESISTOR(2),
    .NORESET("DISABLE"),
    .ODIV_MUXC0("DIV"),
    .ODIV_MUXC1("DIV"),
    .ODIV_MUXC2("DIV"),
    .ODIV_MUXC3("DIV"),
    .ODIV_MUXC4("DIV"),
    .OFFSET_MODE("EXT"),
    .PLLC2RST_ENA("DISABLE"),
    .PLLC34RST_ENA("DISABLE"),
    .PLLMRST_ENA("DISABLE"),
    .PLLRST_ENA("ENABLE"),
    .PLL_LOCK_MODE(0),
    .PREDIV_MUXC0("VCO"),
    .PREDIV_MUXC1("VCO"),
    .PREDIV_MUXC2("VCO"),
    .PREDIV_MUXC3("VCO"),
    .PREDIV_MUXC4("VCO"),
    .PREDIV_MUXC5("VCO"),
    .PREDIV_MUXC6("VCO"),
    .PU_INTP("DISABLE"),
    .REFCLK_DIV(1),
    .REFCLK_SEL("INTERNAL"),
    .SSC_AMP("0.000000"),
    .SSC_ENABLE("DISABLE"),
    .SSC_FREQ_DIV(0),
    .SSC_MODE("Down"),
    .SSC_RNGE(0),
    .STDBY_ENABLE("DISABLE"),
    .STDBY_VCO_ENA("DISABLE"),
    .SYNC_ENABLE("DISABLE"),
    .VCO_NORESET("DISABLE"))
    \U_PLL/pll_inst  (
    .daddr(6'b000000),
    .dclk(1'b0),
    .dcs(1'b0),
    .di(8'b00000000),
    .dsm_refclk(1'b0),
    .dsm_rst(1'b0),
    .dwe(1'b0),
    .fbclk(1'b0),
    .frac_offset_valid(1'b0),
    .psclk(1'b0),
    .psclksel(3'b000),
    .psdown(1'b0),
    .psstep(1'b0),
    .refclk(clkin_pad),
    .reset(1'b0),
    .ssc_en(1'b0),
    .stdby(1'b0),
    .clkc({open_n229,open_n230,open_n231,open_n232,clk25m,clk100m_keep,open_n233}),
    .extlock(rstn));  // al_ip/PLL.v(92)
  EF2_PHY_PAD #(
    //.LOCATION("P70"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u100 (
    .ipad(limit_r[5]),
    .di(limit_r_pad[5]));  // CPLD_SOC_AHB_TOP.v(6)
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1000 (
    .a(_al_u995_o),
    .b(_al_u997_o),
    .c(_al_u999_o),
    .o(\PWM7/n0_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1001 (
    .a(\PWM7/n0_lutinv ),
    .b(\PWM7/stopreq ),
    .o(\PWM7/n1 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1002 (
    .a(\PWM7/n0_lutinv ),
    .b(\PWM7/n11 ),
    .o(\PWM7/mux3_b0_sel_is_3_o ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1003 (
    .a(\PWM7/n0_lutinv ),
    .b(\PWM7/n12 [9]),
    .c(freq7[9]),
    .o(\PWM7/n13 [9]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1004 (
    .a(\PWM7/n0_lutinv ),
    .b(\PWM7/n12 [8]),
    .c(freq7[8]),
    .o(\PWM7/n13 [8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1005 (
    .a(\PWM7/n0_lutinv ),
    .b(\PWM7/n12 [7]),
    .c(freq7[7]),
    .o(\PWM7/n13 [7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1006 (
    .a(\PWM7/n0_lutinv ),
    .b(\PWM7/n12 [6]),
    .c(freq7[6]),
    .o(\PWM7/n13 [6]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1007 (
    .a(\PWM7/n0_lutinv ),
    .b(\PWM7/n12 [5]),
    .c(freq7[5]),
    .o(\PWM7/n13 [5]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1008 (
    .a(\PWM7/n0_lutinv ),
    .b(\PWM7/n12 [4]),
    .c(freq7[4]),
    .o(\PWM7/n13 [4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1009 (
    .a(\PWM7/n0_lutinv ),
    .b(\PWM7/n12 [3]),
    .c(freq7[3]),
    .o(\PWM7/n13 [3]));
  EF2_PHY_PAD #(
    //.LOCATION("P59"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u101 (
    .ipad(limit_r[4]),
    .di(limit_r_pad[4]));  // CPLD_SOC_AHB_TOP.v(6)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1010 (
    .a(\PWM7/n0_lutinv ),
    .b(\PWM7/n12 [26]),
    .c(freq7[26]),
    .o(\PWM7/n13 [26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1011 (
    .a(\PWM7/n0_lutinv ),
    .b(\PWM7/n12 [25]),
    .c(freq7[25]),
    .o(\PWM7/n13 [25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1012 (
    .a(\PWM7/n0_lutinv ),
    .b(\PWM7/n12 [24]),
    .c(freq7[24]),
    .o(\PWM7/n13 [24]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1013 (
    .a(\PWM7/n0_lutinv ),
    .b(\PWM7/n12 [23]),
    .c(freq7[23]),
    .o(\PWM7/n13 [23]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1014 (
    .a(\PWM7/n0_lutinv ),
    .b(\PWM7/n12 [22]),
    .c(freq7[22]),
    .o(\PWM7/n13 [22]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1015 (
    .a(\PWM7/n0_lutinv ),
    .b(\PWM7/n12 [21]),
    .c(freq7[21]),
    .o(\PWM7/n13 [21]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1016 (
    .a(\PWM7/n0_lutinv ),
    .b(\PWM7/n12 [20]),
    .c(freq7[20]),
    .o(\PWM7/n13 [20]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1017 (
    .a(\PWM7/n0_lutinv ),
    .b(\PWM7/n12 [2]),
    .c(freq7[2]),
    .o(\PWM7/n13 [2]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1018 (
    .a(\PWM7/n0_lutinv ),
    .b(\PWM7/n12 [19]),
    .c(freq7[19]),
    .o(\PWM7/n13 [19]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1019 (
    .a(\PWM7/n0_lutinv ),
    .b(\PWM7/n12 [18]),
    .c(freq7[18]),
    .o(\PWM7/n13 [18]));
  EF2_PHY_PAD #(
    //.LOCATION("P57"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u102 (
    .ipad(limit_r[3]),
    .di(limit_r_pad[3]));  // CPLD_SOC_AHB_TOP.v(6)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1020 (
    .a(\PWM7/n0_lutinv ),
    .b(\PWM7/n12 [17]),
    .c(freq7[17]),
    .o(\PWM7/n13 [17]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1021 (
    .a(\PWM7/n0_lutinv ),
    .b(\PWM7/n12 [16]),
    .c(freq7[16]),
    .o(\PWM7/n13 [16]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1022 (
    .a(\PWM7/n0_lutinv ),
    .b(\PWM7/n12 [15]),
    .c(freq7[15]),
    .o(\PWM7/n13 [15]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1023 (
    .a(\PWM7/n0_lutinv ),
    .b(\PWM7/n12 [14]),
    .c(freq7[14]),
    .o(\PWM7/n13 [14]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1024 (
    .a(\PWM7/n0_lutinv ),
    .b(\PWM7/n12 [13]),
    .c(freq7[13]),
    .o(\PWM7/n13 [13]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1025 (
    .a(\PWM7/n0_lutinv ),
    .b(\PWM7/n12 [12]),
    .c(freq7[12]),
    .o(\PWM7/n13 [12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1026 (
    .a(\PWM7/n0_lutinv ),
    .b(\PWM7/n12 [11]),
    .c(freq7[11]),
    .o(\PWM7/n13 [11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1027 (
    .a(\PWM7/n0_lutinv ),
    .b(\PWM7/n12 [10]),
    .c(freq7[10]),
    .o(\PWM7/n13 [10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1028 (
    .a(\PWM7/n0_lutinv ),
    .b(\PWM7/n12 [1]),
    .c(freq7[1]),
    .o(\PWM7/n13 [1]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1029 (
    .a(\PWM7/n0_lutinv ),
    .b(\PWM7/n12 [0]),
    .c(freq7[0]),
    .o(\PWM7/n13 [0]));
  EF2_PHY_PAD #(
    //.LOCATION("P55"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u103 (
    .ipad(limit_r[2]),
    .di(limit_r_pad[2]));  // CPLD_SOC_AHB_TOP.v(6)
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1030 (
    .a(\PWM8/FreCnt [23]),
    .b(\PWM8/FreCnt [24]),
    .c(\PWM8/FreCnt [25]),
    .d(\PWM8/FreCnt [26]),
    .o(_al_u1030_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u1031 (
    .a(_al_u1030_o),
    .b(\PWM8/FreCnt [3]),
    .c(\PWM8/FreCnt [4]),
    .d(\PWM8/FreCnt [5]),
    .e(\PWM8/FreCnt [6]),
    .o(_al_u1031_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u1032 (
    .a(_al_u1031_o),
    .b(\PWM8/FreCnt [7]),
    .c(\PWM8/FreCnt [8]),
    .d(\PWM8/FreCnt [9]),
    .o(_al_u1032_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1033 (
    .a(\PWM8/FreCnt [0]),
    .b(\PWM8/FreCnt [1]),
    .c(\PWM8/FreCnt [10]),
    .d(\PWM8/FreCnt [11]),
    .o(_al_u1033_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u1034 (
    .a(_al_u1033_o),
    .b(\PWM8/FreCnt [12]),
    .c(\PWM8/FreCnt [13]),
    .d(\PWM8/FreCnt [14]),
    .e(\PWM8/FreCnt [15]),
    .o(_al_u1034_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1035 (
    .a(\PWM8/FreCnt [16]),
    .b(\PWM8/FreCnt [17]),
    .c(\PWM8/FreCnt [18]),
    .d(\PWM8/FreCnt [19]),
    .o(_al_u1035_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u1036 (
    .a(_al_u1035_o),
    .b(\PWM8/FreCnt [2]),
    .c(\PWM8/FreCnt [20]),
    .d(\PWM8/FreCnt [21]),
    .e(\PWM8/FreCnt [22]),
    .o(_al_u1036_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1037 (
    .a(_al_u1032_o),
    .b(_al_u1034_o),
    .c(_al_u1036_o),
    .o(\PWM8/n0_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1038 (
    .a(\PWM8/n0_lutinv ),
    .b(\PWM8/stopreq ),
    .o(\PWM8/n1 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1039 (
    .a(\PWM8/n0_lutinv ),
    .b(\PWM8/n11 ),
    .o(\PWM8/mux3_b0_sel_is_3_o ));
  EF2_PHY_PAD #(
    //.LOCATION("P49"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u104 (
    .ipad(limit_r[1]),
    .di(limit_r_pad[1]));  // CPLD_SOC_AHB_TOP.v(6)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1040 (
    .a(\PWM8/n0_lutinv ),
    .b(\PWM8/n12 [9]),
    .c(freq8[9]),
    .o(\PWM8/n13 [9]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1041 (
    .a(\PWM8/n0_lutinv ),
    .b(\PWM8/n12 [8]),
    .c(freq8[8]),
    .o(\PWM8/n13 [8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1042 (
    .a(\PWM8/n0_lutinv ),
    .b(\PWM8/n12 [7]),
    .c(freq8[7]),
    .o(\PWM8/n13 [7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1043 (
    .a(\PWM8/n0_lutinv ),
    .b(\PWM8/n12 [6]),
    .c(freq8[6]),
    .o(\PWM8/n13 [6]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1044 (
    .a(\PWM8/n0_lutinv ),
    .b(\PWM8/n12 [5]),
    .c(freq8[5]),
    .o(\PWM8/n13 [5]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1045 (
    .a(\PWM8/n0_lutinv ),
    .b(\PWM8/n12 [4]),
    .c(freq8[4]),
    .o(\PWM8/n13 [4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1046 (
    .a(\PWM8/n0_lutinv ),
    .b(\PWM8/n12 [3]),
    .c(freq8[3]),
    .o(\PWM8/n13 [3]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1047 (
    .a(\PWM8/n0_lutinv ),
    .b(\PWM8/n12 [26]),
    .c(freq8[26]),
    .o(\PWM8/n13 [26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1048 (
    .a(\PWM8/n0_lutinv ),
    .b(\PWM8/n12 [25]),
    .c(freq8[25]),
    .o(\PWM8/n13 [25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1049 (
    .a(\PWM8/n0_lutinv ),
    .b(\PWM8/n12 [24]),
    .c(freq8[24]),
    .o(\PWM8/n13 [24]));
  EF2_PHY_PAD #(
    //.LOCATION("P40"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u105 (
    .ipad(limit_r[0]),
    .di(limit_r_pad[0]));  // CPLD_SOC_AHB_TOP.v(6)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1050 (
    .a(\PWM8/n0_lutinv ),
    .b(\PWM8/n12 [23]),
    .c(freq8[23]),
    .o(\PWM8/n13 [23]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1051 (
    .a(\PWM8/n0_lutinv ),
    .b(\PWM8/n12 [22]),
    .c(freq8[22]),
    .o(\PWM8/n13 [22]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1052 (
    .a(\PWM8/n0_lutinv ),
    .b(\PWM8/n12 [21]),
    .c(freq8[21]),
    .o(\PWM8/n13 [21]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1053 (
    .a(\PWM8/n0_lutinv ),
    .b(\PWM8/n12 [20]),
    .c(freq8[20]),
    .o(\PWM8/n13 [20]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1054 (
    .a(\PWM8/n0_lutinv ),
    .b(\PWM8/n12 [2]),
    .c(freq8[2]),
    .o(\PWM8/n13 [2]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1055 (
    .a(\PWM8/n0_lutinv ),
    .b(\PWM8/n12 [19]),
    .c(freq8[19]),
    .o(\PWM8/n13 [19]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1056 (
    .a(\PWM8/n0_lutinv ),
    .b(\PWM8/n12 [18]),
    .c(freq8[18]),
    .o(\PWM8/n13 [18]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1057 (
    .a(\PWM8/n0_lutinv ),
    .b(\PWM8/n12 [17]),
    .c(freq8[17]),
    .o(\PWM8/n13 [17]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1058 (
    .a(\PWM8/n0_lutinv ),
    .b(\PWM8/n12 [16]),
    .c(freq8[16]),
    .o(\PWM8/n13 [16]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1059 (
    .a(\PWM8/n0_lutinv ),
    .b(\PWM8/n12 [15]),
    .c(freq8[15]),
    .o(\PWM8/n13 [15]));
  EF2_PHY_PAD #(
    //.LOCATION("P111"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u106 (
    .do({open_n382,open_n383,open_n384,pwm_pad[15]}),
    .opad(pwm[15]));  // CPLD_SOC_AHB_TOP.v(7)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1060 (
    .a(\PWM8/n0_lutinv ),
    .b(\PWM8/n12 [14]),
    .c(freq8[14]),
    .o(\PWM8/n13 [14]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1061 (
    .a(\PWM8/n0_lutinv ),
    .b(\PWM8/n12 [13]),
    .c(freq8[13]),
    .o(\PWM8/n13 [13]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1062 (
    .a(\PWM8/n0_lutinv ),
    .b(\PWM8/n12 [12]),
    .c(freq8[12]),
    .o(\PWM8/n13 [12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1063 (
    .a(\PWM8/n0_lutinv ),
    .b(\PWM8/n12 [11]),
    .c(freq8[11]),
    .o(\PWM8/n13 [11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1064 (
    .a(\PWM8/n0_lutinv ),
    .b(\PWM8/n12 [10]),
    .c(freq8[10]),
    .o(\PWM8/n13 [10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1065 (
    .a(\PWM8/n0_lutinv ),
    .b(\PWM8/n12 [1]),
    .c(freq8[1]),
    .o(\PWM8/n13 [1]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1066 (
    .a(\PWM8/n0_lutinv ),
    .b(\PWM8/n12 [0]),
    .c(freq8[0]),
    .o(\PWM8/n13 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1067 (
    .a(\PWM9/FreCnt [23]),
    .b(\PWM9/FreCnt [24]),
    .c(\PWM9/FreCnt [25]),
    .d(\PWM9/FreCnt [26]),
    .o(_al_u1067_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u1068 (
    .a(_al_u1067_o),
    .b(\PWM9/FreCnt [3]),
    .c(\PWM9/FreCnt [4]),
    .d(\PWM9/FreCnt [5]),
    .e(\PWM9/FreCnt [6]),
    .o(_al_u1068_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u1069 (
    .a(_al_u1068_o),
    .b(\PWM9/FreCnt [7]),
    .c(\PWM9/FreCnt [8]),
    .d(\PWM9/FreCnt [9]),
    .o(_al_u1069_o));
  EF2_PHY_PAD #(
    //.LOCATION("P112"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u107 (
    .do({open_n405,open_n406,open_n407,pwm_pad[14]}),
    .opad(pwm[14]));  // CPLD_SOC_AHB_TOP.v(7)
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1070 (
    .a(\PWM9/FreCnt [0]),
    .b(\PWM9/FreCnt [1]),
    .c(\PWM9/FreCnt [10]),
    .d(\PWM9/FreCnt [11]),
    .o(_al_u1070_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u1071 (
    .a(_al_u1070_o),
    .b(\PWM9/FreCnt [12]),
    .c(\PWM9/FreCnt [13]),
    .d(\PWM9/FreCnt [14]),
    .e(\PWM9/FreCnt [15]),
    .o(_al_u1071_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1072 (
    .a(\PWM9/FreCnt [16]),
    .b(\PWM9/FreCnt [17]),
    .c(\PWM9/FreCnt [18]),
    .d(\PWM9/FreCnt [19]),
    .o(_al_u1072_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u1073 (
    .a(_al_u1072_o),
    .b(\PWM9/FreCnt [2]),
    .c(\PWM9/FreCnt [20]),
    .d(\PWM9/FreCnt [21]),
    .e(\PWM9/FreCnt [22]),
    .o(_al_u1073_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1074 (
    .a(_al_u1069_o),
    .b(_al_u1071_o),
    .c(_al_u1073_o),
    .o(\PWM9/n0_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1075 (
    .a(\PWM9/n0_lutinv ),
    .b(\PWM9/stopreq ),
    .o(\PWM9/n1 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1076 (
    .a(\PWM9/n0_lutinv ),
    .b(\PWM9/n11 ),
    .o(\PWM9/mux3_b0_sel_is_3_o ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1077 (
    .a(\PWM9/n0_lutinv ),
    .b(\PWM9/n12 [9]),
    .c(freq9[9]),
    .o(\PWM9/n13 [9]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1078 (
    .a(\PWM9/n0_lutinv ),
    .b(\PWM9/n12 [8]),
    .c(freq9[8]),
    .o(\PWM9/n13 [8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1079 (
    .a(\PWM9/n0_lutinv ),
    .b(\PWM9/n12 [7]),
    .c(freq9[7]),
    .o(\PWM9/n13 [7]));
  EF2_PHY_PAD #(
    //.LOCATION("P115"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u108 (
    .do({open_n428,open_n429,open_n430,pwm_pad[13]}),
    .opad(pwm[13]));  // CPLD_SOC_AHB_TOP.v(7)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1080 (
    .a(\PWM9/n0_lutinv ),
    .b(\PWM9/n12 [6]),
    .c(freq9[6]),
    .o(\PWM9/n13 [6]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1081 (
    .a(\PWM9/n0_lutinv ),
    .b(\PWM9/n12 [5]),
    .c(freq9[5]),
    .o(\PWM9/n13 [5]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1082 (
    .a(\PWM9/n0_lutinv ),
    .b(\PWM9/n12 [4]),
    .c(freq9[4]),
    .o(\PWM9/n13 [4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1083 (
    .a(\PWM9/n0_lutinv ),
    .b(\PWM9/n12 [3]),
    .c(freq9[3]),
    .o(\PWM9/n13 [3]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1084 (
    .a(\PWM9/n0_lutinv ),
    .b(\PWM9/n12 [26]),
    .c(freq9[26]),
    .o(\PWM9/n13 [26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1085 (
    .a(\PWM9/n0_lutinv ),
    .b(\PWM9/n12 [25]),
    .c(freq9[25]),
    .o(\PWM9/n13 [25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1086 (
    .a(\PWM9/n0_lutinv ),
    .b(\PWM9/n12 [24]),
    .c(freq9[24]),
    .o(\PWM9/n13 [24]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1087 (
    .a(\PWM9/n0_lutinv ),
    .b(\PWM9/n12 [23]),
    .c(freq9[23]),
    .o(\PWM9/n13 [23]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1088 (
    .a(\PWM9/n0_lutinv ),
    .b(\PWM9/n12 [22]),
    .c(freq9[22]),
    .o(\PWM9/n13 [22]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1089 (
    .a(\PWM9/n0_lutinv ),
    .b(\PWM9/n12 [21]),
    .c(freq9[21]),
    .o(\PWM9/n13 [21]));
  EF2_PHY_PAD #(
    //.LOCATION("P117"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u109 (
    .do({open_n451,open_n452,open_n453,pwm_pad[12]}),
    .opad(pwm[12]));  // CPLD_SOC_AHB_TOP.v(7)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1090 (
    .a(\PWM9/n0_lutinv ),
    .b(\PWM9/n12 [20]),
    .c(freq9[20]),
    .o(\PWM9/n13 [20]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1091 (
    .a(\PWM9/n0_lutinv ),
    .b(\PWM9/n12 [2]),
    .c(freq9[2]),
    .o(\PWM9/n13 [2]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1092 (
    .a(\PWM9/n0_lutinv ),
    .b(\PWM9/n12 [19]),
    .c(freq9[19]),
    .o(\PWM9/n13 [19]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1093 (
    .a(\PWM9/n0_lutinv ),
    .b(\PWM9/n12 [18]),
    .c(freq9[18]),
    .o(\PWM9/n13 [18]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1094 (
    .a(\PWM9/n0_lutinv ),
    .b(\PWM9/n12 [17]),
    .c(freq9[17]),
    .o(\PWM9/n13 [17]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1095 (
    .a(\PWM9/n0_lutinv ),
    .b(\PWM9/n12 [16]),
    .c(freq9[16]),
    .o(\PWM9/n13 [16]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1096 (
    .a(\PWM9/n0_lutinv ),
    .b(\PWM9/n12 [15]),
    .c(freq9[15]),
    .o(\PWM9/n13 [15]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1097 (
    .a(\PWM9/n0_lutinv ),
    .b(\PWM9/n12 [14]),
    .c(freq9[14]),
    .o(\PWM9/n13 [14]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1098 (
    .a(\PWM9/n0_lutinv ),
    .b(\PWM9/n12 [13]),
    .c(freq9[13]),
    .o(\PWM9/n13 [13]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1099 (
    .a(\PWM9/n0_lutinv ),
    .b(\PWM9/n12 [12]),
    .c(freq9[12]),
    .o(\PWM9/n13 [12]));
  EF2_PHY_PAD #(
    //.LOCATION("P52"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u110 (
    .do({open_n474,open_n475,open_n476,pwm_pad[11]}),
    .opad(pwm[11]));  // CPLD_SOC_AHB_TOP.v(7)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1100 (
    .a(\PWM9/n0_lutinv ),
    .b(\PWM9/n12 [11]),
    .c(freq9[11]),
    .o(\PWM9/n13 [11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1101 (
    .a(\PWM9/n0_lutinv ),
    .b(\PWM9/n12 [10]),
    .c(freq9[10]),
    .o(\PWM9/n13 [10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1102 (
    .a(\PWM9/n0_lutinv ),
    .b(\PWM9/n12 [1]),
    .c(freq9[1]),
    .o(\PWM9/n13 [1]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1103 (
    .a(\PWM9/n0_lutinv ),
    .b(\PWM9/n12 [0]),
    .c(freq9[0]),
    .o(\PWM9/n13 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1104 (
    .a(\PWMA/FreCnt [23]),
    .b(\PWMA/FreCnt [24]),
    .c(\PWMA/FreCnt [25]),
    .d(\PWMA/FreCnt [26]),
    .o(_al_u1104_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u1105 (
    .a(_al_u1104_o),
    .b(\PWMA/FreCnt [3]),
    .c(\PWMA/FreCnt [4]),
    .d(\PWMA/FreCnt [5]),
    .e(\PWMA/FreCnt [6]),
    .o(_al_u1105_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u1106 (
    .a(_al_u1105_o),
    .b(\PWMA/FreCnt [7]),
    .c(\PWMA/FreCnt [8]),
    .d(\PWMA/FreCnt [9]),
    .o(_al_u1106_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1107 (
    .a(\PWMA/FreCnt [0]),
    .b(\PWMA/FreCnt [1]),
    .c(\PWMA/FreCnt [10]),
    .d(\PWMA/FreCnt [11]),
    .o(_al_u1107_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u1108 (
    .a(_al_u1107_o),
    .b(\PWMA/FreCnt [12]),
    .c(\PWMA/FreCnt [13]),
    .d(\PWMA/FreCnt [14]),
    .e(\PWMA/FreCnt [15]),
    .o(_al_u1108_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1109 (
    .a(\PWMA/FreCnt [16]),
    .b(\PWMA/FreCnt [17]),
    .c(\PWMA/FreCnt [18]),
    .d(\PWMA/FreCnt [19]),
    .o(_al_u1109_o));
  EF2_PHY_PAD #(
    //.LOCATION("P47"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u111 (
    .do({open_n497,open_n498,open_n499,pwm_pad[10]}),
    .opad(pwm[10]));  // CPLD_SOC_AHB_TOP.v(7)
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u1110 (
    .a(_al_u1109_o),
    .b(\PWMA/FreCnt [2]),
    .c(\PWMA/FreCnt [20]),
    .d(\PWMA/FreCnt [21]),
    .e(\PWMA/FreCnt [22]),
    .o(_al_u1110_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1111 (
    .a(_al_u1106_o),
    .b(_al_u1108_o),
    .c(_al_u1110_o),
    .o(\PWMA/n0_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1112 (
    .a(\PWMA/n0_lutinv ),
    .b(\PWMA/stopreq ),
    .o(\PWMA/n1 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1113 (
    .a(\PWMA/n0_lutinv ),
    .b(\PWMA/n11 ),
    .o(\PWMA/mux3_b0_sel_is_3_o ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1114 (
    .a(\PWMA/n0_lutinv ),
    .b(\PWMA/n12 [9]),
    .c(freqA[9]),
    .o(\PWMA/n13 [9]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1115 (
    .a(\PWMA/n0_lutinv ),
    .b(\PWMA/n12 [8]),
    .c(freqA[8]),
    .o(\PWMA/n13 [8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1116 (
    .a(\PWMA/n0_lutinv ),
    .b(\PWMA/n12 [7]),
    .c(freqA[7]),
    .o(\PWMA/n13 [7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1117 (
    .a(\PWMA/n0_lutinv ),
    .b(\PWMA/n12 [6]),
    .c(freqA[6]),
    .o(\PWMA/n13 [6]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1118 (
    .a(\PWMA/n0_lutinv ),
    .b(\PWMA/n12 [5]),
    .c(freqA[5]),
    .o(\PWMA/n13 [5]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1119 (
    .a(\PWMA/n0_lutinv ),
    .b(\PWMA/n12 [4]),
    .c(freqA[4]),
    .o(\PWMA/n13 [4]));
  EF2_PHY_PAD #(
    //.LOCATION("P44"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u112 (
    .do({open_n520,open_n521,open_n522,pwm_pad[9]}),
    .opad(pwm[9]));  // CPLD_SOC_AHB_TOP.v(7)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1120 (
    .a(\PWMA/n0_lutinv ),
    .b(\PWMA/n12 [3]),
    .c(freqA[3]),
    .o(\PWMA/n13 [3]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1121 (
    .a(\PWMA/n0_lutinv ),
    .b(\PWMA/n12 [26]),
    .c(freqA[26]),
    .o(\PWMA/n13 [26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1122 (
    .a(\PWMA/n0_lutinv ),
    .b(\PWMA/n12 [25]),
    .c(freqA[25]),
    .o(\PWMA/n13 [25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1123 (
    .a(\PWMA/n0_lutinv ),
    .b(\PWMA/n12 [24]),
    .c(freqA[24]),
    .o(\PWMA/n13 [24]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1124 (
    .a(\PWMA/n0_lutinv ),
    .b(\PWMA/n12 [23]),
    .c(freqA[23]),
    .o(\PWMA/n13 [23]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1125 (
    .a(\PWMA/n0_lutinv ),
    .b(\PWMA/n12 [22]),
    .c(freqA[22]),
    .o(\PWMA/n13 [22]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1126 (
    .a(\PWMA/n0_lutinv ),
    .b(\PWMA/n12 [21]),
    .c(freqA[21]),
    .o(\PWMA/n13 [21]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1127 (
    .a(\PWMA/n0_lutinv ),
    .b(\PWMA/n12 [20]),
    .c(freqA[20]),
    .o(\PWMA/n13 [20]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1128 (
    .a(\PWMA/n0_lutinv ),
    .b(\PWMA/n12 [2]),
    .c(freqA[2]),
    .o(\PWMA/n13 [2]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1129 (
    .a(\PWMA/n0_lutinv ),
    .b(\PWMA/n12 [19]),
    .c(freqA[19]),
    .o(\PWMA/n13 [19]));
  EF2_PHY_SPAD #(
    //.LOCATION("P107"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("16"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u113 (
    .do({open_n544,pwm_pad[8]}),
    .ts(1'b1),
    .opad(pwm[8]));  // CPLD_SOC_AHB_TOP.v(7)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1130 (
    .a(\PWMA/n0_lutinv ),
    .b(\PWMA/n12 [18]),
    .c(freqA[18]),
    .o(\PWMA/n13 [18]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1131 (
    .a(\PWMA/n0_lutinv ),
    .b(\PWMA/n12 [17]),
    .c(freqA[17]),
    .o(\PWMA/n13 [17]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1132 (
    .a(\PWMA/n0_lutinv ),
    .b(\PWMA/n12 [16]),
    .c(freqA[16]),
    .o(\PWMA/n13 [16]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1133 (
    .a(\PWMA/n0_lutinv ),
    .b(\PWMA/n12 [15]),
    .c(freqA[15]),
    .o(\PWMA/n13 [15]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1134 (
    .a(\PWMA/n0_lutinv ),
    .b(\PWMA/n12 [14]),
    .c(freqA[14]),
    .o(\PWMA/n13 [14]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1135 (
    .a(\PWMA/n0_lutinv ),
    .b(\PWMA/n12 [13]),
    .c(freqA[13]),
    .o(\PWMA/n13 [13]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1136 (
    .a(\PWMA/n0_lutinv ),
    .b(\PWMA/n12 [12]),
    .c(freqA[12]),
    .o(\PWMA/n13 [12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1137 (
    .a(\PWMA/n0_lutinv ),
    .b(\PWMA/n12 [11]),
    .c(freqA[11]),
    .o(\PWMA/n13 [11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1138 (
    .a(\PWMA/n0_lutinv ),
    .b(\PWMA/n12 [10]),
    .c(freqA[10]),
    .o(\PWMA/n13 [10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1139 (
    .a(\PWMA/n0_lutinv ),
    .b(\PWMA/n12 [1]),
    .c(freqA[1]),
    .o(\PWMA/n13 [1]));
  EF2_PHY_PAD #(
    //.LOCATION("P113"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u114 (
    .do({open_n552,open_n553,open_n554,pwm_pad[7]}),
    .opad(pwm[7]));  // CPLD_SOC_AHB_TOP.v(7)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1140 (
    .a(\PWMA/n0_lutinv ),
    .b(\PWMA/n12 [0]),
    .c(freqA[0]),
    .o(\PWMA/n13 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1141 (
    .a(\PWMB/FreCnt [23]),
    .b(\PWMB/FreCnt [24]),
    .c(\PWMB/FreCnt [25]),
    .d(\PWMB/FreCnt [26]),
    .o(_al_u1141_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u1142 (
    .a(_al_u1141_o),
    .b(\PWMB/FreCnt [3]),
    .c(\PWMB/FreCnt [4]),
    .d(\PWMB/FreCnt [5]),
    .e(\PWMB/FreCnt [6]),
    .o(_al_u1142_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u1143 (
    .a(_al_u1142_o),
    .b(\PWMB/FreCnt [7]),
    .c(\PWMB/FreCnt [8]),
    .d(\PWMB/FreCnt [9]),
    .o(_al_u1143_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1144 (
    .a(\PWMB/FreCnt [0]),
    .b(\PWMB/FreCnt [1]),
    .c(\PWMB/FreCnt [10]),
    .d(\PWMB/FreCnt [11]),
    .o(_al_u1144_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u1145 (
    .a(_al_u1144_o),
    .b(\PWMB/FreCnt [12]),
    .c(\PWMB/FreCnt [13]),
    .d(\PWMB/FreCnt [14]),
    .e(\PWMB/FreCnt [15]),
    .o(_al_u1145_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1146 (
    .a(\PWMB/FreCnt [16]),
    .b(\PWMB/FreCnt [17]),
    .c(\PWMB/FreCnt [18]),
    .d(\PWMB/FreCnt [19]),
    .o(_al_u1146_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u1147 (
    .a(_al_u1146_o),
    .b(\PWMB/FreCnt [2]),
    .c(\PWMB/FreCnt [20]),
    .d(\PWMB/FreCnt [21]),
    .e(\PWMB/FreCnt [22]),
    .o(_al_u1147_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1148 (
    .a(_al_u1143_o),
    .b(_al_u1145_o),
    .c(_al_u1147_o),
    .o(\PWMB/n0_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1149 (
    .a(\PWMB/n0_lutinv ),
    .b(\PWMB/stopreq ),
    .o(\PWMB/n1 ));
  EF2_PHY_PAD #(
    //.LOCATION("P121"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u115 (
    .do({open_n575,open_n576,open_n577,pwm_pad[6]}),
    .opad(pwm[6]));  // CPLD_SOC_AHB_TOP.v(7)
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1150 (
    .a(\PWMB/n0_lutinv ),
    .b(\PWMB/n11 ),
    .o(\PWMB/mux3_b0_sel_is_3_o ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1151 (
    .a(\PWMB/n0_lutinv ),
    .b(\PWMB/n12 [9]),
    .c(freqB[9]),
    .o(\PWMB/n13 [9]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1152 (
    .a(\PWMB/n0_lutinv ),
    .b(\PWMB/n12 [8]),
    .c(freqB[8]),
    .o(\PWMB/n13 [8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1153 (
    .a(\PWMB/n0_lutinv ),
    .b(\PWMB/n12 [7]),
    .c(freqB[7]),
    .o(\PWMB/n13 [7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1154 (
    .a(\PWMB/n0_lutinv ),
    .b(\PWMB/n12 [6]),
    .c(freqB[6]),
    .o(\PWMB/n13 [6]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1155 (
    .a(\PWMB/n0_lutinv ),
    .b(\PWMB/n12 [5]),
    .c(freqB[5]),
    .o(\PWMB/n13 [5]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1156 (
    .a(\PWMB/n0_lutinv ),
    .b(\PWMB/n12 [4]),
    .c(freqB[4]),
    .o(\PWMB/n13 [4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1157 (
    .a(\PWMB/n0_lutinv ),
    .b(\PWMB/n12 [3]),
    .c(freqB[3]),
    .o(\PWMB/n13 [3]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1158 (
    .a(\PWMB/n0_lutinv ),
    .b(\PWMB/n12 [26]),
    .c(freqB[26]),
    .o(\PWMB/n13 [26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1159 (
    .a(\PWMB/n0_lutinv ),
    .b(\PWMB/n12 [25]),
    .c(freqB[25]),
    .o(\PWMB/n13 [25]));
  EF2_PHY_SPAD #(
    //.LOCATION("P25"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("16"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u116 (
    .do({open_n599,pwm_pad[5]}),
    .ts(1'b1),
    .opad(pwm[5]));  // CPLD_SOC_AHB_TOP.v(7)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1160 (
    .a(\PWMB/n0_lutinv ),
    .b(\PWMB/n12 [24]),
    .c(freqB[24]),
    .o(\PWMB/n13 [24]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1161 (
    .a(\PWMB/n0_lutinv ),
    .b(\PWMB/n12 [23]),
    .c(freqB[23]),
    .o(\PWMB/n13 [23]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1162 (
    .a(\PWMB/n0_lutinv ),
    .b(\PWMB/n12 [22]),
    .c(freqB[22]),
    .o(\PWMB/n13 [22]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1163 (
    .a(\PWMB/n0_lutinv ),
    .b(\PWMB/n12 [21]),
    .c(freqB[21]),
    .o(\PWMB/n13 [21]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1164 (
    .a(\PWMB/n0_lutinv ),
    .b(\PWMB/n12 [20]),
    .c(freqB[20]),
    .o(\PWMB/n13 [20]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1165 (
    .a(\PWMB/n0_lutinv ),
    .b(\PWMB/n12 [2]),
    .c(freqB[2]),
    .o(\PWMB/n13 [2]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1166 (
    .a(\PWMB/n0_lutinv ),
    .b(\PWMB/n12 [19]),
    .c(freqB[19]),
    .o(\PWMB/n13 [19]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1167 (
    .a(\PWMB/n0_lutinv ),
    .b(\PWMB/n12 [18]),
    .c(freqB[18]),
    .o(\PWMB/n13 [18]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1168 (
    .a(\PWMB/n0_lutinv ),
    .b(\PWMB/n12 [17]),
    .c(freqB[17]),
    .o(\PWMB/n13 [17]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1169 (
    .a(\PWMB/n0_lutinv ),
    .b(\PWMB/n12 [16]),
    .c(freqB[16]),
    .o(\PWMB/n13 [16]));
  EF2_PHY_PAD #(
    //.LOCATION("P125"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u117 (
    .do({open_n607,open_n608,open_n609,pwm_pad[4]}),
    .opad(pwm[4]));  // CPLD_SOC_AHB_TOP.v(7)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1170 (
    .a(\PWMB/n0_lutinv ),
    .b(\PWMB/n12 [15]),
    .c(freqB[15]),
    .o(\PWMB/n13 [15]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1171 (
    .a(\PWMB/n0_lutinv ),
    .b(\PWMB/n12 [14]),
    .c(freqB[14]),
    .o(\PWMB/n13 [14]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1172 (
    .a(\PWMB/n0_lutinv ),
    .b(\PWMB/n12 [13]),
    .c(freqB[13]),
    .o(\PWMB/n13 [13]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1173 (
    .a(\PWMB/n0_lutinv ),
    .b(\PWMB/n12 [12]),
    .c(freqB[12]),
    .o(\PWMB/n13 [12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1174 (
    .a(\PWMB/n0_lutinv ),
    .b(\PWMB/n12 [11]),
    .c(freqB[11]),
    .o(\PWMB/n13 [11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1175 (
    .a(\PWMB/n0_lutinv ),
    .b(\PWMB/n12 [10]),
    .c(freqB[10]),
    .o(\PWMB/n13 [10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1176 (
    .a(\PWMB/n0_lutinv ),
    .b(\PWMB/n12 [1]),
    .c(freqB[1]),
    .o(\PWMB/n13 [1]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1177 (
    .a(\PWMB/n0_lutinv ),
    .b(\PWMB/n12 [0]),
    .c(freqB[0]),
    .o(\PWMB/n13 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1178 (
    .a(\PWMC/FreCnt [23]),
    .b(\PWMC/FreCnt [24]),
    .c(\PWMC/FreCnt [25]),
    .d(\PWMC/FreCnt [26]),
    .o(_al_u1178_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u1179 (
    .a(_al_u1178_o),
    .b(\PWMC/FreCnt [3]),
    .c(\PWMC/FreCnt [4]),
    .d(\PWMC/FreCnt [5]),
    .e(\PWMC/FreCnt [6]),
    .o(_al_u1179_o));
  EF2_PHY_PAD #(
    //.LOCATION("P126"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u118 (
    .do({open_n630,open_n631,open_n632,pwm_pad[3]}),
    .opad(pwm[3]));  // CPLD_SOC_AHB_TOP.v(7)
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u1180 (
    .a(_al_u1179_o),
    .b(\PWMC/FreCnt [7]),
    .c(\PWMC/FreCnt [8]),
    .d(\PWMC/FreCnt [9]),
    .o(_al_u1180_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1181 (
    .a(\PWMC/FreCnt [0]),
    .b(\PWMC/FreCnt [1]),
    .c(\PWMC/FreCnt [10]),
    .d(\PWMC/FreCnt [11]),
    .o(_al_u1181_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u1182 (
    .a(_al_u1181_o),
    .b(\PWMC/FreCnt [12]),
    .c(\PWMC/FreCnt [13]),
    .d(\PWMC/FreCnt [14]),
    .e(\PWMC/FreCnt [15]),
    .o(_al_u1182_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1183 (
    .a(\PWMC/FreCnt [16]),
    .b(\PWMC/FreCnt [17]),
    .c(\PWMC/FreCnt [18]),
    .d(\PWMC/FreCnt [19]),
    .o(_al_u1183_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u1184 (
    .a(_al_u1183_o),
    .b(\PWMC/FreCnt [2]),
    .c(\PWMC/FreCnt [20]),
    .d(\PWMC/FreCnt [21]),
    .e(\PWMC/FreCnt [22]),
    .o(_al_u1184_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1185 (
    .a(_al_u1180_o),
    .b(_al_u1182_o),
    .c(_al_u1184_o),
    .o(\PWMC/n0_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1186 (
    .a(\PWMC/n0_lutinv ),
    .b(\PWMC/stopreq ),
    .o(\PWMC/n1 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1187 (
    .a(\PWMC/n0_lutinv ),
    .b(\PWMC/n11 ),
    .o(\PWMC/mux3_b0_sel_is_3_o ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1188 (
    .a(\PWMC/n0_lutinv ),
    .b(\PWMC/n12 [9]),
    .c(freqC[9]),
    .o(\PWMC/n13 [9]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1189 (
    .a(\PWMC/n0_lutinv ),
    .b(\PWMC/n12 [8]),
    .c(freqC[8]),
    .o(\PWMC/n13 [8]));
  EF2_PHY_PAD #(
    //.LOCATION("P127"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u119 (
    .do({open_n653,open_n654,open_n655,pwm_pad[2]}),
    .opad(pwm[2]));  // CPLD_SOC_AHB_TOP.v(7)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1190 (
    .a(\PWMC/n0_lutinv ),
    .b(\PWMC/n12 [7]),
    .c(freqC[7]),
    .o(\PWMC/n13 [7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1191 (
    .a(\PWMC/n0_lutinv ),
    .b(\PWMC/n12 [6]),
    .c(freqC[6]),
    .o(\PWMC/n13 [6]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1192 (
    .a(\PWMC/n0_lutinv ),
    .b(\PWMC/n12 [5]),
    .c(freqC[5]),
    .o(\PWMC/n13 [5]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1193 (
    .a(\PWMC/n0_lutinv ),
    .b(\PWMC/n12 [4]),
    .c(freqC[4]),
    .o(\PWMC/n13 [4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1194 (
    .a(\PWMC/n0_lutinv ),
    .b(\PWMC/n12 [3]),
    .c(freqC[3]),
    .o(\PWMC/n13 [3]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1195 (
    .a(\PWMC/n0_lutinv ),
    .b(\PWMC/n12 [26]),
    .c(freqC[26]),
    .o(\PWMC/n13 [26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1196 (
    .a(\PWMC/n0_lutinv ),
    .b(\PWMC/n12 [25]),
    .c(freqC[25]),
    .o(\PWMC/n13 [25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1197 (
    .a(\PWMC/n0_lutinv ),
    .b(\PWMC/n12 [24]),
    .c(freqC[24]),
    .o(\PWMC/n13 [24]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1198 (
    .a(\PWMC/n0_lutinv ),
    .b(\PWMC/n12 [23]),
    .c(freqC[23]),
    .o(\PWMC/n13 [23]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1199 (
    .a(\PWMC/n0_lutinv ),
    .b(\PWMC/n12 [22]),
    .c(freqC[22]),
    .o(\PWMC/n13 [22]));
  EF2_PHY_PAD #(
    //.LOCATION("P128"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u120 (
    .do({open_n676,open_n677,open_n678,pwm_pad[1]}),
    .opad(pwm[1]));  // CPLD_SOC_AHB_TOP.v(7)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1200 (
    .a(\PWMC/n0_lutinv ),
    .b(\PWMC/n12 [21]),
    .c(freqC[21]),
    .o(\PWMC/n13 [21]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1201 (
    .a(\PWMC/n0_lutinv ),
    .b(\PWMC/n12 [20]),
    .c(freqC[20]),
    .o(\PWMC/n13 [20]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1202 (
    .a(\PWMC/n0_lutinv ),
    .b(\PWMC/n12 [2]),
    .c(freqC[2]),
    .o(\PWMC/n13 [2]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1203 (
    .a(\PWMC/n0_lutinv ),
    .b(\PWMC/n12 [19]),
    .c(freqC[19]),
    .o(\PWMC/n13 [19]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1204 (
    .a(\PWMC/n0_lutinv ),
    .b(\PWMC/n12 [18]),
    .c(freqC[18]),
    .o(\PWMC/n13 [18]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1205 (
    .a(\PWMC/n0_lutinv ),
    .b(\PWMC/n12 [17]),
    .c(freqC[17]),
    .o(\PWMC/n13 [17]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1206 (
    .a(\PWMC/n0_lutinv ),
    .b(\PWMC/n12 [16]),
    .c(freqC[16]),
    .o(\PWMC/n13 [16]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1207 (
    .a(\PWMC/n0_lutinv ),
    .b(\PWMC/n12 [15]),
    .c(freqC[15]),
    .o(\PWMC/n13 [15]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1208 (
    .a(\PWMC/n0_lutinv ),
    .b(\PWMC/n12 [14]),
    .c(freqC[14]),
    .o(\PWMC/n13 [14]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1209 (
    .a(\PWMC/n0_lutinv ),
    .b(\PWMC/n12 [13]),
    .c(freqC[13]),
    .o(\PWMC/n13 [13]));
  EF2_PHY_PAD #(
    //.LOCATION("P141"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u121 (
    .do({open_n699,open_n700,open_n701,pwm_pad[0]}),
    .opad(pwm[0]));  // CPLD_SOC_AHB_TOP.v(7)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1210 (
    .a(\PWMC/n0_lutinv ),
    .b(\PWMC/n12 [12]),
    .c(freqC[12]),
    .o(\PWMC/n13 [12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1211 (
    .a(\PWMC/n0_lutinv ),
    .b(\PWMC/n12 [11]),
    .c(freqC[11]),
    .o(\PWMC/n13 [11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1212 (
    .a(\PWMC/n0_lutinv ),
    .b(\PWMC/n12 [10]),
    .c(freqC[10]),
    .o(\PWMC/n13 [10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1213 (
    .a(\PWMC/n0_lutinv ),
    .b(\PWMC/n12 [1]),
    .c(freqC[1]),
    .o(\PWMC/n13 [1]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1214 (
    .a(\PWMC/n0_lutinv ),
    .b(\PWMC/n12 [0]),
    .c(freqC[0]),
    .o(\PWMC/n13 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1215 (
    .a(\PWMD/FreCnt [23]),
    .b(\PWMD/FreCnt [24]),
    .c(\PWMD/FreCnt [25]),
    .d(\PWMD/FreCnt [26]),
    .o(_al_u1215_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u1216 (
    .a(_al_u1215_o),
    .b(\PWMD/FreCnt [3]),
    .c(\PWMD/FreCnt [4]),
    .d(\PWMD/FreCnt [5]),
    .e(\PWMD/FreCnt [6]),
    .o(_al_u1216_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u1217 (
    .a(_al_u1216_o),
    .b(\PWMD/FreCnt [7]),
    .c(\PWMD/FreCnt [8]),
    .d(\PWMD/FreCnt [9]),
    .o(_al_u1217_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1218 (
    .a(\PWMD/FreCnt [0]),
    .b(\PWMD/FreCnt [1]),
    .c(\PWMD/FreCnt [10]),
    .d(\PWMD/FreCnt [11]),
    .o(_al_u1218_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u1219 (
    .a(_al_u1218_o),
    .b(\PWMD/FreCnt [12]),
    .c(\PWMD/FreCnt [13]),
    .d(\PWMD/FreCnt [14]),
    .e(\PWMD/FreCnt [15]),
    .o(_al_u1219_o));
  EF2_PHY_PAD #(
    //.LOCATION("P38"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u122 (
    .ipad(rst_n),
    .di(rst_n_pad));  // CPLD_SOC_AHB_TOP.v(4)
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1220 (
    .a(\PWMD/FreCnt [16]),
    .b(\PWMD/FreCnt [17]),
    .c(\PWMD/FreCnt [18]),
    .d(\PWMD/FreCnt [19]),
    .o(_al_u1220_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u1221 (
    .a(_al_u1220_o),
    .b(\PWMD/FreCnt [2]),
    .c(\PWMD/FreCnt [20]),
    .d(\PWMD/FreCnt [21]),
    .e(\PWMD/FreCnt [22]),
    .o(_al_u1221_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1222 (
    .a(_al_u1217_o),
    .b(_al_u1219_o),
    .c(_al_u1221_o),
    .o(\PWMD/n0_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1223 (
    .a(\PWMD/n0_lutinv ),
    .b(\PWMD/stopreq ),
    .o(\PWMD/n1 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1224 (
    .a(\PWMD/n0_lutinv ),
    .b(\PWMD/n11 ),
    .o(\PWMD/mux3_b0_sel_is_3_o ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1225 (
    .a(\PWMD/n0_lutinv ),
    .b(\PWMD/n12 [9]),
    .c(freqD[9]),
    .o(\PWMD/n13 [9]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1226 (
    .a(\PWMD/n0_lutinv ),
    .b(\PWMD/n12 [8]),
    .c(freqD[8]),
    .o(\PWMD/n13 [8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1227 (
    .a(\PWMD/n0_lutinv ),
    .b(\PWMD/n12 [7]),
    .c(freqD[7]),
    .o(\PWMD/n13 [7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1228 (
    .a(\PWMD/n0_lutinv ),
    .b(\PWMD/n12 [6]),
    .c(freqD[6]),
    .o(\PWMD/n13 [6]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1229 (
    .a(\PWMD/n0_lutinv ),
    .b(\PWMD/n12 [5]),
    .c(freqD[5]),
    .o(\PWMD/n13 [5]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1230 (
    .a(\PWMD/n0_lutinv ),
    .b(\PWMD/n12 [4]),
    .c(freqD[4]),
    .o(\PWMD/n13 [4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1231 (
    .a(\PWMD/n0_lutinv ),
    .b(\PWMD/n12 [3]),
    .c(freqD[3]),
    .o(\PWMD/n13 [3]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1232 (
    .a(\PWMD/n0_lutinv ),
    .b(\PWMD/n12 [26]),
    .c(freqD[26]),
    .o(\PWMD/n13 [26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1233 (
    .a(\PWMD/n0_lutinv ),
    .b(\PWMD/n12 [25]),
    .c(freqD[25]),
    .o(\PWMD/n13 [25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1234 (
    .a(\PWMD/n0_lutinv ),
    .b(\PWMD/n12 [24]),
    .c(freqD[24]),
    .o(\PWMD/n13 [24]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1235 (
    .a(\PWMD/n0_lutinv ),
    .b(\PWMD/n12 [23]),
    .c(freqD[23]),
    .o(\PWMD/n13 [23]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1236 (
    .a(\PWMD/n0_lutinv ),
    .b(\PWMD/n12 [22]),
    .c(freqD[22]),
    .o(\PWMD/n13 [22]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1237 (
    .a(\PWMD/n0_lutinv ),
    .b(\PWMD/n12 [21]),
    .c(freqD[21]),
    .o(\PWMD/n13 [21]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1238 (
    .a(\PWMD/n0_lutinv ),
    .b(\PWMD/n12 [20]),
    .c(freqD[20]),
    .o(\PWMD/n13 [20]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1239 (
    .a(\PWMD/n0_lutinv ),
    .b(\PWMD/n12 [2]),
    .c(freqD[2]),
    .o(\PWMD/n13 [2]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1240 (
    .a(\PWMD/n0_lutinv ),
    .b(\PWMD/n12 [19]),
    .c(freqD[19]),
    .o(\PWMD/n13 [19]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1241 (
    .a(\PWMD/n0_lutinv ),
    .b(\PWMD/n12 [18]),
    .c(freqD[18]),
    .o(\PWMD/n13 [18]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1242 (
    .a(\PWMD/n0_lutinv ),
    .b(\PWMD/n12 [17]),
    .c(freqD[17]),
    .o(\PWMD/n13 [17]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1243 (
    .a(\PWMD/n0_lutinv ),
    .b(\PWMD/n12 [16]),
    .c(freqD[16]),
    .o(\PWMD/n13 [16]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1244 (
    .a(\PWMD/n0_lutinv ),
    .b(\PWMD/n12 [15]),
    .c(freqD[15]),
    .o(\PWMD/n13 [15]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1245 (
    .a(\PWMD/n0_lutinv ),
    .b(\PWMD/n12 [14]),
    .c(freqD[14]),
    .o(\PWMD/n13 [14]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1246 (
    .a(\PWMD/n0_lutinv ),
    .b(\PWMD/n12 [13]),
    .c(freqD[13]),
    .o(\PWMD/n13 [13]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1247 (
    .a(\PWMD/n0_lutinv ),
    .b(\PWMD/n12 [12]),
    .c(freqD[12]),
    .o(\PWMD/n13 [12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1248 (
    .a(\PWMD/n0_lutinv ),
    .b(\PWMD/n12 [11]),
    .c(freqD[11]),
    .o(\PWMD/n13 [11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1249 (
    .a(\PWMD/n0_lutinv ),
    .b(\PWMD/n12 [10]),
    .c(freqD[10]),
    .o(\PWMD/n13 [10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1250 (
    .a(\PWMD/n0_lutinv ),
    .b(\PWMD/n12 [1]),
    .c(freqD[1]),
    .o(\PWMD/n13 [1]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1251 (
    .a(\PWMD/n0_lutinv ),
    .b(\PWMD/n12 [0]),
    .c(freqD[0]),
    .o(\PWMD/n13 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1252 (
    .a(\PWME/FreCnt [23]),
    .b(\PWME/FreCnt [24]),
    .c(\PWME/FreCnt [25]),
    .d(\PWME/FreCnt [26]),
    .o(_al_u1252_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u1253 (
    .a(_al_u1252_o),
    .b(\PWME/FreCnt [3]),
    .c(\PWME/FreCnt [4]),
    .d(\PWME/FreCnt [5]),
    .e(\PWME/FreCnt [6]),
    .o(_al_u1253_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u1254 (
    .a(_al_u1253_o),
    .b(\PWME/FreCnt [7]),
    .c(\PWME/FreCnt [8]),
    .d(\PWME/FreCnt [9]),
    .o(_al_u1254_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1255 (
    .a(\PWME/FreCnt [0]),
    .b(\PWME/FreCnt [1]),
    .c(\PWME/FreCnt [10]),
    .d(\PWME/FreCnt [11]),
    .o(_al_u1255_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u1256 (
    .a(_al_u1255_o),
    .b(\PWME/FreCnt [12]),
    .c(\PWME/FreCnt [13]),
    .d(\PWME/FreCnt [14]),
    .e(\PWME/FreCnt [15]),
    .o(_al_u1256_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1257 (
    .a(\PWME/FreCnt [16]),
    .b(\PWME/FreCnt [17]),
    .c(\PWME/FreCnt [18]),
    .d(\PWME/FreCnt [19]),
    .o(_al_u1257_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u1258 (
    .a(_al_u1257_o),
    .b(\PWME/FreCnt [2]),
    .c(\PWME/FreCnt [20]),
    .d(\PWME/FreCnt [21]),
    .e(\PWME/FreCnt [22]),
    .o(_al_u1258_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1259 (
    .a(_al_u1254_o),
    .b(_al_u1256_o),
    .c(_al_u1258_o),
    .o(\PWME/n0_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1260 (
    .a(\PWME/n0_lutinv ),
    .b(\PWME/stopreq ),
    .o(\PWME/n1 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1261 (
    .a(\PWME/n0_lutinv ),
    .b(\PWME/n11 ),
    .o(\PWME/mux3_b0_sel_is_3_o ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1262 (
    .a(\PWME/n0_lutinv ),
    .b(\PWME/n12 [9]),
    .c(freqE[9]),
    .o(\PWME/n13 [9]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1263 (
    .a(\PWME/n0_lutinv ),
    .b(\PWME/n12 [8]),
    .c(freqE[8]),
    .o(\PWME/n13 [8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1264 (
    .a(\PWME/n0_lutinv ),
    .b(\PWME/n12 [7]),
    .c(freqE[7]),
    .o(\PWME/n13 [7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1265 (
    .a(\PWME/n0_lutinv ),
    .b(\PWME/n12 [6]),
    .c(freqE[6]),
    .o(\PWME/n13 [6]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1266 (
    .a(\PWME/n0_lutinv ),
    .b(\PWME/n12 [5]),
    .c(freqE[5]),
    .o(\PWME/n13 [5]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1267 (
    .a(\PWME/n0_lutinv ),
    .b(\PWME/n12 [4]),
    .c(freqE[4]),
    .o(\PWME/n13 [4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1268 (
    .a(\PWME/n0_lutinv ),
    .b(\PWME/n12 [3]),
    .c(freqE[3]),
    .o(\PWME/n13 [3]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1269 (
    .a(\PWME/n0_lutinv ),
    .b(\PWME/n12 [26]),
    .c(freqE[26]),
    .o(\PWME/n13 [26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1270 (
    .a(\PWME/n0_lutinv ),
    .b(\PWME/n12 [25]),
    .c(freqE[25]),
    .o(\PWME/n13 [25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1271 (
    .a(\PWME/n0_lutinv ),
    .b(\PWME/n12 [24]),
    .c(freqE[24]),
    .o(\PWME/n13 [24]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1272 (
    .a(\PWME/n0_lutinv ),
    .b(\PWME/n12 [23]),
    .c(freqE[23]),
    .o(\PWME/n13 [23]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1273 (
    .a(\PWME/n0_lutinv ),
    .b(\PWME/n12 [22]),
    .c(freqE[22]),
    .o(\PWME/n13 [22]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1274 (
    .a(\PWME/n0_lutinv ),
    .b(\PWME/n12 [21]),
    .c(freqE[21]),
    .o(\PWME/n13 [21]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1275 (
    .a(\PWME/n0_lutinv ),
    .b(\PWME/n12 [20]),
    .c(freqE[20]),
    .o(\PWME/n13 [20]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1276 (
    .a(\PWME/n0_lutinv ),
    .b(\PWME/n12 [2]),
    .c(freqE[2]),
    .o(\PWME/n13 [2]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1277 (
    .a(\PWME/n0_lutinv ),
    .b(\PWME/n12 [19]),
    .c(freqE[19]),
    .o(\PWME/n13 [19]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1278 (
    .a(\PWME/n0_lutinv ),
    .b(\PWME/n12 [18]),
    .c(freqE[18]),
    .o(\PWME/n13 [18]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1279 (
    .a(\PWME/n0_lutinv ),
    .b(\PWME/n12 [17]),
    .c(freqE[17]),
    .o(\PWME/n13 [17]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1280 (
    .a(\PWME/n0_lutinv ),
    .b(\PWME/n12 [16]),
    .c(freqE[16]),
    .o(\PWME/n13 [16]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1281 (
    .a(\PWME/n0_lutinv ),
    .b(\PWME/n12 [15]),
    .c(freqE[15]),
    .o(\PWME/n13 [15]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1282 (
    .a(\PWME/n0_lutinv ),
    .b(\PWME/n12 [14]),
    .c(freqE[14]),
    .o(\PWME/n13 [14]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1283 (
    .a(\PWME/n0_lutinv ),
    .b(\PWME/n12 [13]),
    .c(freqE[13]),
    .o(\PWME/n13 [13]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1284 (
    .a(\PWME/n0_lutinv ),
    .b(\PWME/n12 [12]),
    .c(freqE[12]),
    .o(\PWME/n13 [12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1285 (
    .a(\PWME/n0_lutinv ),
    .b(\PWME/n12 [11]),
    .c(freqE[11]),
    .o(\PWME/n13 [11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1286 (
    .a(\PWME/n0_lutinv ),
    .b(\PWME/n12 [10]),
    .c(freqE[10]),
    .o(\PWME/n13 [10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1287 (
    .a(\PWME/n0_lutinv ),
    .b(\PWME/n12 [1]),
    .c(freqE[1]),
    .o(\PWME/n13 [1]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1288 (
    .a(\PWME/n0_lutinv ),
    .b(\PWME/n12 [0]),
    .c(freqE[0]),
    .o(\PWME/n13 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1289 (
    .a(\PWMF/FreCnt [23]),
    .b(\PWMF/FreCnt [24]),
    .c(\PWMF/FreCnt [25]),
    .d(\PWMF/FreCnt [26]),
    .o(_al_u1289_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u1290 (
    .a(_al_u1289_o),
    .b(\PWMF/FreCnt [3]),
    .c(\PWMF/FreCnt [4]),
    .d(\PWMF/FreCnt [5]),
    .e(\PWMF/FreCnt [6]),
    .o(_al_u1290_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u1291 (
    .a(_al_u1290_o),
    .b(\PWMF/FreCnt [7]),
    .c(\PWMF/FreCnt [8]),
    .d(\PWMF/FreCnt [9]),
    .o(_al_u1291_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1292 (
    .a(\PWMF/FreCnt [0]),
    .b(\PWMF/FreCnt [1]),
    .c(\PWMF/FreCnt [10]),
    .d(\PWMF/FreCnt [11]),
    .o(_al_u1292_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u1293 (
    .a(_al_u1292_o),
    .b(\PWMF/FreCnt [12]),
    .c(\PWMF/FreCnt [13]),
    .d(\PWMF/FreCnt [14]),
    .e(\PWMF/FreCnt [15]),
    .o(_al_u1293_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1294 (
    .a(\PWMF/FreCnt [16]),
    .b(\PWMF/FreCnt [17]),
    .c(\PWMF/FreCnt [18]),
    .d(\PWMF/FreCnt [19]),
    .o(_al_u1294_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u1295 (
    .a(_al_u1294_o),
    .b(\PWMF/FreCnt [2]),
    .c(\PWMF/FreCnt [20]),
    .d(\PWMF/FreCnt [21]),
    .e(\PWMF/FreCnt [22]),
    .o(_al_u1295_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1296 (
    .a(_al_u1291_o),
    .b(_al_u1293_o),
    .c(_al_u1295_o),
    .o(\PWMF/n0_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1297 (
    .a(\PWMF/n0_lutinv ),
    .b(\PWMF/stopreq ),
    .o(\PWMF/n1 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1298 (
    .a(\PWMF/n0_lutinv ),
    .b(\PWMF/n11 ),
    .o(\PWMF/mux3_b0_sel_is_3_o ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1299 (
    .a(\PWMF/n0_lutinv ),
    .b(\PWMF/n12 [9]),
    .c(freqF[9]),
    .o(\PWMF/n13 [9]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1300 (
    .a(\PWMF/n0_lutinv ),
    .b(\PWMF/n12 [8]),
    .c(freqF[8]),
    .o(\PWMF/n13 [8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1301 (
    .a(\PWMF/n0_lutinv ),
    .b(\PWMF/n12 [7]),
    .c(freqF[7]),
    .o(\PWMF/n13 [7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1302 (
    .a(\PWMF/n0_lutinv ),
    .b(\PWMF/n12 [6]),
    .c(freqF[6]),
    .o(\PWMF/n13 [6]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1303 (
    .a(\PWMF/n0_lutinv ),
    .b(\PWMF/n12 [5]),
    .c(freqF[5]),
    .o(\PWMF/n13 [5]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1304 (
    .a(\PWMF/n0_lutinv ),
    .b(\PWMF/n12 [4]),
    .c(freqF[4]),
    .o(\PWMF/n13 [4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1305 (
    .a(\PWMF/n0_lutinv ),
    .b(\PWMF/n12 [3]),
    .c(freqF[3]),
    .o(\PWMF/n13 [3]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1306 (
    .a(\PWMF/n0_lutinv ),
    .b(\PWMF/n12 [26]),
    .c(freqF[26]),
    .o(\PWMF/n13 [26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1307 (
    .a(\PWMF/n0_lutinv ),
    .b(\PWMF/n12 [25]),
    .c(freqF[25]),
    .o(\PWMF/n13 [25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1308 (
    .a(\PWMF/n0_lutinv ),
    .b(\PWMF/n12 [24]),
    .c(freqF[24]),
    .o(\PWMF/n13 [24]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1309 (
    .a(\PWMF/n0_lutinv ),
    .b(\PWMF/n12 [23]),
    .c(freqF[23]),
    .o(\PWMF/n13 [23]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1310 (
    .a(\PWMF/n0_lutinv ),
    .b(\PWMF/n12 [22]),
    .c(freqF[22]),
    .o(\PWMF/n13 [22]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1311 (
    .a(\PWMF/n0_lutinv ),
    .b(\PWMF/n12 [21]),
    .c(freqF[21]),
    .o(\PWMF/n13 [21]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1312 (
    .a(\PWMF/n0_lutinv ),
    .b(\PWMF/n12 [20]),
    .c(freqF[20]),
    .o(\PWMF/n13 [20]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1313 (
    .a(\PWMF/n0_lutinv ),
    .b(\PWMF/n12 [2]),
    .c(freqF[2]),
    .o(\PWMF/n13 [2]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1314 (
    .a(\PWMF/n0_lutinv ),
    .b(\PWMF/n12 [19]),
    .c(freqF[19]),
    .o(\PWMF/n13 [19]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1315 (
    .a(\PWMF/n0_lutinv ),
    .b(\PWMF/n12 [18]),
    .c(freqF[18]),
    .o(\PWMF/n13 [18]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1316 (
    .a(\PWMF/n0_lutinv ),
    .b(\PWMF/n12 [17]),
    .c(freqF[17]),
    .o(\PWMF/n13 [17]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1317 (
    .a(\PWMF/n0_lutinv ),
    .b(\PWMF/n12 [16]),
    .c(freqF[16]),
    .o(\PWMF/n13 [16]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1318 (
    .a(\PWMF/n0_lutinv ),
    .b(\PWMF/n12 [15]),
    .c(freqF[15]),
    .o(\PWMF/n13 [15]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1319 (
    .a(\PWMF/n0_lutinv ),
    .b(\PWMF/n12 [14]),
    .c(freqF[14]),
    .o(\PWMF/n13 [14]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1320 (
    .a(\PWMF/n0_lutinv ),
    .b(\PWMF/n12 [13]),
    .c(freqF[13]),
    .o(\PWMF/n13 [13]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1321 (
    .a(\PWMF/n0_lutinv ),
    .b(\PWMF/n12 [12]),
    .c(freqF[12]),
    .o(\PWMF/n13 [12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1322 (
    .a(\PWMF/n0_lutinv ),
    .b(\PWMF/n12 [11]),
    .c(freqF[11]),
    .o(\PWMF/n13 [11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1323 (
    .a(\PWMF/n0_lutinv ),
    .b(\PWMF/n12 [10]),
    .c(freqF[10]),
    .o(\PWMF/n13 [10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1324 (
    .a(\PWMF/n0_lutinv ),
    .b(\PWMF/n12 [1]),
    .c(freqF[1]),
    .o(\PWMF/n13 [1]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u1325 (
    .a(\PWMF/n0_lutinv ),
    .b(\PWMF/n12 [0]),
    .c(freqF[0]),
    .o(\PWMF/n13 [0]));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u1326 (
    .a(\U_AHB/h2h_hwrite ),
    .b(\U_AHB/h2h_haddr [13]),
    .c(\U_AHB/h2h_haddr [14]),
    .d(\U_AHB/h2h_haddr [8]),
    .o(\U_AHB/n38 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u1327 (
    .a(\U_AHB/h2h_hwrite ),
    .b(\U_AHB/h2h_haddr [13]),
    .c(\U_AHB/h2h_haddr [14]),
    .d(\U_AHB/h2h_haddr [7]),
    .o(\U_AHB/n36 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hdcf0))
    _al_u1328 (
    .a(\U_AHB/n38 ),
    .b(\U_AHB/n36 ),
    .c(gpio_out_pad[9]),
    .d(\U_AHB/h2h_hwdata [9]),
    .o(\U_AHB/n42 [9]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hdcf0))
    _al_u1329 (
    .a(\U_AHB/n38 ),
    .b(\U_AHB/n36 ),
    .c(gpio_out_pad[8]),
    .d(\U_AHB/h2h_hwdata [8]),
    .o(\U_AHB/n42 [8]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hdcf0))
    _al_u1330 (
    .a(\U_AHB/n38 ),
    .b(\U_AHB/n36 ),
    .c(gpio_out_pad[7]),
    .d(\U_AHB/h2h_hwdata [7]),
    .o(\U_AHB/n42 [7]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hdcf0))
    _al_u1331 (
    .a(\U_AHB/n38 ),
    .b(\U_AHB/n36 ),
    .c(gpio_out_pad[6]),
    .d(\U_AHB/h2h_hwdata [6]),
    .o(\U_AHB/n42 [6]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hdcf0))
    _al_u1332 (
    .a(\U_AHB/n38 ),
    .b(\U_AHB/n36 ),
    .c(gpio_out_pad[5]),
    .d(\U_AHB/h2h_hwdata [5]),
    .o(\U_AHB/n42 [5]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hdcf0))
    _al_u1333 (
    .a(\U_AHB/n38 ),
    .b(\U_AHB/n36 ),
    .c(gpio_out_pad[4]),
    .d(\U_AHB/h2h_hwdata [4]),
    .o(\U_AHB/n42 [4]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hdcf0))
    _al_u1334 (
    .a(\U_AHB/n38 ),
    .b(\U_AHB/n36 ),
    .c(gpio_out_pad[31]),
    .d(\U_AHB/h2h_hwdata [31]),
    .o(\U_AHB/n42 [31]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hdcf0))
    _al_u1335 (
    .a(\U_AHB/n38 ),
    .b(\U_AHB/n36 ),
    .c(gpio_out_pad[30]),
    .d(\U_AHB/h2h_hwdata [30]),
    .o(\U_AHB/n42 [30]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hdcf0))
    _al_u1336 (
    .a(\U_AHB/n38 ),
    .b(\U_AHB/n36 ),
    .c(gpio_out_pad[3]),
    .d(\U_AHB/h2h_hwdata [3]),
    .o(\U_AHB/n42 [3]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hdcf0))
    _al_u1337 (
    .a(\U_AHB/n38 ),
    .b(\U_AHB/n36 ),
    .c(gpio_out_pad[29]),
    .d(\U_AHB/h2h_hwdata [29]),
    .o(\U_AHB/n42 [29]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hdcf0))
    _al_u1338 (
    .a(\U_AHB/n38 ),
    .b(\U_AHB/n36 ),
    .c(gpio_out_pad[28]),
    .d(\U_AHB/h2h_hwdata [28]),
    .o(\U_AHB/n42 [28]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hdcf0))
    _al_u1339 (
    .a(\U_AHB/n38 ),
    .b(\U_AHB/n36 ),
    .c(gpio_out_pad[27]),
    .d(\U_AHB/h2h_hwdata [27]),
    .o(\U_AHB/n42 [27]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hdcf0))
    _al_u1340 (
    .a(\U_AHB/n38 ),
    .b(\U_AHB/n36 ),
    .c(gpio_out_pad[26]),
    .d(\U_AHB/h2h_hwdata [26]),
    .o(\U_AHB/n42 [26]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hdcf0))
    _al_u1341 (
    .a(\U_AHB/n38 ),
    .b(\U_AHB/n36 ),
    .c(gpio_out_pad[25]),
    .d(\U_AHB/h2h_hwdata [25]),
    .o(\U_AHB/n42 [25]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hdcf0))
    _al_u1342 (
    .a(\U_AHB/n38 ),
    .b(\U_AHB/n36 ),
    .c(gpio_out_pad[24]),
    .d(\U_AHB/h2h_hwdata [24]),
    .o(\U_AHB/n42 [24]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hdcf0))
    _al_u1343 (
    .a(\U_AHB/n38 ),
    .b(\U_AHB/n36 ),
    .c(gpio_out_pad[23]),
    .d(\U_AHB/h2h_hwdata [23]),
    .o(\U_AHB/n42 [23]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hdcf0))
    _al_u1344 (
    .a(\U_AHB/n38 ),
    .b(\U_AHB/n36 ),
    .c(gpio_out_pad[22]),
    .d(\U_AHB/h2h_hwdata [22]),
    .o(\U_AHB/n42 [22]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hdcf0))
    _al_u1345 (
    .a(\U_AHB/n38 ),
    .b(\U_AHB/n36 ),
    .c(gpio_out_pad[21]),
    .d(\U_AHB/h2h_hwdata [21]),
    .o(\U_AHB/n42 [21]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hdcf0))
    _al_u1346 (
    .a(\U_AHB/n38 ),
    .b(\U_AHB/n36 ),
    .c(gpio_out_pad[20]),
    .d(\U_AHB/h2h_hwdata [20]),
    .o(\U_AHB/n42 [20]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hdcf0))
    _al_u1347 (
    .a(\U_AHB/n38 ),
    .b(\U_AHB/n36 ),
    .c(gpio_out_pad[2]),
    .d(\U_AHB/h2h_hwdata [2]),
    .o(\U_AHB/n42 [2]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hdcf0))
    _al_u1348 (
    .a(\U_AHB/n38 ),
    .b(\U_AHB/n36 ),
    .c(gpio_out_pad[19]),
    .d(\U_AHB/h2h_hwdata [19]),
    .o(\U_AHB/n42 [19]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hdcf0))
    _al_u1349 (
    .a(\U_AHB/n38 ),
    .b(\U_AHB/n36 ),
    .c(gpio_out_pad[18]),
    .d(\U_AHB/h2h_hwdata [18]),
    .o(\U_AHB/n42 [18]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hdcf0))
    _al_u1350 (
    .a(\U_AHB/n38 ),
    .b(\U_AHB/n36 ),
    .c(gpio_out_pad[17]),
    .d(\U_AHB/h2h_hwdata [17]),
    .o(\U_AHB/n42 [17]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hdcf0))
    _al_u1351 (
    .a(\U_AHB/n38 ),
    .b(\U_AHB/n36 ),
    .c(gpio_out_pad[16]),
    .d(\U_AHB/h2h_hwdata [16]),
    .o(\U_AHB/n42 [16]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hdcf0))
    _al_u1352 (
    .a(\U_AHB/n38 ),
    .b(\U_AHB/n36 ),
    .c(gpio_out_pad[15]),
    .d(\U_AHB/h2h_hwdata [15]),
    .o(\U_AHB/n42 [15]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hdcf0))
    _al_u1353 (
    .a(\U_AHB/n38 ),
    .b(\U_AHB/n36 ),
    .c(gpio_out_pad[14]),
    .d(\U_AHB/h2h_hwdata [14]),
    .o(\U_AHB/n42 [14]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hdcf0))
    _al_u1354 (
    .a(\U_AHB/n38 ),
    .b(\U_AHB/n36 ),
    .c(gpio_out_pad[13]),
    .d(\U_AHB/h2h_hwdata [13]),
    .o(\U_AHB/n42 [13]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hdcf0))
    _al_u1355 (
    .a(\U_AHB/n38 ),
    .b(\U_AHB/n36 ),
    .c(gpio_out_pad[12]),
    .d(\U_AHB/h2h_hwdata [12]),
    .o(\U_AHB/n42 [12]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hdcf0))
    _al_u1356 (
    .a(\U_AHB/n38 ),
    .b(\U_AHB/n36 ),
    .c(gpio_out_pad[11]),
    .d(\U_AHB/h2h_hwdata [11]),
    .o(\U_AHB/n42 [11]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hdcf0))
    _al_u1357 (
    .a(\U_AHB/n38 ),
    .b(\U_AHB/n36 ),
    .c(gpio_out_pad[10]),
    .d(\U_AHB/h2h_hwdata [10]),
    .o(\U_AHB/n42 [10]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hdcf0))
    _al_u1358 (
    .a(\U_AHB/n38 ),
    .b(\U_AHB/n36 ),
    .c(gpio_out_pad[1]),
    .d(\U_AHB/h2h_hwdata [1]),
    .o(\U_AHB/n42 [1]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hdcf0))
    _al_u1359 (
    .a(\U_AHB/n38 ),
    .b(\U_AHB/n36 ),
    .c(gpio_out_pad[0]),
    .d(\U_AHB/h2h_hwdata [0]),
    .o(\U_AHB/n42 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1360 (
    .a(\PWM0/FreCnt [22]),
    .b(\PWM0/FreCnt [23]),
    .c(\PWM0/FreCntr [22]),
    .d(\PWM0/FreCntr [23]),
    .o(_al_u1360_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1361 (
    .a(_al_u1360_o),
    .b(\PWM0/FreCnt [17]),
    .c(\PWM0/FreCnt [8]),
    .d(\PWM0/FreCntr [17]),
    .e(\PWM0/FreCntr [8]),
    .o(_al_u1361_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1362 (
    .a(\PWM0/FreCnt [6]),
    .b(\PWM0/FreCnt [7]),
    .c(\PWM0/FreCntr [6]),
    .d(\PWM0/FreCntr [7]),
    .o(_al_u1362_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1363 (
    .a(_al_u1362_o),
    .b(\PWM0/FreCnt [4]),
    .c(\PWM0/FreCnt [9]),
    .d(\PWM0/FreCntr [4]),
    .e(\PWM0/FreCntr [9]),
    .o(_al_u1363_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1364 (
    .a(\PWM0/FreCnt [18]),
    .b(\PWM0/FreCnt [5]),
    .c(\PWM0/FreCntr [18]),
    .d(\PWM0/FreCntr [5]),
    .o(_al_u1364_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u1365 (
    .a(_al_u1361_o),
    .b(_al_u1363_o),
    .c(_al_u1364_o),
    .d(\PWM0/FreCnt [3]),
    .e(\PWM0/FreCntr [3]),
    .o(_al_u1365_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u1366 (
    .a(\PWM0/FreCnt [12]),
    .b(\PWM0/FreCnt [15]),
    .c(\PWM0/FreCntr [12]),
    .d(\PWM0/FreCntr [15]),
    .o(_al_u1366_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1367 (
    .a(\PWM0/FreCnt [10]),
    .b(\PWM0/FreCnt [2]),
    .c(\PWM0/FreCntr [10]),
    .d(\PWM0/FreCntr [2]),
    .o(_al_u1367_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D@C))"),
    .INIT(16'h8008))
    _al_u1368 (
    .a(_al_u1366_o),
    .b(_al_u1367_o),
    .c(\PWM0/FreCnt [21]),
    .d(\PWM0/FreCntr [21]),
    .o(_al_u1368_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1369 (
    .a(\PWM0/FreCnt [1]),
    .b(\PWM0/FreCntr [1]),
    .o(_al_u1369_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(E@C)*~(~D*B))"),
    .INIT(32'h50100501))
    _al_u1370 (
    .a(_al_u1369_o),
    .b(\PWM0/FreCnt [12]),
    .c(\PWM0/FreCnt [24]),
    .d(\PWM0/FreCntr [12]),
    .e(\PWM0/FreCntr [24]),
    .o(_al_u1370_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u1371 (
    .a(\PWM0/FreCnt [1]),
    .b(\PWM0/FreCnt [15]),
    .c(\PWM0/FreCntr [1]),
    .d(\PWM0/FreCntr [15]),
    .o(_al_u1371_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u1372 (
    .a(_al_u1368_o),
    .b(_al_u1370_o),
    .c(_al_u1371_o),
    .d(\PWM0/FreCnt [0]),
    .e(\PWM0/FreCntr [0]),
    .o(_al_u1372_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1373 (
    .a(\PWM0/FreCnt [11]),
    .b(\PWM0/FreCnt [25]),
    .c(\PWM0/FreCntr [11]),
    .d(\PWM0/FreCntr [25]),
    .o(_al_u1373_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1374 (
    .a(_al_u1373_o),
    .b(\PWM0/FreCnt [14]),
    .c(\PWM0/FreCnt [20]),
    .d(\PWM0/FreCntr [14]),
    .e(\PWM0/FreCntr [20]),
    .o(_al_u1374_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1375 (
    .a(\PWM0/FreCnt [16]),
    .b(\PWM0/FreCnt [26]),
    .c(\PWM0/FreCntr [16]),
    .d(\PWM0/FreCntr [26]),
    .o(_al_u1375_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1376 (
    .a(_al_u1375_o),
    .b(\PWM0/FreCnt [13]),
    .c(\PWM0/FreCnt [19]),
    .d(\PWM0/FreCntr [13]),
    .e(\PWM0/FreCntr [19]),
    .o(_al_u1376_o));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~(D*C*B*A))"),
    .INIT(32'hffff8000))
    _al_u1377 (
    .a(_al_u1365_o),
    .b(_al_u1372_o),
    .c(_al_u1374_o),
    .d(_al_u1376_o),
    .e(pwm_pad[0]),
    .o(\pwm[0]_d ));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1378 (
    .a(\PWM1/FreCnt [22]),
    .b(\PWM1/FreCnt [23]),
    .c(\PWM1/FreCntr [22]),
    .d(\PWM1/FreCntr [23]),
    .o(_al_u1378_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1379 (
    .a(_al_u1378_o),
    .b(\PWM1/FreCnt [7]),
    .c(\PWM1/FreCnt [9]),
    .d(\PWM1/FreCntr [7]),
    .e(\PWM1/FreCntr [9]),
    .o(_al_u1379_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1380 (
    .a(\PWM1/FreCnt [17]),
    .b(\PWM1/FreCnt [8]),
    .c(\PWM1/FreCntr [17]),
    .d(\PWM1/FreCntr [8]),
    .o(_al_u1380_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1381 (
    .a(_al_u1380_o),
    .b(\PWM1/FreCnt [11]),
    .c(\PWM1/FreCnt [24]),
    .d(\PWM1/FreCntr [11]),
    .e(\PWM1/FreCntr [24]),
    .o(_al_u1381_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1382 (
    .a(\PWM1/FreCnt [18]),
    .b(\PWM1/FreCnt [5]),
    .c(\PWM1/FreCntr [18]),
    .d(\PWM1/FreCntr [5]),
    .o(_al_u1382_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u1383 (
    .a(_al_u1379_o),
    .b(_al_u1381_o),
    .c(_al_u1382_o),
    .d(\PWM1/FreCnt [4]),
    .e(\PWM1/FreCntr [4]),
    .o(_al_u1383_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1384 (
    .a(\PWM1/FreCnt [0]),
    .b(\PWM1/FreCnt [10]),
    .c(\PWM1/FreCntr [0]),
    .d(\PWM1/FreCntr [10]),
    .o(_al_u1384_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u1385 (
    .a(\PWM1/FreCnt [12]),
    .b(\PWM1/FreCnt [15]),
    .c(\PWM1/FreCntr [12]),
    .d(\PWM1/FreCntr [15]),
    .o(_al_u1385_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D@C))"),
    .INIT(16'h8008))
    _al_u1386 (
    .a(_al_u1384_o),
    .b(_al_u1385_o),
    .c(\PWM1/FreCnt [21]),
    .d(\PWM1/FreCntr [21]),
    .o(_al_u1386_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u1387 (
    .a(\PWM1/FreCnt [12]),
    .b(\PWM1/FreCnt [15]),
    .c(\PWM1/FreCntr [12]),
    .d(\PWM1/FreCntr [15]),
    .o(_al_u1387_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1388 (
    .a(\PWM1/FreCnt [1]),
    .b(\PWM1/FreCnt [3]),
    .c(\PWM1/FreCntr [1]),
    .d(\PWM1/FreCntr [3]),
    .o(_al_u1388_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u1389 (
    .a(_al_u1386_o),
    .b(_al_u1387_o),
    .c(_al_u1388_o),
    .d(\PWM1/FreCnt [6]),
    .e(\PWM1/FreCntr [6]),
    .o(_al_u1389_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1390 (
    .a(\PWM1/FreCnt [14]),
    .b(\PWM1/FreCnt [25]),
    .c(\PWM1/FreCntr [14]),
    .d(\PWM1/FreCntr [25]),
    .o(_al_u1390_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1391 (
    .a(_al_u1390_o),
    .b(\PWM1/FreCnt [20]),
    .c(\PWM1/FreCnt [26]),
    .d(\PWM1/FreCntr [20]),
    .e(\PWM1/FreCntr [26]),
    .o(_al_u1391_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1392 (
    .a(\PWM1/FreCnt [13]),
    .b(\PWM1/FreCnt [16]),
    .c(\PWM1/FreCntr [13]),
    .d(\PWM1/FreCntr [16]),
    .o(_al_u1392_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1393 (
    .a(_al_u1392_o),
    .b(\PWM1/FreCnt [19]),
    .c(\PWM1/FreCnt [2]),
    .d(\PWM1/FreCntr [19]),
    .e(\PWM1/FreCntr [2]),
    .o(_al_u1393_o));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~(D*C*B*A))"),
    .INIT(32'hffff8000))
    _al_u1394 (
    .a(_al_u1383_o),
    .b(_al_u1389_o),
    .c(_al_u1391_o),
    .d(_al_u1393_o),
    .e(pwm_pad[1]),
    .o(\pwm[1]_d ));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1395 (
    .a(\PWM2/FreCnt [22]),
    .b(\PWM2/FreCnt [23]),
    .c(\PWM2/FreCntr [22]),
    .d(\PWM2/FreCntr [23]),
    .o(_al_u1395_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1396 (
    .a(_al_u1395_o),
    .b(\PWM2/FreCnt [17]),
    .c(\PWM2/FreCnt [8]),
    .d(\PWM2/FreCntr [17]),
    .e(\PWM2/FreCntr [8]),
    .o(_al_u1396_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1397 (
    .a(\PWM2/FreCnt [6]),
    .b(\PWM2/FreCnt [7]),
    .c(\PWM2/FreCntr [6]),
    .d(\PWM2/FreCntr [7]),
    .o(_al_u1397_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1398 (
    .a(_al_u1397_o),
    .b(\PWM2/FreCnt [11]),
    .c(\PWM2/FreCnt [9]),
    .d(\PWM2/FreCntr [11]),
    .e(\PWM2/FreCntr [9]),
    .o(_al_u1398_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1399 (
    .a(\PWM2/FreCnt [18]),
    .b(\PWM2/FreCnt [5]),
    .c(\PWM2/FreCntr [18]),
    .d(\PWM2/FreCntr [5]),
    .o(_al_u1399_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u1400 (
    .a(_al_u1396_o),
    .b(_al_u1398_o),
    .c(_al_u1399_o),
    .d(\PWM2/FreCnt [4]),
    .e(\PWM2/FreCntr [4]),
    .o(_al_u1400_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u1401 (
    .a(\PWM2/FreCnt [12]),
    .b(\PWM2/FreCnt [15]),
    .c(\PWM2/FreCntr [12]),
    .d(\PWM2/FreCntr [15]),
    .o(_al_u1401_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1402 (
    .a(\PWM2/FreCnt [10]),
    .b(\PWM2/FreCnt [3]),
    .c(\PWM2/FreCntr [10]),
    .d(\PWM2/FreCntr [3]),
    .o(_al_u1402_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D@C))"),
    .INIT(16'h8008))
    _al_u1403 (
    .a(_al_u1401_o),
    .b(_al_u1402_o),
    .c(\PWM2/FreCnt [21]),
    .d(\PWM2/FreCntr [21]),
    .o(_al_u1403_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1404 (
    .a(\PWM2/FreCnt [1]),
    .b(\PWM2/FreCntr [1]),
    .o(_al_u1404_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(E@C)*~(~D*B))"),
    .INIT(32'h50100501))
    _al_u1405 (
    .a(_al_u1404_o),
    .b(\PWM2/FreCnt [12]),
    .c(\PWM2/FreCnt [24]),
    .d(\PWM2/FreCntr [12]),
    .e(\PWM2/FreCntr [24]),
    .o(_al_u1405_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u1406 (
    .a(\PWM2/FreCnt [1]),
    .b(\PWM2/FreCnt [15]),
    .c(\PWM2/FreCntr [1]),
    .d(\PWM2/FreCntr [15]),
    .o(_al_u1406_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u1407 (
    .a(_al_u1403_o),
    .b(_al_u1405_o),
    .c(_al_u1406_o),
    .d(\PWM2/FreCnt [0]),
    .e(\PWM2/FreCntr [0]),
    .o(_al_u1407_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1408 (
    .a(\PWM2/FreCnt [14]),
    .b(\PWM2/FreCnt [25]),
    .c(\PWM2/FreCntr [14]),
    .d(\PWM2/FreCntr [25]),
    .o(_al_u1408_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1409 (
    .a(_al_u1408_o),
    .b(\PWM2/FreCnt [20]),
    .c(\PWM2/FreCnt [26]),
    .d(\PWM2/FreCntr [20]),
    .e(\PWM2/FreCntr [26]),
    .o(_al_u1409_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1410 (
    .a(\PWM2/FreCnt [13]),
    .b(\PWM2/FreCnt [16]),
    .c(\PWM2/FreCntr [13]),
    .d(\PWM2/FreCntr [16]),
    .o(_al_u1410_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1411 (
    .a(_al_u1410_o),
    .b(\PWM2/FreCnt [19]),
    .c(\PWM2/FreCnt [2]),
    .d(\PWM2/FreCntr [19]),
    .e(\PWM2/FreCntr [2]),
    .o(_al_u1411_o));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~(D*C*B*A))"),
    .INIT(32'hffff8000))
    _al_u1412 (
    .a(_al_u1400_o),
    .b(_al_u1407_o),
    .c(_al_u1409_o),
    .d(_al_u1411_o),
    .e(pwm_pad[2]),
    .o(\pwm[2]_d ));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1413 (
    .a(\PWM3/FreCnt [16]),
    .b(\PWM3/FreCnt [3]),
    .c(\PWM3/FreCntr [16]),
    .d(\PWM3/FreCntr [3]),
    .o(_al_u1413_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1414 (
    .a(_al_u1413_o),
    .b(\PWM3/FreCnt [18]),
    .c(\PWM3/FreCnt [5]),
    .d(\PWM3/FreCntr [18]),
    .e(\PWM3/FreCntr [5]),
    .o(_al_u1414_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1415 (
    .a(\PWM3/FreCnt [22]),
    .b(\PWM3/FreCnt [23]),
    .c(\PWM3/FreCntr [22]),
    .d(\PWM3/FreCntr [23]),
    .o(_al_u1415_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1416 (
    .a(_al_u1415_o),
    .b(\PWM3/FreCnt [17]),
    .c(\PWM3/FreCnt [8]),
    .d(\PWM3/FreCntr [17]),
    .e(\PWM3/FreCntr [8]),
    .o(_al_u1416_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1417 (
    .a(\PWM3/FreCnt [20]),
    .b(\PWM3/FreCnt [26]),
    .c(\PWM3/FreCntr [20]),
    .d(\PWM3/FreCntr [26]),
    .o(_al_u1417_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u1418 (
    .a(_al_u1414_o),
    .b(_al_u1416_o),
    .c(_al_u1417_o),
    .d(\PWM3/FreCnt [14]),
    .e(\PWM3/FreCntr [14]),
    .o(_al_u1418_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u1419 (
    .a(\PWM3/FreCnt [12]),
    .b(\PWM3/FreCnt [15]),
    .c(\PWM3/FreCntr [12]),
    .d(\PWM3/FreCntr [15]),
    .o(_al_u1419_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u1420 (
    .a(_al_u1419_o),
    .b(\PWM3/FreCnt [6]),
    .c(\PWM3/FreCntr [6]),
    .o(_al_u1420_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1421 (
    .a(\PWM3/FreCnt [0]),
    .b(\PWM3/FreCnt [24]),
    .c(\PWM3/FreCntr [0]),
    .d(\PWM3/FreCntr [24]),
    .o(_al_u1421_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1422 (
    .a(_al_u1421_o),
    .b(\PWM3/FreCnt [13]),
    .c(\PWM3/FreCnt [19]),
    .d(\PWM3/FreCntr [13]),
    .e(\PWM3/FreCntr [19]),
    .o(_al_u1422_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u1423 (
    .a(\PWM3/FreCnt [12]),
    .b(\PWM3/FreCnt [15]),
    .c(\PWM3/FreCntr [12]),
    .d(\PWM3/FreCntr [15]),
    .o(_al_u1423_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u1424 (
    .a(_al_u1420_o),
    .b(_al_u1422_o),
    .c(_al_u1423_o),
    .d(\PWM3/FreCnt [21]),
    .e(\PWM3/FreCntr [21]),
    .o(_al_u1424_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1425 (
    .a(\PWM3/FreCnt [7]),
    .b(\PWM3/FreCnt [9]),
    .c(\PWM3/FreCntr [7]),
    .d(\PWM3/FreCntr [9]),
    .o(_al_u1425_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1426 (
    .a(_al_u1425_o),
    .b(\PWM3/FreCnt [11]),
    .c(\PWM3/FreCnt [4]),
    .d(\PWM3/FreCntr [11]),
    .e(\PWM3/FreCntr [4]),
    .o(_al_u1426_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1427 (
    .a(\PWM3/FreCnt [2]),
    .b(\PWM3/FreCnt [25]),
    .c(\PWM3/FreCntr [2]),
    .d(\PWM3/FreCntr [25]),
    .o(_al_u1427_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1428 (
    .a(_al_u1427_o),
    .b(\PWM3/FreCnt [1]),
    .c(\PWM3/FreCnt [10]),
    .d(\PWM3/FreCntr [1]),
    .e(\PWM3/FreCntr [10]),
    .o(_al_u1428_o));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~(D*C*B*A))"),
    .INIT(32'hffff8000))
    _al_u1429 (
    .a(_al_u1418_o),
    .b(_al_u1424_o),
    .c(_al_u1426_o),
    .d(_al_u1428_o),
    .e(pwm_pad[3]),
    .o(\pwm[3]_d ));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1430 (
    .a(\PWM4/FreCnt [16]),
    .b(\PWM4/FreCnt [4]),
    .c(\PWM4/FreCntr [16]),
    .d(\PWM4/FreCntr [4]),
    .o(_al_u1430_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1431 (
    .a(_al_u1430_o),
    .b(\PWM4/FreCnt [18]),
    .c(\PWM4/FreCnt [5]),
    .d(\PWM4/FreCntr [18]),
    .e(\PWM4/FreCntr [5]),
    .o(_al_u1431_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1432 (
    .a(\PWM4/FreCnt [22]),
    .b(\PWM4/FreCnt [23]),
    .c(\PWM4/FreCntr [22]),
    .d(\PWM4/FreCntr [23]),
    .o(_al_u1432_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1433 (
    .a(_al_u1432_o),
    .b(\PWM4/FreCnt [17]),
    .c(\PWM4/FreCnt [8]),
    .d(\PWM4/FreCntr [17]),
    .e(\PWM4/FreCntr [8]),
    .o(_al_u1433_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1434 (
    .a(\PWM4/FreCnt [20]),
    .b(\PWM4/FreCnt [26]),
    .c(\PWM4/FreCntr [20]),
    .d(\PWM4/FreCntr [26]),
    .o(_al_u1434_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u1435 (
    .a(_al_u1431_o),
    .b(_al_u1433_o),
    .c(_al_u1434_o),
    .d(\PWM4/FreCnt [14]),
    .e(\PWM4/FreCntr [14]),
    .o(_al_u1435_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u1436 (
    .a(\PWM4/FreCnt [12]),
    .b(\PWM4/FreCnt [15]),
    .c(\PWM4/FreCntr [12]),
    .d(\PWM4/FreCntr [15]),
    .o(_al_u1436_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u1437 (
    .a(_al_u1436_o),
    .b(\PWM4/FreCnt [6]),
    .c(\PWM4/FreCntr [6]),
    .o(_al_u1437_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1438 (
    .a(\PWM4/FreCnt [0]),
    .b(\PWM4/FreCnt [24]),
    .c(\PWM4/FreCntr [0]),
    .d(\PWM4/FreCntr [24]),
    .o(_al_u1438_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1439 (
    .a(_al_u1438_o),
    .b(\PWM4/FreCnt [13]),
    .c(\PWM4/FreCnt [19]),
    .d(\PWM4/FreCntr [13]),
    .e(\PWM4/FreCntr [19]),
    .o(_al_u1439_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u1440 (
    .a(\PWM4/FreCnt [12]),
    .b(\PWM4/FreCnt [15]),
    .c(\PWM4/FreCntr [12]),
    .d(\PWM4/FreCntr [15]),
    .o(_al_u1440_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u1441 (
    .a(_al_u1437_o),
    .b(_al_u1439_o),
    .c(_al_u1440_o),
    .d(\PWM4/FreCnt [21]),
    .e(\PWM4/FreCntr [21]),
    .o(_al_u1441_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1442 (
    .a(\PWM4/FreCnt [7]),
    .b(\PWM4/FreCnt [9]),
    .c(\PWM4/FreCntr [7]),
    .d(\PWM4/FreCntr [9]),
    .o(_al_u1442_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1443 (
    .a(_al_u1442_o),
    .b(\PWM4/FreCnt [11]),
    .c(\PWM4/FreCnt [25]),
    .d(\PWM4/FreCntr [11]),
    .e(\PWM4/FreCntr [25]),
    .o(_al_u1443_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1444 (
    .a(\PWM4/FreCnt [2]),
    .b(\PWM4/FreCnt [3]),
    .c(\PWM4/FreCntr [2]),
    .d(\PWM4/FreCntr [3]),
    .o(_al_u1444_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1445 (
    .a(_al_u1444_o),
    .b(\PWM4/FreCnt [1]),
    .c(\PWM4/FreCnt [10]),
    .d(\PWM4/FreCntr [1]),
    .e(\PWM4/FreCntr [10]),
    .o(_al_u1445_o));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~(D*C*B*A))"),
    .INIT(32'hffff8000))
    _al_u1446 (
    .a(_al_u1435_o),
    .b(_al_u1441_o),
    .c(_al_u1443_o),
    .d(_al_u1445_o),
    .e(pwm_pad[4]),
    .o(\pwm[4]_d ));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1447 (
    .a(\PWM5/FreCnt [16]),
    .b(\PWM5/FreCnt [4]),
    .c(\PWM5/FreCntr [16]),
    .d(\PWM5/FreCntr [4]),
    .o(_al_u1447_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1448 (
    .a(_al_u1447_o),
    .b(\PWM5/FreCnt [18]),
    .c(\PWM5/FreCnt [5]),
    .d(\PWM5/FreCntr [18]),
    .e(\PWM5/FreCntr [5]),
    .o(_al_u1448_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1449 (
    .a(\PWM5/FreCnt [22]),
    .b(\PWM5/FreCnt [23]),
    .c(\PWM5/FreCntr [22]),
    .d(\PWM5/FreCntr [23]),
    .o(_al_u1449_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1450 (
    .a(_al_u1449_o),
    .b(\PWM5/FreCnt [17]),
    .c(\PWM5/FreCnt [8]),
    .d(\PWM5/FreCntr [17]),
    .e(\PWM5/FreCntr [8]),
    .o(_al_u1450_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1451 (
    .a(\PWM5/FreCnt [20]),
    .b(\PWM5/FreCnt [26]),
    .c(\PWM5/FreCntr [20]),
    .d(\PWM5/FreCntr [26]),
    .o(_al_u1451_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u1452 (
    .a(_al_u1448_o),
    .b(_al_u1450_o),
    .c(_al_u1451_o),
    .d(\PWM5/FreCnt [14]),
    .e(\PWM5/FreCntr [14]),
    .o(_al_u1452_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u1453 (
    .a(\PWM5/FreCnt [12]),
    .b(\PWM5/FreCnt [15]),
    .c(\PWM5/FreCntr [12]),
    .d(\PWM5/FreCntr [15]),
    .o(_al_u1453_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u1454 (
    .a(_al_u1453_o),
    .b(\PWM5/FreCnt [6]),
    .c(\PWM5/FreCntr [6]),
    .o(_al_u1454_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1455 (
    .a(\PWM5/FreCnt [0]),
    .b(\PWM5/FreCnt [24]),
    .c(\PWM5/FreCntr [0]),
    .d(\PWM5/FreCntr [24]),
    .o(_al_u1455_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1456 (
    .a(_al_u1455_o),
    .b(\PWM5/FreCnt [13]),
    .c(\PWM5/FreCnt [19]),
    .d(\PWM5/FreCntr [13]),
    .e(\PWM5/FreCntr [19]),
    .o(_al_u1456_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u1457 (
    .a(\PWM5/FreCnt [12]),
    .b(\PWM5/FreCnt [15]),
    .c(\PWM5/FreCntr [12]),
    .d(\PWM5/FreCntr [15]),
    .o(_al_u1457_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u1458 (
    .a(_al_u1454_o),
    .b(_al_u1456_o),
    .c(_al_u1457_o),
    .d(\PWM5/FreCnt [21]),
    .e(\PWM5/FreCntr [21]),
    .o(_al_u1458_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1459 (
    .a(\PWM5/FreCnt [7]),
    .b(\PWM5/FreCnt [9]),
    .c(\PWM5/FreCntr [7]),
    .d(\PWM5/FreCntr [9]),
    .o(_al_u1459_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1460 (
    .a(_al_u1459_o),
    .b(\PWM5/FreCnt [11]),
    .c(\PWM5/FreCnt [25]),
    .d(\PWM5/FreCntr [11]),
    .e(\PWM5/FreCntr [25]),
    .o(_al_u1460_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1461 (
    .a(\PWM5/FreCnt [2]),
    .b(\PWM5/FreCnt [3]),
    .c(\PWM5/FreCntr [2]),
    .d(\PWM5/FreCntr [3]),
    .o(_al_u1461_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1462 (
    .a(_al_u1461_o),
    .b(\PWM5/FreCnt [1]),
    .c(\PWM5/FreCnt [10]),
    .d(\PWM5/FreCntr [1]),
    .e(\PWM5/FreCntr [10]),
    .o(_al_u1462_o));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~(D*C*B*A))"),
    .INIT(32'hffff8000))
    _al_u1463 (
    .a(_al_u1452_o),
    .b(_al_u1458_o),
    .c(_al_u1460_o),
    .d(_al_u1462_o),
    .e(pwm_pad[5]),
    .o(\pwm[5]_d ));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1464 (
    .a(\PWM6/FreCnt [16]),
    .b(\PWM6/FreCnt [4]),
    .c(\PWM6/FreCntr [16]),
    .d(\PWM6/FreCntr [4]),
    .o(_al_u1464_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1465 (
    .a(_al_u1464_o),
    .b(\PWM6/FreCnt [18]),
    .c(\PWM6/FreCnt [5]),
    .d(\PWM6/FreCntr [18]),
    .e(\PWM6/FreCntr [5]),
    .o(_al_u1465_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1466 (
    .a(\PWM6/FreCnt [22]),
    .b(\PWM6/FreCnt [23]),
    .c(\PWM6/FreCntr [22]),
    .d(\PWM6/FreCntr [23]),
    .o(_al_u1466_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1467 (
    .a(_al_u1466_o),
    .b(\PWM6/FreCnt [24]),
    .c(\PWM6/FreCnt [7]),
    .d(\PWM6/FreCntr [24]),
    .e(\PWM6/FreCntr [7]),
    .o(_al_u1467_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1468 (
    .a(\PWM6/FreCnt [20]),
    .b(\PWM6/FreCnt [26]),
    .c(\PWM6/FreCntr [20]),
    .d(\PWM6/FreCntr [26]),
    .o(_al_u1468_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u1469 (
    .a(_al_u1465_o),
    .b(_al_u1467_o),
    .c(_al_u1468_o),
    .d(\PWM6/FreCnt [14]),
    .e(\PWM6/FreCntr [14]),
    .o(_al_u1469_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1470 (
    .a(\PWM6/FreCnt [1]),
    .b(\PWM6/FreCnt [21]),
    .c(\PWM6/FreCntr [1]),
    .d(\PWM6/FreCntr [21]),
    .o(_al_u1470_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1471 (
    .a(_al_u1470_o),
    .b(\PWM6/FreCnt [12]),
    .c(\PWM6/FreCnt [15]),
    .d(\PWM6/FreCntr [12]),
    .e(\PWM6/FreCntr [15]),
    .o(_al_u1471_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1472 (
    .a(\PWM6/FreCnt [0]),
    .b(\PWM6/FreCnt [10]),
    .c(\PWM6/FreCntr [0]),
    .d(\PWM6/FreCntr [10]),
    .o(_al_u1472_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1473 (
    .a(_al_u1472_o),
    .b(\PWM6/FreCnt [13]),
    .c(\PWM6/FreCnt [19]),
    .d(\PWM6/FreCntr [13]),
    .e(\PWM6/FreCntr [19]),
    .o(_al_u1473_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1474 (
    .a(\PWM6/FreCnt [17]),
    .b(\PWM6/FreCnt [9]),
    .c(\PWM6/FreCntr [17]),
    .d(\PWM6/FreCntr [9]),
    .o(_al_u1474_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1475 (
    .a(_al_u1474_o),
    .b(\PWM6/FreCnt [6]),
    .c(\PWM6/FreCnt [8]),
    .d(\PWM6/FreCntr [6]),
    .e(\PWM6/FreCntr [8]),
    .o(_al_u1475_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1476 (
    .a(\PWM6/FreCnt [11]),
    .b(\PWM6/FreCnt [25]),
    .c(\PWM6/FreCntr [11]),
    .d(\PWM6/FreCntr [25]),
    .o(_al_u1476_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1477 (
    .a(_al_u1476_o),
    .b(\PWM6/FreCnt [2]),
    .c(\PWM6/FreCnt [3]),
    .d(\PWM6/FreCntr [2]),
    .e(\PWM6/FreCntr [3]),
    .o(_al_u1477_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    _al_u1478 (
    .a(_al_u1469_o),
    .b(_al_u1471_o),
    .c(_al_u1473_o),
    .d(_al_u1475_o),
    .e(_al_u1477_o),
    .o(\PWM6/n18_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u1479 (
    .a(\PWM6/n18_lutinv ),
    .b(pwm_pad[6]),
    .o(\pwm[6]_d ));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1480 (
    .a(\PWM7/FreCnt [22]),
    .b(\PWM7/FreCnt [23]),
    .c(\PWM7/FreCntr [22]),
    .d(\PWM7/FreCntr [23]),
    .o(_al_u1480_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1481 (
    .a(_al_u1480_o),
    .b(\PWM7/FreCnt [17]),
    .c(\PWM7/FreCnt [8]),
    .d(\PWM7/FreCntr [17]),
    .e(\PWM7/FreCntr [8]),
    .o(_al_u1481_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1482 (
    .a(\PWM7/FreCnt [6]),
    .b(\PWM7/FreCnt [7]),
    .c(\PWM7/FreCntr [6]),
    .d(\PWM7/FreCntr [7]),
    .o(_al_u1482_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1483 (
    .a(_al_u1482_o),
    .b(\PWM7/FreCnt [4]),
    .c(\PWM7/FreCnt [9]),
    .d(\PWM7/FreCntr [4]),
    .e(\PWM7/FreCntr [9]),
    .o(_al_u1483_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1484 (
    .a(\PWM7/FreCnt [18]),
    .b(\PWM7/FreCnt [5]),
    .c(\PWM7/FreCntr [18]),
    .d(\PWM7/FreCntr [5]),
    .o(_al_u1484_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u1485 (
    .a(_al_u1481_o),
    .b(_al_u1483_o),
    .c(_al_u1484_o),
    .d(\PWM7/FreCnt [3]),
    .e(\PWM7/FreCntr [3]),
    .o(_al_u1485_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u1486 (
    .a(\PWM7/FreCnt [12]),
    .b(\PWM7/FreCnt [15]),
    .c(\PWM7/FreCntr [12]),
    .d(\PWM7/FreCntr [15]),
    .o(_al_u1486_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1487 (
    .a(\PWM7/FreCnt [10]),
    .b(\PWM7/FreCnt [2]),
    .c(\PWM7/FreCntr [10]),
    .d(\PWM7/FreCntr [2]),
    .o(_al_u1487_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D@C))"),
    .INIT(16'h8008))
    _al_u1488 (
    .a(_al_u1486_o),
    .b(_al_u1487_o),
    .c(\PWM7/FreCnt [21]),
    .d(\PWM7/FreCntr [21]),
    .o(_al_u1488_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1489 (
    .a(\PWM7/FreCnt [1]),
    .b(\PWM7/FreCntr [1]),
    .o(_al_u1489_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(E@C)*~(~D*B))"),
    .INIT(32'h50100501))
    _al_u1490 (
    .a(_al_u1489_o),
    .b(\PWM7/FreCnt [12]),
    .c(\PWM7/FreCnt [24]),
    .d(\PWM7/FreCntr [12]),
    .e(\PWM7/FreCntr [24]),
    .o(_al_u1490_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u1491 (
    .a(\PWM7/FreCnt [1]),
    .b(\PWM7/FreCnt [15]),
    .c(\PWM7/FreCntr [1]),
    .d(\PWM7/FreCntr [15]),
    .o(_al_u1491_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u1492 (
    .a(_al_u1488_o),
    .b(_al_u1490_o),
    .c(_al_u1491_o),
    .d(\PWM7/FreCnt [0]),
    .e(\PWM7/FreCntr [0]),
    .o(_al_u1492_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1493 (
    .a(\PWM7/FreCnt [11]),
    .b(\PWM7/FreCnt [25]),
    .c(\PWM7/FreCntr [11]),
    .d(\PWM7/FreCntr [25]),
    .o(_al_u1493_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1494 (
    .a(_al_u1493_o),
    .b(\PWM7/FreCnt [14]),
    .c(\PWM7/FreCnt [20]),
    .d(\PWM7/FreCntr [14]),
    .e(\PWM7/FreCntr [20]),
    .o(_al_u1494_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1495 (
    .a(\PWM7/FreCnt [16]),
    .b(\PWM7/FreCnt [26]),
    .c(\PWM7/FreCntr [16]),
    .d(\PWM7/FreCntr [26]),
    .o(_al_u1495_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1496 (
    .a(_al_u1495_o),
    .b(\PWM7/FreCnt [13]),
    .c(\PWM7/FreCnt [19]),
    .d(\PWM7/FreCntr [13]),
    .e(\PWM7/FreCntr [19]),
    .o(_al_u1496_o));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~(D*C*B*A))"),
    .INIT(32'hffff8000))
    _al_u1497 (
    .a(_al_u1485_o),
    .b(_al_u1492_o),
    .c(_al_u1494_o),
    .d(_al_u1496_o),
    .e(pwm_pad[7]),
    .o(\pwm[7]_d ));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1498 (
    .a(\PWM8/FreCnt [22]),
    .b(\PWM8/FreCnt [23]),
    .c(\PWM8/FreCntr [22]),
    .d(\PWM8/FreCntr [23]),
    .o(_al_u1498_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1499 (
    .a(_al_u1498_o),
    .b(\PWM8/FreCnt [17]),
    .c(\PWM8/FreCnt [8]),
    .d(\PWM8/FreCntr [17]),
    .e(\PWM8/FreCntr [8]),
    .o(_al_u1499_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1500 (
    .a(\PWM8/FreCnt [6]),
    .b(\PWM8/FreCnt [7]),
    .c(\PWM8/FreCntr [6]),
    .d(\PWM8/FreCntr [7]),
    .o(_al_u1500_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1501 (
    .a(_al_u1500_o),
    .b(\PWM8/FreCnt [4]),
    .c(\PWM8/FreCnt [9]),
    .d(\PWM8/FreCntr [4]),
    .e(\PWM8/FreCntr [9]),
    .o(_al_u1501_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1502 (
    .a(\PWM8/FreCnt [18]),
    .b(\PWM8/FreCnt [5]),
    .c(\PWM8/FreCntr [18]),
    .d(\PWM8/FreCntr [5]),
    .o(_al_u1502_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u1503 (
    .a(_al_u1499_o),
    .b(_al_u1501_o),
    .c(_al_u1502_o),
    .d(\PWM8/FreCnt [3]),
    .e(\PWM8/FreCntr [3]),
    .o(_al_u1503_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u1504 (
    .a(\PWM8/FreCnt [12]),
    .b(\PWM8/FreCnt [15]),
    .c(\PWM8/FreCntr [12]),
    .d(\PWM8/FreCntr [15]),
    .o(_al_u1504_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1505 (
    .a(\PWM8/FreCnt [10]),
    .b(\PWM8/FreCnt [2]),
    .c(\PWM8/FreCntr [10]),
    .d(\PWM8/FreCntr [2]),
    .o(_al_u1505_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D@C))"),
    .INIT(16'h8008))
    _al_u1506 (
    .a(_al_u1504_o),
    .b(_al_u1505_o),
    .c(\PWM8/FreCnt [21]),
    .d(\PWM8/FreCntr [21]),
    .o(_al_u1506_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1507 (
    .a(\PWM8/FreCnt [1]),
    .b(\PWM8/FreCntr [1]),
    .o(_al_u1507_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(E@C)*~(~D*B))"),
    .INIT(32'h50100501))
    _al_u1508 (
    .a(_al_u1507_o),
    .b(\PWM8/FreCnt [12]),
    .c(\PWM8/FreCnt [24]),
    .d(\PWM8/FreCntr [12]),
    .e(\PWM8/FreCntr [24]),
    .o(_al_u1508_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u1509 (
    .a(\PWM8/FreCnt [1]),
    .b(\PWM8/FreCnt [15]),
    .c(\PWM8/FreCntr [1]),
    .d(\PWM8/FreCntr [15]),
    .o(_al_u1509_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u1510 (
    .a(_al_u1506_o),
    .b(_al_u1508_o),
    .c(_al_u1509_o),
    .d(\PWM8/FreCnt [0]),
    .e(\PWM8/FreCntr [0]),
    .o(_al_u1510_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1511 (
    .a(\PWM8/FreCnt [11]),
    .b(\PWM8/FreCnt [25]),
    .c(\PWM8/FreCntr [11]),
    .d(\PWM8/FreCntr [25]),
    .o(_al_u1511_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1512 (
    .a(_al_u1511_o),
    .b(\PWM8/FreCnt [14]),
    .c(\PWM8/FreCnt [20]),
    .d(\PWM8/FreCntr [14]),
    .e(\PWM8/FreCntr [20]),
    .o(_al_u1512_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1513 (
    .a(\PWM8/FreCnt [16]),
    .b(\PWM8/FreCnt [26]),
    .c(\PWM8/FreCntr [16]),
    .d(\PWM8/FreCntr [26]),
    .o(_al_u1513_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1514 (
    .a(_al_u1513_o),
    .b(\PWM8/FreCnt [13]),
    .c(\PWM8/FreCnt [19]),
    .d(\PWM8/FreCntr [13]),
    .e(\PWM8/FreCntr [19]),
    .o(_al_u1514_o));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~(D*C*B*A))"),
    .INIT(32'hffff8000))
    _al_u1515 (
    .a(_al_u1503_o),
    .b(_al_u1510_o),
    .c(_al_u1512_o),
    .d(_al_u1514_o),
    .e(pwm_pad[8]),
    .o(\pwm[8]_d ));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1516 (
    .a(\PWM9/FreCnt [16]),
    .b(\PWM9/FreCnt [3]),
    .c(\PWM9/FreCntr [16]),
    .d(\PWM9/FreCntr [3]),
    .o(_al_u1516_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1517 (
    .a(_al_u1516_o),
    .b(\PWM9/FreCnt [18]),
    .c(\PWM9/FreCnt [5]),
    .d(\PWM9/FreCntr [18]),
    .e(\PWM9/FreCntr [5]),
    .o(_al_u1517_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1518 (
    .a(\PWM9/FreCnt [22]),
    .b(\PWM9/FreCnt [23]),
    .c(\PWM9/FreCntr [22]),
    .d(\PWM9/FreCntr [23]),
    .o(_al_u1518_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1519 (
    .a(_al_u1518_o),
    .b(\PWM9/FreCnt [17]),
    .c(\PWM9/FreCnt [8]),
    .d(\PWM9/FreCntr [17]),
    .e(\PWM9/FreCntr [8]),
    .o(_al_u1519_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1520 (
    .a(\PWM9/FreCnt [20]),
    .b(\PWM9/FreCnt [26]),
    .c(\PWM9/FreCntr [20]),
    .d(\PWM9/FreCntr [26]),
    .o(_al_u1520_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u1521 (
    .a(_al_u1517_o),
    .b(_al_u1519_o),
    .c(_al_u1520_o),
    .d(\PWM9/FreCnt [14]),
    .e(\PWM9/FreCntr [14]),
    .o(_al_u1521_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u1522 (
    .a(\PWM9/FreCnt [12]),
    .b(\PWM9/FreCnt [15]),
    .c(\PWM9/FreCntr [12]),
    .d(\PWM9/FreCntr [15]),
    .o(_al_u1522_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u1523 (
    .a(_al_u1522_o),
    .b(\PWM9/FreCnt [6]),
    .c(\PWM9/FreCntr [6]),
    .o(_al_u1523_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1524 (
    .a(\PWM9/FreCnt [0]),
    .b(\PWM9/FreCnt [24]),
    .c(\PWM9/FreCntr [0]),
    .d(\PWM9/FreCntr [24]),
    .o(_al_u1524_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1525 (
    .a(_al_u1524_o),
    .b(\PWM9/FreCnt [13]),
    .c(\PWM9/FreCnt [19]),
    .d(\PWM9/FreCntr [13]),
    .e(\PWM9/FreCntr [19]),
    .o(_al_u1525_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u1526 (
    .a(\PWM9/FreCnt [12]),
    .b(\PWM9/FreCnt [15]),
    .c(\PWM9/FreCntr [12]),
    .d(\PWM9/FreCntr [15]),
    .o(_al_u1526_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u1527 (
    .a(_al_u1523_o),
    .b(_al_u1525_o),
    .c(_al_u1526_o),
    .d(\PWM9/FreCnt [21]),
    .e(\PWM9/FreCntr [21]),
    .o(_al_u1527_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1528 (
    .a(\PWM9/FreCnt [7]),
    .b(\PWM9/FreCnt [9]),
    .c(\PWM9/FreCntr [7]),
    .d(\PWM9/FreCntr [9]),
    .o(_al_u1528_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1529 (
    .a(_al_u1528_o),
    .b(\PWM9/FreCnt [11]),
    .c(\PWM9/FreCnt [4]),
    .d(\PWM9/FreCntr [11]),
    .e(\PWM9/FreCntr [4]),
    .o(_al_u1529_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1530 (
    .a(\PWM9/FreCnt [2]),
    .b(\PWM9/FreCnt [25]),
    .c(\PWM9/FreCntr [2]),
    .d(\PWM9/FreCntr [25]),
    .o(_al_u1530_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1531 (
    .a(_al_u1530_o),
    .b(\PWM9/FreCnt [1]),
    .c(\PWM9/FreCnt [10]),
    .d(\PWM9/FreCntr [1]),
    .e(\PWM9/FreCntr [10]),
    .o(_al_u1531_o));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~(D*C*B*A))"),
    .INIT(32'hffff8000))
    _al_u1532 (
    .a(_al_u1521_o),
    .b(_al_u1527_o),
    .c(_al_u1529_o),
    .d(_al_u1531_o),
    .e(pwm_pad[9]),
    .o(\pwm[9]_d ));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1533 (
    .a(\PWMA/FreCnt [22]),
    .b(\PWMA/FreCnt [23]),
    .c(\PWMA/FreCntr [22]),
    .d(\PWMA/FreCntr [23]),
    .o(_al_u1533_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1534 (
    .a(_al_u1533_o),
    .b(\PWMA/FreCnt [17]),
    .c(\PWMA/FreCnt [8]),
    .d(\PWMA/FreCntr [17]),
    .e(\PWMA/FreCntr [8]),
    .o(_al_u1534_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1535 (
    .a(\PWMA/FreCnt [6]),
    .b(\PWMA/FreCnt [7]),
    .c(\PWMA/FreCntr [6]),
    .d(\PWMA/FreCntr [7]),
    .o(_al_u1535_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1536 (
    .a(_al_u1535_o),
    .b(\PWMA/FreCnt [11]),
    .c(\PWMA/FreCnt [9]),
    .d(\PWMA/FreCntr [11]),
    .e(\PWMA/FreCntr [9]),
    .o(_al_u1536_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1537 (
    .a(\PWMA/FreCnt [18]),
    .b(\PWMA/FreCnt [5]),
    .c(\PWMA/FreCntr [18]),
    .d(\PWMA/FreCntr [5]),
    .o(_al_u1537_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u1538 (
    .a(_al_u1534_o),
    .b(_al_u1536_o),
    .c(_al_u1537_o),
    .d(\PWMA/FreCnt [4]),
    .e(\PWMA/FreCntr [4]),
    .o(_al_u1538_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u1539 (
    .a(\PWMA/FreCnt [12]),
    .b(\PWMA/FreCnt [15]),
    .c(\PWMA/FreCntr [12]),
    .d(\PWMA/FreCntr [15]),
    .o(_al_u1539_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1540 (
    .a(\PWMA/FreCnt [10]),
    .b(\PWMA/FreCnt [3]),
    .c(\PWMA/FreCntr [10]),
    .d(\PWMA/FreCntr [3]),
    .o(_al_u1540_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D@C))"),
    .INIT(16'h8008))
    _al_u1541 (
    .a(_al_u1539_o),
    .b(_al_u1540_o),
    .c(\PWMA/FreCnt [21]),
    .d(\PWMA/FreCntr [21]),
    .o(_al_u1541_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1542 (
    .a(\PWMA/FreCnt [1]),
    .b(\PWMA/FreCntr [1]),
    .o(_al_u1542_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(E@C)*~(~D*B))"),
    .INIT(32'h50100501))
    _al_u1543 (
    .a(_al_u1542_o),
    .b(\PWMA/FreCnt [12]),
    .c(\PWMA/FreCnt [24]),
    .d(\PWMA/FreCntr [12]),
    .e(\PWMA/FreCntr [24]),
    .o(_al_u1543_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u1544 (
    .a(\PWMA/FreCnt [1]),
    .b(\PWMA/FreCnt [15]),
    .c(\PWMA/FreCntr [1]),
    .d(\PWMA/FreCntr [15]),
    .o(_al_u1544_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u1545 (
    .a(_al_u1541_o),
    .b(_al_u1543_o),
    .c(_al_u1544_o),
    .d(\PWMA/FreCnt [0]),
    .e(\PWMA/FreCntr [0]),
    .o(_al_u1545_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1546 (
    .a(\PWMA/FreCnt [14]),
    .b(\PWMA/FreCnt [25]),
    .c(\PWMA/FreCntr [14]),
    .d(\PWMA/FreCntr [25]),
    .o(_al_u1546_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1547 (
    .a(_al_u1546_o),
    .b(\PWMA/FreCnt [20]),
    .c(\PWMA/FreCnt [26]),
    .d(\PWMA/FreCntr [20]),
    .e(\PWMA/FreCntr [26]),
    .o(_al_u1547_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1548 (
    .a(\PWMA/FreCnt [13]),
    .b(\PWMA/FreCnt [16]),
    .c(\PWMA/FreCntr [13]),
    .d(\PWMA/FreCntr [16]),
    .o(_al_u1548_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1549 (
    .a(_al_u1548_o),
    .b(\PWMA/FreCnt [19]),
    .c(\PWMA/FreCnt [2]),
    .d(\PWMA/FreCntr [19]),
    .e(\PWMA/FreCntr [2]),
    .o(_al_u1549_o));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~(D*C*B*A))"),
    .INIT(32'hffff8000))
    _al_u1550 (
    .a(_al_u1538_o),
    .b(_al_u1545_o),
    .c(_al_u1547_o),
    .d(_al_u1549_o),
    .e(pwm_pad[10]),
    .o(\pwm[10]_d ));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1551 (
    .a(\PWMB/FreCnt [16]),
    .b(\PWMB/FreCnt [3]),
    .c(\PWMB/FreCntr [16]),
    .d(\PWMB/FreCntr [3]),
    .o(_al_u1551_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1552 (
    .a(_al_u1551_o),
    .b(\PWMB/FreCnt [18]),
    .c(\PWMB/FreCnt [5]),
    .d(\PWMB/FreCntr [18]),
    .e(\PWMB/FreCntr [5]),
    .o(_al_u1552_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1553 (
    .a(\PWMB/FreCnt [22]),
    .b(\PWMB/FreCnt [23]),
    .c(\PWMB/FreCntr [22]),
    .d(\PWMB/FreCntr [23]),
    .o(_al_u1553_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1554 (
    .a(_al_u1553_o),
    .b(\PWMB/FreCnt [17]),
    .c(\PWMB/FreCnt [8]),
    .d(\PWMB/FreCntr [17]),
    .e(\PWMB/FreCntr [8]),
    .o(_al_u1554_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1555 (
    .a(\PWMB/FreCnt [20]),
    .b(\PWMB/FreCnt [26]),
    .c(\PWMB/FreCntr [20]),
    .d(\PWMB/FreCntr [26]),
    .o(_al_u1555_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u1556 (
    .a(_al_u1552_o),
    .b(_al_u1554_o),
    .c(_al_u1555_o),
    .d(\PWMB/FreCnt [14]),
    .e(\PWMB/FreCntr [14]),
    .o(_al_u1556_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u1557 (
    .a(\PWMB/FreCnt [12]),
    .b(\PWMB/FreCnt [15]),
    .c(\PWMB/FreCntr [12]),
    .d(\PWMB/FreCntr [15]),
    .o(_al_u1557_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u1558 (
    .a(_al_u1557_o),
    .b(\PWMB/FreCnt [6]),
    .c(\PWMB/FreCntr [6]),
    .o(_al_u1558_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1559 (
    .a(\PWMB/FreCnt [0]),
    .b(\PWMB/FreCnt [24]),
    .c(\PWMB/FreCntr [0]),
    .d(\PWMB/FreCntr [24]),
    .o(_al_u1559_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1560 (
    .a(_al_u1559_o),
    .b(\PWMB/FreCnt [13]),
    .c(\PWMB/FreCnt [19]),
    .d(\PWMB/FreCntr [13]),
    .e(\PWMB/FreCntr [19]),
    .o(_al_u1560_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u1561 (
    .a(\PWMB/FreCnt [12]),
    .b(\PWMB/FreCnt [15]),
    .c(\PWMB/FreCntr [12]),
    .d(\PWMB/FreCntr [15]),
    .o(_al_u1561_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u1562 (
    .a(_al_u1558_o),
    .b(_al_u1560_o),
    .c(_al_u1561_o),
    .d(\PWMB/FreCnt [21]),
    .e(\PWMB/FreCntr [21]),
    .o(_al_u1562_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1563 (
    .a(\PWMB/FreCnt [7]),
    .b(\PWMB/FreCnt [9]),
    .c(\PWMB/FreCntr [7]),
    .d(\PWMB/FreCntr [9]),
    .o(_al_u1563_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1564 (
    .a(_al_u1563_o),
    .b(\PWMB/FreCnt [11]),
    .c(\PWMB/FreCnt [4]),
    .d(\PWMB/FreCntr [11]),
    .e(\PWMB/FreCntr [4]),
    .o(_al_u1564_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1565 (
    .a(\PWMB/FreCnt [2]),
    .b(\PWMB/FreCnt [25]),
    .c(\PWMB/FreCntr [2]),
    .d(\PWMB/FreCntr [25]),
    .o(_al_u1565_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1566 (
    .a(_al_u1565_o),
    .b(\PWMB/FreCnt [1]),
    .c(\PWMB/FreCnt [10]),
    .d(\PWMB/FreCntr [1]),
    .e(\PWMB/FreCntr [10]),
    .o(_al_u1566_o));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~(D*C*B*A))"),
    .INIT(32'hffff8000))
    _al_u1567 (
    .a(_al_u1556_o),
    .b(_al_u1562_o),
    .c(_al_u1564_o),
    .d(_al_u1566_o),
    .e(pwm_pad[11]),
    .o(\pwm[11]_d ));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1568 (
    .a(\PWMC/FreCnt [16]),
    .b(\PWMC/FreCnt [4]),
    .c(\PWMC/FreCntr [16]),
    .d(\PWMC/FreCntr [4]),
    .o(_al_u1568_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1569 (
    .a(_al_u1568_o),
    .b(\PWMC/FreCnt [18]),
    .c(\PWMC/FreCnt [5]),
    .d(\PWMC/FreCntr [18]),
    .e(\PWMC/FreCntr [5]),
    .o(_al_u1569_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1570 (
    .a(\PWMC/FreCnt [22]),
    .b(\PWMC/FreCnt [23]),
    .c(\PWMC/FreCntr [22]),
    .d(\PWMC/FreCntr [23]),
    .o(_al_u1570_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1571 (
    .a(_al_u1570_o),
    .b(\PWMC/FreCnt [7]),
    .c(\PWMC/FreCnt [9]),
    .d(\PWMC/FreCntr [7]),
    .e(\PWMC/FreCntr [9]),
    .o(_al_u1571_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1572 (
    .a(\PWMC/FreCnt [20]),
    .b(\PWMC/FreCnt [26]),
    .c(\PWMC/FreCntr [20]),
    .d(\PWMC/FreCntr [26]),
    .o(_al_u1572_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u1573 (
    .a(_al_u1569_o),
    .b(_al_u1571_o),
    .c(_al_u1572_o),
    .d(\PWMC/FreCnt [14]),
    .e(\PWMC/FreCntr [14]),
    .o(_al_u1573_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u1574 (
    .a(\PWMC/FreCnt [15]),
    .b(\PWMC/FreCnt [21]),
    .c(\PWMC/FreCntr [15]),
    .d(\PWMC/FreCntr [21]),
    .o(_al_u1574_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u1575 (
    .a(_al_u1574_o),
    .b(\PWMC/FreCnt [1]),
    .c(\PWMC/FreCntr [1]),
    .o(_al_u1575_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1576 (
    .a(\PWMC/FreCnt [0]),
    .b(\PWMC/FreCnt [10]),
    .c(\PWMC/FreCntr [0]),
    .d(\PWMC/FreCntr [10]),
    .o(_al_u1576_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1577 (
    .a(_al_u1576_o),
    .b(\PWMC/FreCnt [13]),
    .c(\PWMC/FreCnt [19]),
    .d(\PWMC/FreCntr [13]),
    .e(\PWMC/FreCntr [19]),
    .o(_al_u1577_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u1578 (
    .a(\PWMC/FreCnt [15]),
    .b(\PWMC/FreCnt [21]),
    .c(\PWMC/FreCntr [15]),
    .d(\PWMC/FreCntr [21]),
    .o(_al_u1578_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u1579 (
    .a(_al_u1575_o),
    .b(_al_u1577_o),
    .c(_al_u1578_o),
    .d(\PWMC/FreCnt [12]),
    .e(\PWMC/FreCntr [12]),
    .o(_al_u1579_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1580 (
    .a(\PWMC/FreCnt [17]),
    .b(\PWMC/FreCnt [6]),
    .c(\PWMC/FreCntr [17]),
    .d(\PWMC/FreCntr [6]),
    .o(_al_u1580_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1581 (
    .a(_al_u1580_o),
    .b(\PWMC/FreCnt [24]),
    .c(\PWMC/FreCnt [8]),
    .d(\PWMC/FreCntr [24]),
    .e(\PWMC/FreCntr [8]),
    .o(_al_u1581_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1582 (
    .a(\PWMC/FreCnt [11]),
    .b(\PWMC/FreCnt [25]),
    .c(\PWMC/FreCntr [11]),
    .d(\PWMC/FreCntr [25]),
    .o(_al_u1582_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1583 (
    .a(_al_u1582_o),
    .b(\PWMC/FreCnt [2]),
    .c(\PWMC/FreCnt [3]),
    .d(\PWMC/FreCntr [2]),
    .e(\PWMC/FreCntr [3]),
    .o(_al_u1583_o));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~(D*C*B*A))"),
    .INIT(32'hffff8000))
    _al_u1584 (
    .a(_al_u1573_o),
    .b(_al_u1579_o),
    .c(_al_u1581_o),
    .d(_al_u1583_o),
    .e(pwm_pad[12]),
    .o(\pwm[12]_d ));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1585 (
    .a(\PWMD/FreCnt [16]),
    .b(\PWMD/FreCnt [4]),
    .c(\PWMD/FreCntr [16]),
    .d(\PWMD/FreCntr [4]),
    .o(_al_u1585_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1586 (
    .a(_al_u1585_o),
    .b(\PWMD/FreCnt [18]),
    .c(\PWMD/FreCnt [5]),
    .d(\PWMD/FreCntr [18]),
    .e(\PWMD/FreCntr [5]),
    .o(_al_u1586_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1587 (
    .a(\PWMD/FreCnt [22]),
    .b(\PWMD/FreCnt [23]),
    .c(\PWMD/FreCntr [22]),
    .d(\PWMD/FreCntr [23]),
    .o(_al_u1587_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1588 (
    .a(_al_u1587_o),
    .b(\PWMD/FreCnt [17]),
    .c(\PWMD/FreCnt [8]),
    .d(\PWMD/FreCntr [17]),
    .e(\PWMD/FreCntr [8]),
    .o(_al_u1588_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1589 (
    .a(\PWMD/FreCnt [20]),
    .b(\PWMD/FreCnt [26]),
    .c(\PWMD/FreCntr [20]),
    .d(\PWMD/FreCntr [26]),
    .o(_al_u1589_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u1590 (
    .a(_al_u1586_o),
    .b(_al_u1588_o),
    .c(_al_u1589_o),
    .d(\PWMD/FreCnt [14]),
    .e(\PWMD/FreCntr [14]),
    .o(_al_u1590_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u1591 (
    .a(\PWMD/FreCnt [12]),
    .b(\PWMD/FreCnt [15]),
    .c(\PWMD/FreCntr [12]),
    .d(\PWMD/FreCntr [15]),
    .o(_al_u1591_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u1592 (
    .a(_al_u1591_o),
    .b(\PWMD/FreCnt [6]),
    .c(\PWMD/FreCntr [6]),
    .o(_al_u1592_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1593 (
    .a(\PWMD/FreCnt [0]),
    .b(\PWMD/FreCnt [24]),
    .c(\PWMD/FreCntr [0]),
    .d(\PWMD/FreCntr [24]),
    .o(_al_u1593_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1594 (
    .a(_al_u1593_o),
    .b(\PWMD/FreCnt [13]),
    .c(\PWMD/FreCnt [19]),
    .d(\PWMD/FreCntr [13]),
    .e(\PWMD/FreCntr [19]),
    .o(_al_u1594_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u1595 (
    .a(\PWMD/FreCnt [12]),
    .b(\PWMD/FreCnt [15]),
    .c(\PWMD/FreCntr [12]),
    .d(\PWMD/FreCntr [15]),
    .o(_al_u1595_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u1596 (
    .a(_al_u1592_o),
    .b(_al_u1594_o),
    .c(_al_u1595_o),
    .d(\PWMD/FreCnt [21]),
    .e(\PWMD/FreCntr [21]),
    .o(_al_u1596_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1597 (
    .a(\PWMD/FreCnt [7]),
    .b(\PWMD/FreCnt [9]),
    .c(\PWMD/FreCntr [7]),
    .d(\PWMD/FreCntr [9]),
    .o(_al_u1597_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1598 (
    .a(_al_u1597_o),
    .b(\PWMD/FreCnt [11]),
    .c(\PWMD/FreCnt [25]),
    .d(\PWMD/FreCntr [11]),
    .e(\PWMD/FreCntr [25]),
    .o(_al_u1598_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1599 (
    .a(\PWMD/FreCnt [2]),
    .b(\PWMD/FreCnt [3]),
    .c(\PWMD/FreCntr [2]),
    .d(\PWMD/FreCntr [3]),
    .o(_al_u1599_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1600 (
    .a(_al_u1599_o),
    .b(\PWMD/FreCnt [1]),
    .c(\PWMD/FreCnt [10]),
    .d(\PWMD/FreCntr [1]),
    .e(\PWMD/FreCntr [10]),
    .o(_al_u1600_o));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~(D*C*B*A))"),
    .INIT(32'hffff8000))
    _al_u1601 (
    .a(_al_u1590_o),
    .b(_al_u1596_o),
    .c(_al_u1598_o),
    .d(_al_u1600_o),
    .e(pwm_pad[13]),
    .o(\pwm[13]_d ));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1602 (
    .a(\PWME/FreCnt [22]),
    .b(\PWME/FreCnt [23]),
    .c(\PWME/FreCntr [22]),
    .d(\PWME/FreCntr [23]),
    .o(_al_u1602_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1603 (
    .a(_al_u1602_o),
    .b(\PWME/FreCnt [17]),
    .c(\PWME/FreCnt [8]),
    .d(\PWME/FreCntr [17]),
    .e(\PWME/FreCntr [8]),
    .o(_al_u1603_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1604 (
    .a(\PWME/FreCnt [6]),
    .b(\PWME/FreCnt [7]),
    .c(\PWME/FreCntr [6]),
    .d(\PWME/FreCntr [7]),
    .o(_al_u1604_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1605 (
    .a(_al_u1604_o),
    .b(\PWME/FreCnt [11]),
    .c(\PWME/FreCnt [9]),
    .d(\PWME/FreCntr [11]),
    .e(\PWME/FreCntr [9]),
    .o(_al_u1605_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1606 (
    .a(\PWME/FreCnt [18]),
    .b(\PWME/FreCnt [5]),
    .c(\PWME/FreCntr [18]),
    .d(\PWME/FreCntr [5]),
    .o(_al_u1606_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u1607 (
    .a(_al_u1603_o),
    .b(_al_u1605_o),
    .c(_al_u1606_o),
    .d(\PWME/FreCnt [4]),
    .e(\PWME/FreCntr [4]),
    .o(_al_u1607_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u1608 (
    .a(\PWME/FreCnt [12]),
    .b(\PWME/FreCnt [15]),
    .c(\PWME/FreCntr [12]),
    .d(\PWME/FreCntr [15]),
    .o(_al_u1608_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1609 (
    .a(\PWME/FreCnt [10]),
    .b(\PWME/FreCnt [3]),
    .c(\PWME/FreCntr [10]),
    .d(\PWME/FreCntr [3]),
    .o(_al_u1609_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D@C))"),
    .INIT(16'h8008))
    _al_u1610 (
    .a(_al_u1608_o),
    .b(_al_u1609_o),
    .c(\PWME/FreCnt [21]),
    .d(\PWME/FreCntr [21]),
    .o(_al_u1610_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1611 (
    .a(\PWME/FreCnt [1]),
    .b(\PWME/FreCntr [1]),
    .o(_al_u1611_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(E@C)*~(~D*B))"),
    .INIT(32'h50100501))
    _al_u1612 (
    .a(_al_u1611_o),
    .b(\PWME/FreCnt [12]),
    .c(\PWME/FreCnt [24]),
    .d(\PWME/FreCntr [12]),
    .e(\PWME/FreCntr [24]),
    .o(_al_u1612_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u1613 (
    .a(\PWME/FreCnt [1]),
    .b(\PWME/FreCnt [15]),
    .c(\PWME/FreCntr [1]),
    .d(\PWME/FreCntr [15]),
    .o(_al_u1613_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u1614 (
    .a(_al_u1610_o),
    .b(_al_u1612_o),
    .c(_al_u1613_o),
    .d(\PWME/FreCnt [0]),
    .e(\PWME/FreCntr [0]),
    .o(_al_u1614_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1615 (
    .a(\PWME/FreCnt [14]),
    .b(\PWME/FreCnt [25]),
    .c(\PWME/FreCntr [14]),
    .d(\PWME/FreCntr [25]),
    .o(_al_u1615_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1616 (
    .a(_al_u1615_o),
    .b(\PWME/FreCnt [20]),
    .c(\PWME/FreCnt [26]),
    .d(\PWME/FreCntr [20]),
    .e(\PWME/FreCntr [26]),
    .o(_al_u1616_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1617 (
    .a(\PWME/FreCnt [13]),
    .b(\PWME/FreCnt [16]),
    .c(\PWME/FreCntr [13]),
    .d(\PWME/FreCntr [16]),
    .o(_al_u1617_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1618 (
    .a(_al_u1617_o),
    .b(\PWME/FreCnt [19]),
    .c(\PWME/FreCnt [2]),
    .d(\PWME/FreCntr [19]),
    .e(\PWME/FreCntr [2]),
    .o(_al_u1618_o));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~(D*C*B*A))"),
    .INIT(32'hffff8000))
    _al_u1619 (
    .a(_al_u1607_o),
    .b(_al_u1614_o),
    .c(_al_u1616_o),
    .d(_al_u1618_o),
    .e(pwm_pad[14]),
    .o(\pwm[14]_d ));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1620 (
    .a(\PWMF/FreCnt [22]),
    .b(\PWMF/FreCnt [23]),
    .c(\PWMF/FreCntr [22]),
    .d(\PWMF/FreCntr [23]),
    .o(_al_u1620_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1621 (
    .a(_al_u1620_o),
    .b(\PWMF/FreCnt [17]),
    .c(\PWMF/FreCnt [8]),
    .d(\PWMF/FreCntr [17]),
    .e(\PWMF/FreCntr [8]),
    .o(_al_u1621_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1622 (
    .a(\PWMF/FreCnt [6]),
    .b(\PWMF/FreCnt [7]),
    .c(\PWMF/FreCntr [6]),
    .d(\PWMF/FreCntr [7]),
    .o(_al_u1622_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1623 (
    .a(_al_u1622_o),
    .b(\PWMF/FreCnt [4]),
    .c(\PWMF/FreCnt [9]),
    .d(\PWMF/FreCntr [4]),
    .e(\PWMF/FreCntr [9]),
    .o(_al_u1623_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1624 (
    .a(\PWMF/FreCnt [18]),
    .b(\PWMF/FreCnt [5]),
    .c(\PWMF/FreCntr [18]),
    .d(\PWMF/FreCntr [5]),
    .o(_al_u1624_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u1625 (
    .a(_al_u1621_o),
    .b(_al_u1623_o),
    .c(_al_u1624_o),
    .d(\PWMF/FreCnt [3]),
    .e(\PWMF/FreCntr [3]),
    .o(_al_u1625_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u1626 (
    .a(\PWMF/FreCnt [12]),
    .b(\PWMF/FreCnt [15]),
    .c(\PWMF/FreCntr [12]),
    .d(\PWMF/FreCntr [15]),
    .o(_al_u1626_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1627 (
    .a(\PWMF/FreCnt [10]),
    .b(\PWMF/FreCnt [2]),
    .c(\PWMF/FreCntr [10]),
    .d(\PWMF/FreCntr [2]),
    .o(_al_u1627_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D@C))"),
    .INIT(16'h8008))
    _al_u1628 (
    .a(_al_u1626_o),
    .b(_al_u1627_o),
    .c(\PWMF/FreCnt [21]),
    .d(\PWMF/FreCntr [21]),
    .o(_al_u1628_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1629 (
    .a(\PWMF/FreCnt [1]),
    .b(\PWMF/FreCntr [1]),
    .o(_al_u1629_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(E@C)*~(~D*B))"),
    .INIT(32'h50100501))
    _al_u1630 (
    .a(_al_u1629_o),
    .b(\PWMF/FreCnt [12]),
    .c(\PWMF/FreCnt [24]),
    .d(\PWMF/FreCntr [12]),
    .e(\PWMF/FreCntr [24]),
    .o(_al_u1630_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u1631 (
    .a(\PWMF/FreCnt [1]),
    .b(\PWMF/FreCnt [15]),
    .c(\PWMF/FreCntr [1]),
    .d(\PWMF/FreCntr [15]),
    .o(_al_u1631_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u1632 (
    .a(_al_u1628_o),
    .b(_al_u1630_o),
    .c(_al_u1631_o),
    .d(\PWMF/FreCnt [0]),
    .e(\PWMF/FreCntr [0]),
    .o(_al_u1632_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1633 (
    .a(\PWMF/FreCnt [11]),
    .b(\PWMF/FreCnt [25]),
    .c(\PWMF/FreCntr [11]),
    .d(\PWMF/FreCntr [25]),
    .o(_al_u1633_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1634 (
    .a(_al_u1633_o),
    .b(\PWMF/FreCnt [14]),
    .c(\PWMF/FreCnt [20]),
    .d(\PWMF/FreCntr [14]),
    .e(\PWMF/FreCntr [20]),
    .o(_al_u1634_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1635 (
    .a(\PWMF/FreCnt [16]),
    .b(\PWMF/FreCnt [26]),
    .c(\PWMF/FreCntr [16]),
    .d(\PWMF/FreCntr [26]),
    .o(_al_u1635_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1636 (
    .a(_al_u1635_o),
    .b(\PWMF/FreCnt [13]),
    .c(\PWMF/FreCnt [19]),
    .d(\PWMF/FreCntr [13]),
    .e(\PWMF/FreCntr [19]),
    .o(_al_u1636_o));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~(D*C*B*A))"),
    .INIT(32'hffff8000))
    _al_u1637 (
    .a(_al_u1625_o),
    .b(_al_u1632_o),
    .c(_al_u1634_o),
    .d(_al_u1636_o),
    .e(pwm_pad[15]),
    .o(\pwm[15]_d ));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*~A)"),
    .INIT(32'h00000001))
    _al_u1638 (
    .a(timer[28]),
    .b(timer[29]),
    .c(timer[30]),
    .d(timer[31]),
    .e(timer[9]),
    .o(_al_u1638_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1639 (
    .a(timer[20]),
    .b(timer[21]),
    .c(timer[22]),
    .d(timer[23]),
    .o(_al_u1639_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*B*A)"),
    .INIT(32'h00000008))
    _al_u1640 (
    .a(_al_u1638_o),
    .b(_al_u1639_o),
    .c(timer[10]),
    .d(timer[11]),
    .e(timer[8]),
    .o(_al_u1640_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1641 (
    .a(timer[0]),
    .b(timer[1]),
    .c(timer[2]),
    .d(timer[3]),
    .o(_al_u1641_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*D*C*B*A)"),
    .INIT(32'h00008000))
    _al_u1642 (
    .a(_al_u1641_o),
    .b(timer[4]),
    .c(timer[5]),
    .d(timer[6]),
    .e(timer[7]),
    .o(_al_u1642_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u1643 (
    .a(timer[12]),
    .b(timer[13]),
    .c(timer[16]),
    .d(timer[17]),
    .o(_al_u1643_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*C*~B*A)"),
    .INIT(32'h00000020))
    _al_u1644 (
    .a(_al_u1643_o),
    .b(timer[24]),
    .c(timer[25]),
    .d(timer[26]),
    .e(timer[27]),
    .o(_al_u1644_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u1645 (
    .a(timer[14]),
    .b(timer[15]),
    .c(timer[18]),
    .d(timer[19]),
    .o(_al_u1645_o));
  AL_MAP_LUT4 #(
    .EQN("~(D*C*B*A)"),
    .INIT(16'h7fff))
    _al_u1646 (
    .a(_al_u1640_o),
    .b(_al_u1642_o),
    .c(_al_u1644_o),
    .d(_al_u1645_o),
    .o(n4_neg));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    _al_u1647 (
    .a(_al_u1638_o),
    .b(timer[10]),
    .c(timer[11]),
    .d(timer[8]),
    .o(_al_u1647_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    _al_u1648 (
    .a(_al_u1641_o),
    .b(timer[4]),
    .c(timer[5]),
    .d(timer[6]),
    .e(timer[7]),
    .o(_al_u1648_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u1649 (
    .a(timer[22]),
    .b(timer[23]),
    .c(timer[26]),
    .d(timer[27]),
    .o(_al_u1649_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*~C*~B*A)"),
    .INIT(32'h02000000))
    _al_u1650 (
    .a(_al_u1649_o),
    .b(timer[12]),
    .c(timer[13]),
    .d(timer[16]),
    .e(timer[17]),
    .o(_al_u1650_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*~B*A)"),
    .INIT(32'h20000000))
    _al_u1651 (
    .a(_al_u1645_o),
    .b(timer[20]),
    .c(timer[21]),
    .d(timer[24]),
    .e(timer[25]),
    .o(_al_u1651_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1652 (
    .a(_al_u1647_o),
    .b(_al_u1648_o),
    .c(_al_u1650_o),
    .d(_al_u1651_o),
    .o(_al_u1652_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1653 (
    .a(_al_u1652_o),
    .b(n2[9]),
    .o(n3[9]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1654 (
    .a(_al_u1652_o),
    .b(n2[8]),
    .o(n3[8]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1655 (
    .a(_al_u1652_o),
    .b(n2[7]),
    .o(n3[7]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1656 (
    .a(_al_u1652_o),
    .b(n2[6]),
    .o(n3[6]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1657 (
    .a(_al_u1652_o),
    .b(n2[5]),
    .o(n3[5]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1658 (
    .a(_al_u1652_o),
    .b(n2[4]),
    .o(n3[4]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1659 (
    .a(_al_u1652_o),
    .b(n2[31]),
    .o(n3[31]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1660 (
    .a(_al_u1652_o),
    .b(n2[30]),
    .o(n3[30]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1661 (
    .a(_al_u1652_o),
    .b(n2[3]),
    .o(n3[3]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1662 (
    .a(_al_u1652_o),
    .b(n2[29]),
    .o(n3[29]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1663 (
    .a(_al_u1652_o),
    .b(n2[28]),
    .o(n3[28]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1664 (
    .a(_al_u1652_o),
    .b(n2[27]),
    .o(n3[27]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1665 (
    .a(_al_u1652_o),
    .b(n2[26]),
    .o(n3[26]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1666 (
    .a(_al_u1652_o),
    .b(n2[25]),
    .o(n3[25]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1667 (
    .a(_al_u1652_o),
    .b(n2[24]),
    .o(n3[24]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1668 (
    .a(_al_u1652_o),
    .b(n2[23]),
    .o(n3[23]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1669 (
    .a(_al_u1652_o),
    .b(n2[22]),
    .o(n3[22]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1670 (
    .a(_al_u1652_o),
    .b(n2[21]),
    .o(n3[21]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1671 (
    .a(_al_u1652_o),
    .b(n2[20]),
    .o(n3[20]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1672 (
    .a(_al_u1652_o),
    .b(n2[2]),
    .o(n3[2]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1673 (
    .a(_al_u1652_o),
    .b(n2[19]),
    .o(n3[19]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1674 (
    .a(_al_u1652_o),
    .b(n2[18]),
    .o(n3[18]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1675 (
    .a(_al_u1652_o),
    .b(n2[17]),
    .o(n3[17]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1676 (
    .a(_al_u1652_o),
    .b(n2[16]),
    .o(n3[16]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1677 (
    .a(_al_u1652_o),
    .b(n2[15]),
    .o(n3[15]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1678 (
    .a(_al_u1652_o),
    .b(n2[14]),
    .o(n3[14]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1679 (
    .a(_al_u1652_o),
    .b(n2[13]),
    .o(n3[13]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1680 (
    .a(_al_u1652_o),
    .b(n2[12]),
    .o(n3[12]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1681 (
    .a(_al_u1652_o),
    .b(n2[11]),
    .o(n3[11]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1682 (
    .a(_al_u1652_o),
    .b(n2[10]),
    .o(n3[10]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1683 (
    .a(_al_u1652_o),
    .b(n2[1]),
    .o(n3[1]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1684 (
    .a(_al_u1652_o),
    .b(n2[0]),
    .o(n3[0]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1685 (
    .a(\PWM0/n0_lutinv ),
    .b(pwm_state_read[0]),
    .o(\PWM0/n24 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1686 (
    .a(pnumcnt0[18]),
    .b(pnumcnt0[19]),
    .c(pnumcnt0[1]),
    .d(pnumcnt0[20]),
    .o(_al_u1686_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u1687 (
    .a(_al_u1686_o),
    .b(pnumcnt0[21]),
    .c(pnumcnt0[22]),
    .d(pnumcnt0[23]),
    .e(pnumcnt0[2]),
    .o(_al_u1687_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u1688 (
    .a(_al_u1687_o),
    .b(pnumcnt0[6]),
    .c(pnumcnt0[7]),
    .d(pnumcnt0[8]),
    .e(pnumcnt0[9]),
    .o(_al_u1688_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1689 (
    .a(pnumcnt0[10]),
    .b(pnumcnt0[11]),
    .c(pnumcnt0[12]),
    .d(pnumcnt0[13]),
    .o(_al_u1689_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u1690 (
    .a(_al_u1689_o),
    .b(pnumcnt0[14]),
    .c(pnumcnt0[15]),
    .d(pnumcnt0[16]),
    .e(pnumcnt0[17]),
    .o(_al_u1690_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u1691 (
    .a(pnumcnt0[3]),
    .b(pnumcnt0[4]),
    .c(pnumcnt0[5]),
    .o(_al_u1691_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u1692 (
    .a(_al_u1688_o),
    .b(_al_u1690_o),
    .c(_al_u1691_o),
    .d(pnumcnt0[0]),
    .o(\PWM0/n25_neg_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1693 (
    .a(\PWM0/n24 ),
    .b(\PWM0/n25_neg_lutinv ),
    .c(\PWM0/n26 [9]),
    .d(\PWM0/pnumr [9]),
    .o(_al_u1693_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1694 (
    .a(_al_u1693_o),
    .b(\PWM0/n24 ),
    .c(pnumcnt0[9]),
    .d(\PWM0/pnumr [9]),
    .e(pwm_start_stop[16]),
    .o(\PWM0/n31 [9]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1695 (
    .a(\PWM0/n24 ),
    .b(\PWM0/n25_neg_lutinv ),
    .c(\PWM0/n26 [8]),
    .d(\PWM0/pnumr [8]),
    .o(_al_u1695_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1696 (
    .a(_al_u1695_o),
    .b(\PWM0/n24 ),
    .c(pnumcnt0[8]),
    .d(\PWM0/pnumr [8]),
    .e(pwm_start_stop[16]),
    .o(\PWM0/n31 [8]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1697 (
    .a(\PWM0/n24 ),
    .b(\PWM0/n25_neg_lutinv ),
    .c(\PWM0/n26 [7]),
    .d(\PWM0/pnumr [7]),
    .o(_al_u1697_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1698 (
    .a(_al_u1697_o),
    .b(\PWM0/n24 ),
    .c(pnumcnt0[7]),
    .d(\PWM0/pnumr [7]),
    .e(pwm_start_stop[16]),
    .o(\PWM0/n31 [7]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1699 (
    .a(\PWM0/n24 ),
    .b(\PWM0/n25_neg_lutinv ),
    .c(\PWM0/n26 [6]),
    .d(\PWM0/pnumr [6]),
    .o(_al_u1699_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1700 (
    .a(_al_u1699_o),
    .b(\PWM0/n24 ),
    .c(pnumcnt0[6]),
    .d(\PWM0/pnumr [6]),
    .e(pwm_start_stop[16]),
    .o(\PWM0/n31 [6]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1701 (
    .a(\PWM0/n24 ),
    .b(\PWM0/n25_neg_lutinv ),
    .c(\PWM0/n26 [5]),
    .d(\PWM0/pnumr [5]),
    .o(_al_u1701_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1702 (
    .a(_al_u1701_o),
    .b(\PWM0/n24 ),
    .c(pnumcnt0[5]),
    .d(\PWM0/pnumr [5]),
    .e(pwm_start_stop[16]),
    .o(\PWM0/n31 [5]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1703 (
    .a(\PWM0/n24 ),
    .b(\PWM0/n25_neg_lutinv ),
    .c(\PWM0/n26 [4]),
    .d(\PWM0/pnumr [4]),
    .o(_al_u1703_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1704 (
    .a(_al_u1703_o),
    .b(\PWM0/n24 ),
    .c(pnumcnt0[4]),
    .d(\PWM0/pnumr [4]),
    .e(pwm_start_stop[16]),
    .o(\PWM0/n31 [4]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1705 (
    .a(\PWM0/n24 ),
    .b(\PWM0/n25_neg_lutinv ),
    .c(\PWM0/n26 [3]),
    .d(\PWM0/pnumr [3]),
    .o(_al_u1705_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1706 (
    .a(_al_u1705_o),
    .b(\PWM0/n24 ),
    .c(pnumcnt0[3]),
    .d(\PWM0/pnumr [3]),
    .e(pwm_start_stop[16]),
    .o(\PWM0/n31 [3]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1707 (
    .a(\PWM0/n24 ),
    .b(\PWM0/n25_neg_lutinv ),
    .c(\PWM0/n26 [23]),
    .d(\PWM0/pnumr [23]),
    .o(_al_u1707_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1708 (
    .a(_al_u1707_o),
    .b(\PWM0/n24 ),
    .c(pnumcnt0[23]),
    .d(\PWM0/pnumr [23]),
    .e(pwm_start_stop[16]),
    .o(\PWM0/n31 [23]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1709 (
    .a(\PWM0/n24 ),
    .b(\PWM0/n25_neg_lutinv ),
    .c(\PWM0/n26 [22]),
    .d(\PWM0/pnumr [22]),
    .o(_al_u1709_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1710 (
    .a(_al_u1709_o),
    .b(\PWM0/n24 ),
    .c(pnumcnt0[22]),
    .d(\PWM0/pnumr [22]),
    .e(pwm_start_stop[16]),
    .o(\PWM0/n31 [22]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1711 (
    .a(\PWM0/n24 ),
    .b(\PWM0/n25_neg_lutinv ),
    .c(\PWM0/n26 [21]),
    .d(\PWM0/pnumr [21]),
    .o(_al_u1711_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1712 (
    .a(_al_u1711_o),
    .b(\PWM0/n24 ),
    .c(pnumcnt0[21]),
    .d(\PWM0/pnumr [21]),
    .e(pwm_start_stop[16]),
    .o(\PWM0/n31 [21]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1713 (
    .a(\PWM0/n24 ),
    .b(\PWM0/n25_neg_lutinv ),
    .c(\PWM0/n26 [20]),
    .d(\PWM0/pnumr [20]),
    .o(_al_u1713_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1714 (
    .a(_al_u1713_o),
    .b(\PWM0/n24 ),
    .c(pnumcnt0[20]),
    .d(\PWM0/pnumr [20]),
    .e(pwm_start_stop[16]),
    .o(\PWM0/n31 [20]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1715 (
    .a(\PWM0/n24 ),
    .b(\PWM0/n25_neg_lutinv ),
    .c(\PWM0/n26 [2]),
    .d(\PWM0/pnumr [2]),
    .o(_al_u1715_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1716 (
    .a(_al_u1715_o),
    .b(\PWM0/n24 ),
    .c(pnumcnt0[2]),
    .d(\PWM0/pnumr [2]),
    .e(pwm_start_stop[16]),
    .o(\PWM0/n31 [2]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1717 (
    .a(\PWM0/n24 ),
    .b(\PWM0/n25_neg_lutinv ),
    .c(\PWM0/n26 [19]),
    .d(\PWM0/pnumr [19]),
    .o(_al_u1717_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1718 (
    .a(_al_u1717_o),
    .b(\PWM0/n24 ),
    .c(pnumcnt0[19]),
    .d(\PWM0/pnumr [19]),
    .e(pwm_start_stop[16]),
    .o(\PWM0/n31 [19]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1719 (
    .a(\PWM0/n24 ),
    .b(\PWM0/n25_neg_lutinv ),
    .c(\PWM0/n26 [18]),
    .d(\PWM0/pnumr [18]),
    .o(_al_u1719_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1720 (
    .a(_al_u1719_o),
    .b(\PWM0/n24 ),
    .c(pnumcnt0[18]),
    .d(\PWM0/pnumr [18]),
    .e(pwm_start_stop[16]),
    .o(\PWM0/n31 [18]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1721 (
    .a(\PWM0/n24 ),
    .b(\PWM0/n25_neg_lutinv ),
    .c(\PWM0/n26 [17]),
    .d(\PWM0/pnumr [17]),
    .o(_al_u1721_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1722 (
    .a(_al_u1721_o),
    .b(\PWM0/n24 ),
    .c(pnumcnt0[17]),
    .d(\PWM0/pnumr [17]),
    .e(pwm_start_stop[16]),
    .o(\PWM0/n31 [17]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1723 (
    .a(\PWM0/n24 ),
    .b(\PWM0/n25_neg_lutinv ),
    .c(\PWM0/n26 [16]),
    .d(\PWM0/pnumr [16]),
    .o(_al_u1723_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1724 (
    .a(_al_u1723_o),
    .b(\PWM0/n24 ),
    .c(pnumcnt0[16]),
    .d(\PWM0/pnumr [16]),
    .e(pwm_start_stop[16]),
    .o(\PWM0/n31 [16]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1725 (
    .a(\PWM0/n24 ),
    .b(\PWM0/n25_neg_lutinv ),
    .c(\PWM0/n26 [15]),
    .d(\PWM0/pnumr [15]),
    .o(_al_u1725_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1726 (
    .a(_al_u1725_o),
    .b(\PWM0/n24 ),
    .c(pnumcnt0[15]),
    .d(\PWM0/pnumr [15]),
    .e(pwm_start_stop[16]),
    .o(\PWM0/n31 [15]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1727 (
    .a(\PWM0/n24 ),
    .b(\PWM0/n25_neg_lutinv ),
    .c(\PWM0/n26 [14]),
    .d(\PWM0/pnumr [14]),
    .o(_al_u1727_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1728 (
    .a(_al_u1727_o),
    .b(\PWM0/n24 ),
    .c(pnumcnt0[14]),
    .d(\PWM0/pnumr [14]),
    .e(pwm_start_stop[16]),
    .o(\PWM0/n31 [14]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1729 (
    .a(\PWM0/n24 ),
    .b(\PWM0/n25_neg_lutinv ),
    .c(\PWM0/n26 [13]),
    .d(\PWM0/pnumr [13]),
    .o(_al_u1729_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u173 (
    .a(pwm_state_read[0]),
    .b(pwm_start_stop[16]),
    .o(\PWM0/n11 ));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1730 (
    .a(_al_u1729_o),
    .b(\PWM0/n24 ),
    .c(pnumcnt0[13]),
    .d(\PWM0/pnumr [13]),
    .e(pwm_start_stop[16]),
    .o(\PWM0/n31 [13]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1731 (
    .a(\PWM0/n24 ),
    .b(\PWM0/n25_neg_lutinv ),
    .c(\PWM0/n26 [12]),
    .d(\PWM0/pnumr [12]),
    .o(_al_u1731_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1732 (
    .a(_al_u1731_o),
    .b(\PWM0/n24 ),
    .c(pnumcnt0[12]),
    .d(\PWM0/pnumr [12]),
    .e(pwm_start_stop[16]),
    .o(\PWM0/n31 [12]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1733 (
    .a(\PWM0/n24 ),
    .b(\PWM0/n25_neg_lutinv ),
    .c(\PWM0/n26 [11]),
    .d(\PWM0/pnumr [11]),
    .o(_al_u1733_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1734 (
    .a(_al_u1733_o),
    .b(\PWM0/n24 ),
    .c(pnumcnt0[11]),
    .d(\PWM0/pnumr [11]),
    .e(pwm_start_stop[16]),
    .o(\PWM0/n31 [11]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1735 (
    .a(\PWM0/n24 ),
    .b(\PWM0/n25_neg_lutinv ),
    .c(\PWM0/n26 [10]),
    .d(\PWM0/pnumr [10]),
    .o(_al_u1735_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1736 (
    .a(_al_u1735_o),
    .b(\PWM0/n24 ),
    .c(pnumcnt0[10]),
    .d(\PWM0/pnumr [10]),
    .e(pwm_start_stop[16]),
    .o(\PWM0/n31 [10]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1737 (
    .a(\PWM0/n24 ),
    .b(\PWM0/n25_neg_lutinv ),
    .c(\PWM0/n26 [1]),
    .d(\PWM0/pnumr [1]),
    .o(_al_u1737_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1738 (
    .a(_al_u1737_o),
    .b(\PWM0/n24 ),
    .c(pnumcnt0[1]),
    .d(\PWM0/pnumr [1]),
    .e(pwm_start_stop[16]),
    .o(\PWM0/n31 [1]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1739 (
    .a(\PWM0/n24 ),
    .b(\PWM0/n25_neg_lutinv ),
    .c(\PWM0/n26 [0]),
    .d(\PWM0/pnumr [0]),
    .o(_al_u1739_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u174 (
    .a(pwm_state_read[1]),
    .b(pwm_start_stop[17]),
    .o(\PWM1/n11 ));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1740 (
    .a(_al_u1739_o),
    .b(\PWM0/n24 ),
    .c(pnumcnt0[0]),
    .d(\PWM0/pnumr [0]),
    .e(pwm_start_stop[16]),
    .o(\PWM0/n31 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u1741 (
    .a(\PWM0/FreCnt [0]),
    .b(\PWM0/FreCnt [8]),
    .c(\PWM0/FreCntr [1]),
    .d(\PWM0/FreCntr [9]),
    .o(_al_u1741_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*~C)*~(D*~B))"),
    .INIT(32'h80a088aa))
    _al_u1742 (
    .a(_al_u1741_o),
    .b(\PWM0/FreCnt [12]),
    .c(\PWM0/FreCnt [5]),
    .d(\PWM0/FreCntr [13]),
    .e(\PWM0/FreCntr [6]),
    .o(_al_u1742_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u1743 (
    .a(\PWM0/FreCnt [12]),
    .b(\PWM0/FreCnt [8]),
    .c(\PWM0/FreCntr [13]),
    .d(\PWM0/FreCntr [9]),
    .o(_al_u1743_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D@C))"),
    .INIT(16'h8008))
    _al_u1744 (
    .a(_al_u1742_o),
    .b(_al_u1743_o),
    .c(\PWM0/FreCnt [9]),
    .d(\PWM0/FreCntr [10]),
    .o(_al_u1744_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u1745 (
    .a(\PWM0/FreCnt [19]),
    .b(\PWM0/FreCnt [3]),
    .c(\PWM0/FreCntr [20]),
    .d(\PWM0/FreCntr [4]),
    .o(_al_u1745_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*~C)*~(D*~B))"),
    .INIT(32'h80a088aa))
    _al_u1746 (
    .a(_al_u1745_o),
    .b(\PWM0/FreCnt [13]),
    .c(\PWM0/FreCnt [25]),
    .d(\PWM0/FreCntr [14]),
    .e(\PWM0/FreCntr [26]),
    .o(_al_u1746_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u1747 (
    .a(\PWM0/FreCnt [15]),
    .b(\PWM0/FreCnt [7]),
    .c(\PWM0/FreCntr [16]),
    .d(\PWM0/FreCntr [8]),
    .o(_al_u1747_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u1748 (
    .a(_al_u1744_o),
    .b(_al_u1746_o),
    .c(_al_u1747_o),
    .d(\PWM0/FreCnt [6]),
    .e(\PWM0/FreCntr [7]),
    .o(_al_u1748_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1749 (
    .a(\PWM0/FreCnt [14]),
    .b(\PWM0/FreCnt [4]),
    .c(\PWM0/FreCntr [15]),
    .d(\PWM0/FreCntr [5]),
    .o(_al_u1749_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u175 (
    .a(pwm_state_read[2]),
    .b(pwm_start_stop[18]),
    .o(\PWM2/n11 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u1750 (
    .a(_al_u1749_o),
    .b(\PWM0/FreCnt [21]),
    .c(\PWM0/FreCntr [22]),
    .o(_al_u1750_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1751 (
    .a(\PWM0/FreCnt [18]),
    .b(\PWM0/FreCnt [2]),
    .c(\PWM0/FreCntr [19]),
    .d(\PWM0/FreCntr [3]),
    .o(_al_u1751_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1752 (
    .a(_al_u1751_o),
    .b(\PWM0/FreCnt [20]),
    .c(\PWM0/FreCnt [22]),
    .d(\PWM0/FreCntr [21]),
    .e(\PWM0/FreCntr [23]),
    .o(_al_u1752_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1753 (
    .a(\PWM0/FreCnt [13]),
    .b(\PWM0/FreCntr [14]),
    .o(_al_u1753_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(E*~C)*~(D@B))"),
    .INIT(32'h40104411))
    _al_u1754 (
    .a(_al_u1753_o),
    .b(\PWM0/FreCnt [10]),
    .c(\PWM0/FreCnt [16]),
    .d(\PWM0/FreCntr [11]),
    .e(\PWM0/FreCntr [17]),
    .o(_al_u1754_o));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(~E*B)*~(D@A))"),
    .INIT(32'h0a050201))
    _al_u1755 (
    .a(\PWM0/FreCnt [11]),
    .b(\PWM0/FreCnt [16]),
    .c(\PWM0/FreCnt [26]),
    .d(\PWM0/FreCntr [12]),
    .e(\PWM0/FreCntr [17]),
    .o(_al_u1755_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1756 (
    .a(_al_u1750_o),
    .b(_al_u1752_o),
    .c(_al_u1754_o),
    .d(_al_u1755_o),
    .o(_al_u1756_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u1757 (
    .a(\PWM0/FreCnt [1]),
    .b(\PWM0/FreCnt [25]),
    .c(\PWM0/FreCntr [2]),
    .d(\PWM0/FreCntr [26]),
    .o(_al_u1757_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*~C)*~(D*~B))"),
    .INIT(32'h80a088aa))
    _al_u1758 (
    .a(_al_u1757_o),
    .b(\PWM0/FreCnt [17]),
    .c(\PWM0/FreCnt [19]),
    .d(\PWM0/FreCntr [18]),
    .e(\PWM0/FreCntr [20]),
    .o(_al_u1758_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u1759 (
    .a(\PWM0/FreCnt [5]),
    .b(\PWM0/FreCnt [7]),
    .c(\PWM0/FreCntr [6]),
    .d(\PWM0/FreCntr [8]),
    .o(_al_u1759_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u176 (
    .a(pwm_state_read[3]),
    .b(pwm_start_stop[19]),
    .o(\PWM3/n11 ));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*~C))"),
    .INIT(16'h8088))
    _al_u1760 (
    .a(_al_u1758_o),
    .b(_al_u1759_o),
    .c(\PWM0/FreCnt [23]),
    .d(\PWM0/FreCntr [24]),
    .o(_al_u1760_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u1761 (
    .a(\PWM0/FreCnt [1]),
    .b(\PWM0/FreCnt [23]),
    .c(\PWM0/FreCntr [2]),
    .d(\PWM0/FreCntr [24]),
    .o(_al_u1761_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*C)*~(~D*B))"),
    .INIT(32'haa220a02))
    _al_u1762 (
    .a(_al_u1761_o),
    .b(\PWM0/FreCnt [15]),
    .c(\PWM0/FreCnt [17]),
    .d(\PWM0/FreCntr [16]),
    .e(\PWM0/FreCntr [18]),
    .o(_al_u1762_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1763 (
    .a(\PWM0/FreCnt [3]),
    .b(\PWM0/FreCntr [4]),
    .o(_al_u1763_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(E@C)*~(D*~B))"),
    .INIT(32'h40500405))
    _al_u1764 (
    .a(_al_u1763_o),
    .b(\PWM0/FreCnt [0]),
    .c(\PWM0/FreCnt [24]),
    .d(\PWM0/FreCntr [1]),
    .e(\PWM0/FreCntr [25]),
    .o(_al_u1764_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    _al_u1765 (
    .a(_al_u1748_o),
    .b(_al_u1756_o),
    .c(_al_u1760_o),
    .d(_al_u1762_o),
    .e(_al_u1764_o),
    .o(_al_u1765_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1766 (
    .a(_al_u1765_o),
    .b(pwm_state_read[0]),
    .o(\PWM0/u14_sel_is_1_o ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1767 (
    .a(\PWM1/n0_lutinv ),
    .b(pwm_state_read[1]),
    .o(\PWM1/n24 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1768 (
    .a(pnumcnt1[18]),
    .b(pnumcnt1[19]),
    .c(pnumcnt1[1]),
    .d(pnumcnt1[20]),
    .o(_al_u1768_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u1769 (
    .a(_al_u1768_o),
    .b(pnumcnt1[21]),
    .c(pnumcnt1[22]),
    .d(pnumcnt1[23]),
    .e(pnumcnt1[2]),
    .o(_al_u1769_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u177 (
    .a(pwm_state_read[4]),
    .b(pwm_start_stop[20]),
    .o(\PWM4/n11 ));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u1770 (
    .a(_al_u1769_o),
    .b(pnumcnt1[6]),
    .c(pnumcnt1[7]),
    .d(pnumcnt1[8]),
    .e(pnumcnt1[9]),
    .o(_al_u1770_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1771 (
    .a(pnumcnt1[10]),
    .b(pnumcnt1[11]),
    .c(pnumcnt1[12]),
    .d(pnumcnt1[13]),
    .o(_al_u1771_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u1772 (
    .a(_al_u1771_o),
    .b(pnumcnt1[14]),
    .c(pnumcnt1[15]),
    .d(pnumcnt1[16]),
    .e(pnumcnt1[17]),
    .o(_al_u1772_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u1773 (
    .a(pnumcnt1[3]),
    .b(pnumcnt1[4]),
    .c(pnumcnt1[5]),
    .o(_al_u1773_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u1774 (
    .a(_al_u1770_o),
    .b(_al_u1772_o),
    .c(_al_u1773_o),
    .d(pnumcnt1[0]),
    .o(\PWM1/n25_neg_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1775 (
    .a(\PWM1/n24 ),
    .b(\PWM1/n25_neg_lutinv ),
    .c(\PWM1/n26 [9]),
    .d(\PWM1/pnumr [9]),
    .o(_al_u1775_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1776 (
    .a(_al_u1775_o),
    .b(\PWM1/n24 ),
    .c(pnumcnt1[9]),
    .d(\PWM1/pnumr [9]),
    .e(pwm_start_stop[17]),
    .o(\PWM1/n31 [9]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1777 (
    .a(\PWM1/n24 ),
    .b(\PWM1/n25_neg_lutinv ),
    .c(\PWM1/n26 [8]),
    .d(\PWM1/pnumr [8]),
    .o(_al_u1777_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1778 (
    .a(_al_u1777_o),
    .b(\PWM1/n24 ),
    .c(pnumcnt1[8]),
    .d(\PWM1/pnumr [8]),
    .e(pwm_start_stop[17]),
    .o(\PWM1/n31 [8]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1779 (
    .a(\PWM1/n24 ),
    .b(\PWM1/n25_neg_lutinv ),
    .c(\PWM1/n26 [7]),
    .d(\PWM1/pnumr [7]),
    .o(_al_u1779_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u178 (
    .a(pwm_state_read[5]),
    .b(pwm_start_stop[21]),
    .o(\PWM5/n11 ));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1780 (
    .a(_al_u1779_o),
    .b(\PWM1/n24 ),
    .c(pnumcnt1[7]),
    .d(\PWM1/pnumr [7]),
    .e(pwm_start_stop[17]),
    .o(\PWM1/n31 [7]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1781 (
    .a(\PWM1/n24 ),
    .b(\PWM1/n25_neg_lutinv ),
    .c(\PWM1/n26 [6]),
    .d(\PWM1/pnumr [6]),
    .o(_al_u1781_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1782 (
    .a(_al_u1781_o),
    .b(\PWM1/n24 ),
    .c(pnumcnt1[6]),
    .d(\PWM1/pnumr [6]),
    .e(pwm_start_stop[17]),
    .o(\PWM1/n31 [6]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1783 (
    .a(\PWM1/n24 ),
    .b(\PWM1/n25_neg_lutinv ),
    .c(\PWM1/n26 [5]),
    .d(\PWM1/pnumr [5]),
    .o(_al_u1783_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1784 (
    .a(_al_u1783_o),
    .b(\PWM1/n24 ),
    .c(pnumcnt1[5]),
    .d(\PWM1/pnumr [5]),
    .e(pwm_start_stop[17]),
    .o(\PWM1/n31 [5]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1785 (
    .a(\PWM1/n24 ),
    .b(\PWM1/n25_neg_lutinv ),
    .c(\PWM1/n26 [4]),
    .d(\PWM1/pnumr [4]),
    .o(_al_u1785_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1786 (
    .a(_al_u1785_o),
    .b(\PWM1/n24 ),
    .c(pnumcnt1[4]),
    .d(\PWM1/pnumr [4]),
    .e(pwm_start_stop[17]),
    .o(\PWM1/n31 [4]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1787 (
    .a(\PWM1/n24 ),
    .b(\PWM1/n25_neg_lutinv ),
    .c(\PWM1/n26 [3]),
    .d(\PWM1/pnumr [3]),
    .o(_al_u1787_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1788 (
    .a(_al_u1787_o),
    .b(\PWM1/n24 ),
    .c(pnumcnt1[3]),
    .d(\PWM1/pnumr [3]),
    .e(pwm_start_stop[17]),
    .o(\PWM1/n31 [3]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1789 (
    .a(\PWM1/n24 ),
    .b(\PWM1/n25_neg_lutinv ),
    .c(\PWM1/n26 [23]),
    .d(\PWM1/pnumr [23]),
    .o(_al_u1789_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u179 (
    .a(pwm_state_read[6]),
    .b(pwm_start_stop[22]),
    .o(\PWM6/n11 ));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1790 (
    .a(_al_u1789_o),
    .b(\PWM1/n24 ),
    .c(pnumcnt1[23]),
    .d(\PWM1/pnumr [23]),
    .e(pwm_start_stop[17]),
    .o(\PWM1/n31 [23]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1791 (
    .a(\PWM1/n24 ),
    .b(\PWM1/n25_neg_lutinv ),
    .c(\PWM1/n26 [22]),
    .d(\PWM1/pnumr [22]),
    .o(_al_u1791_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1792 (
    .a(_al_u1791_o),
    .b(\PWM1/n24 ),
    .c(pnumcnt1[22]),
    .d(\PWM1/pnumr [22]),
    .e(pwm_start_stop[17]),
    .o(\PWM1/n31 [22]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1793 (
    .a(\PWM1/n24 ),
    .b(\PWM1/n25_neg_lutinv ),
    .c(\PWM1/n26 [21]),
    .d(\PWM1/pnumr [21]),
    .o(_al_u1793_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1794 (
    .a(_al_u1793_o),
    .b(\PWM1/n24 ),
    .c(pnumcnt1[21]),
    .d(\PWM1/pnumr [21]),
    .e(pwm_start_stop[17]),
    .o(\PWM1/n31 [21]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1795 (
    .a(\PWM1/n24 ),
    .b(\PWM1/n25_neg_lutinv ),
    .c(\PWM1/n26 [20]),
    .d(\PWM1/pnumr [20]),
    .o(_al_u1795_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1796 (
    .a(_al_u1795_o),
    .b(\PWM1/n24 ),
    .c(pnumcnt1[20]),
    .d(\PWM1/pnumr [20]),
    .e(pwm_start_stop[17]),
    .o(\PWM1/n31 [20]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1797 (
    .a(\PWM1/n24 ),
    .b(\PWM1/n25_neg_lutinv ),
    .c(\PWM1/n26 [2]),
    .d(\PWM1/pnumr [2]),
    .o(_al_u1797_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1798 (
    .a(_al_u1797_o),
    .b(\PWM1/n24 ),
    .c(pnumcnt1[2]),
    .d(\PWM1/pnumr [2]),
    .e(pwm_start_stop[17]),
    .o(\PWM1/n31 [2]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1799 (
    .a(\PWM1/n24 ),
    .b(\PWM1/n25_neg_lutinv ),
    .c(\PWM1/n26 [19]),
    .d(\PWM1/pnumr [19]),
    .o(_al_u1799_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u180 (
    .a(pwm_state_read[7]),
    .b(pwm_start_stop[23]),
    .o(\PWM7/n11 ));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1800 (
    .a(_al_u1799_o),
    .b(\PWM1/n24 ),
    .c(pnumcnt1[19]),
    .d(\PWM1/pnumr [19]),
    .e(pwm_start_stop[17]),
    .o(\PWM1/n31 [19]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1801 (
    .a(\PWM1/n24 ),
    .b(\PWM1/n25_neg_lutinv ),
    .c(\PWM1/n26 [18]),
    .d(\PWM1/pnumr [18]),
    .o(_al_u1801_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1802 (
    .a(_al_u1801_o),
    .b(\PWM1/n24 ),
    .c(pnumcnt1[18]),
    .d(\PWM1/pnumr [18]),
    .e(pwm_start_stop[17]),
    .o(\PWM1/n31 [18]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1803 (
    .a(\PWM1/n24 ),
    .b(\PWM1/n25_neg_lutinv ),
    .c(\PWM1/n26 [17]),
    .d(\PWM1/pnumr [17]),
    .o(_al_u1803_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1804 (
    .a(_al_u1803_o),
    .b(\PWM1/n24 ),
    .c(pnumcnt1[17]),
    .d(\PWM1/pnumr [17]),
    .e(pwm_start_stop[17]),
    .o(\PWM1/n31 [17]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1805 (
    .a(\PWM1/n24 ),
    .b(\PWM1/n25_neg_lutinv ),
    .c(\PWM1/n26 [16]),
    .d(\PWM1/pnumr [16]),
    .o(_al_u1805_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1806 (
    .a(_al_u1805_o),
    .b(\PWM1/n24 ),
    .c(pnumcnt1[16]),
    .d(\PWM1/pnumr [16]),
    .e(pwm_start_stop[17]),
    .o(\PWM1/n31 [16]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1807 (
    .a(\PWM1/n24 ),
    .b(\PWM1/n25_neg_lutinv ),
    .c(\PWM1/n26 [15]),
    .d(\PWM1/pnumr [15]),
    .o(_al_u1807_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1808 (
    .a(_al_u1807_o),
    .b(\PWM1/n24 ),
    .c(pnumcnt1[15]),
    .d(\PWM1/pnumr [15]),
    .e(pwm_start_stop[17]),
    .o(\PWM1/n31 [15]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1809 (
    .a(\PWM1/n24 ),
    .b(\PWM1/n25_neg_lutinv ),
    .c(\PWM1/n26 [14]),
    .d(\PWM1/pnumr [14]),
    .o(_al_u1809_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u181 (
    .a(pwm_state_read[8]),
    .b(pwm_start_stop[24]),
    .o(\PWM8/n11 ));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1810 (
    .a(_al_u1809_o),
    .b(\PWM1/n24 ),
    .c(pnumcnt1[14]),
    .d(\PWM1/pnumr [14]),
    .e(pwm_start_stop[17]),
    .o(\PWM1/n31 [14]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1811 (
    .a(\PWM1/n24 ),
    .b(\PWM1/n25_neg_lutinv ),
    .c(\PWM1/n26 [13]),
    .d(\PWM1/pnumr [13]),
    .o(_al_u1811_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1812 (
    .a(_al_u1811_o),
    .b(\PWM1/n24 ),
    .c(pnumcnt1[13]),
    .d(\PWM1/pnumr [13]),
    .e(pwm_start_stop[17]),
    .o(\PWM1/n31 [13]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1813 (
    .a(\PWM1/n24 ),
    .b(\PWM1/n25_neg_lutinv ),
    .c(\PWM1/n26 [12]),
    .d(\PWM1/pnumr [12]),
    .o(_al_u1813_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1814 (
    .a(_al_u1813_o),
    .b(\PWM1/n24 ),
    .c(pnumcnt1[12]),
    .d(\PWM1/pnumr [12]),
    .e(pwm_start_stop[17]),
    .o(\PWM1/n31 [12]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1815 (
    .a(\PWM1/n24 ),
    .b(\PWM1/n25_neg_lutinv ),
    .c(\PWM1/n26 [11]),
    .d(\PWM1/pnumr [11]),
    .o(_al_u1815_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1816 (
    .a(_al_u1815_o),
    .b(\PWM1/n24 ),
    .c(pnumcnt1[11]),
    .d(\PWM1/pnumr [11]),
    .e(pwm_start_stop[17]),
    .o(\PWM1/n31 [11]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1817 (
    .a(\PWM1/n24 ),
    .b(\PWM1/n25_neg_lutinv ),
    .c(\PWM1/n26 [10]),
    .d(\PWM1/pnumr [10]),
    .o(_al_u1817_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1818 (
    .a(_al_u1817_o),
    .b(\PWM1/n24 ),
    .c(pnumcnt1[10]),
    .d(\PWM1/pnumr [10]),
    .e(pwm_start_stop[17]),
    .o(\PWM1/n31 [10]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1819 (
    .a(\PWM1/n24 ),
    .b(\PWM1/n25_neg_lutinv ),
    .c(\PWM1/n26 [1]),
    .d(\PWM1/pnumr [1]),
    .o(_al_u1819_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u182 (
    .a(pwm_state_read[9]),
    .b(pwm_start_stop[25]),
    .o(\PWM9/n11 ));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1820 (
    .a(_al_u1819_o),
    .b(\PWM1/n24 ),
    .c(pnumcnt1[1]),
    .d(\PWM1/pnumr [1]),
    .e(pwm_start_stop[17]),
    .o(\PWM1/n31 [1]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1821 (
    .a(\PWM1/n24 ),
    .b(\PWM1/n25_neg_lutinv ),
    .c(\PWM1/n26 [0]),
    .d(\PWM1/pnumr [0]),
    .o(_al_u1821_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1822 (
    .a(_al_u1821_o),
    .b(\PWM1/n24 ),
    .c(pnumcnt1[0]),
    .d(\PWM1/pnumr [0]),
    .e(pwm_start_stop[17]),
    .o(\PWM1/n31 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u1823 (
    .a(\PWM1/FreCnt [10]),
    .b(\PWM1/FreCnt [17]),
    .c(\PWM1/FreCntr [11]),
    .d(\PWM1/FreCntr [18]),
    .o(_al_u1823_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*~C)*~(~D*B))"),
    .INIT(32'ha020aa22))
    _al_u1824 (
    .a(_al_u1823_o),
    .b(\PWM1/FreCnt [1]),
    .c(\PWM1/FreCnt [23]),
    .d(\PWM1/FreCntr [2]),
    .e(\PWM1/FreCntr [24]),
    .o(_al_u1824_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(~D*B))"),
    .INIT(32'ha0200a02))
    _al_u1825 (
    .a(_al_u1824_o),
    .b(\PWM1/FreCnt [12]),
    .c(\PWM1/FreCnt [14]),
    .d(\PWM1/FreCntr [13]),
    .e(\PWM1/FreCntr [15]),
    .o(_al_u1825_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u1826 (
    .a(\PWM1/FreCnt [12]),
    .b(\PWM1/FreCnt [21]),
    .c(\PWM1/FreCntr [13]),
    .d(\PWM1/FreCntr [22]),
    .o(_al_u1826_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u1827 (
    .a(_al_u1826_o),
    .b(\PWM1/FreCnt [16]),
    .c(\PWM1/FreCntr [17]),
    .o(_al_u1827_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u1828 (
    .a(\PWM1/FreCnt [13]),
    .b(\PWM1/FreCnt [17]),
    .c(\PWM1/FreCntr [14]),
    .d(\PWM1/FreCntr [18]),
    .o(_al_u1828_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u1829 (
    .a(_al_u1825_o),
    .b(_al_u1827_o),
    .c(_al_u1828_o),
    .d(\PWM1/FreCnt [9]),
    .e(\PWM1/FreCntr [10]),
    .o(_al_u1829_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u183 (
    .a(pwm_state_read[10]),
    .b(pwm_start_stop[26]),
    .o(\PWMA/n11 ));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u1830 (
    .a(\PWM1/FreCnt [13]),
    .b(\PWM1/FreCnt [7]),
    .c(\PWM1/FreCntr [14]),
    .d(\PWM1/FreCntr [8]),
    .o(_al_u1830_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*C)*~(D*~B))"),
    .INIT(32'h88aa080a))
    _al_u1831 (
    .a(_al_u1830_o),
    .b(\PWM1/FreCnt [18]),
    .c(\PWM1/FreCnt [23]),
    .d(\PWM1/FreCntr [19]),
    .e(\PWM1/FreCntr [24]),
    .o(_al_u1831_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1832 (
    .a(\PWM1/FreCnt [1]),
    .b(\PWM1/FreCntr [2]),
    .o(_al_u1832_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(~E*C)*~(D@B))"),
    .INIT(32'h44110401))
    _al_u1833 (
    .a(_al_u1832_o),
    .b(\PWM1/FreCnt [5]),
    .c(\PWM1/FreCnt [8]),
    .d(\PWM1/FreCntr [6]),
    .e(\PWM1/FreCntr [9]),
    .o(_al_u1833_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1834 (
    .a(\PWM1/FreCnt [10]),
    .b(\PWM1/FreCntr [11]),
    .o(_al_u1834_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(E*~C)*~(D@B))"),
    .INIT(32'h40104411))
    _al_u1835 (
    .a(_al_u1834_o),
    .b(\PWM1/FreCnt [22]),
    .c(\PWM1/FreCnt [3]),
    .d(\PWM1/FreCntr [23]),
    .e(\PWM1/FreCntr [4]),
    .o(_al_u1835_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1836 (
    .a(\PWM1/FreCnt [18]),
    .b(\PWM1/FreCntr [19]),
    .o(_al_u1836_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(E@C)*~(~D*B))"),
    .INIT(32'h50100501))
    _al_u1837 (
    .a(_al_u1836_o),
    .b(\PWM1/FreCnt [15]),
    .c(\PWM1/FreCnt [20]),
    .d(\PWM1/FreCntr [16]),
    .e(\PWM1/FreCntr [21]),
    .o(_al_u1837_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    _al_u1838 (
    .a(_al_u1829_o),
    .b(_al_u1831_o),
    .c(_al_u1833_o),
    .d(_al_u1835_o),
    .e(_al_u1837_o),
    .o(_al_u1838_o));
  AL_MAP_LUT5 #(
    .EQN("(~B*~(E@C)*~(D*~A))"),
    .INIT(32'h20300203))
    _al_u1839 (
    .a(\PWM1/FreCnt [19]),
    .b(\PWM1/FreCnt [26]),
    .c(\PWM1/FreCnt [4]),
    .d(\PWM1/FreCntr [20]),
    .e(\PWM1/FreCntr [5]),
    .o(_al_u1839_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u184 (
    .a(pwm_state_read[11]),
    .b(pwm_start_stop[27]),
    .o(\PWMB/n11 ));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1840 (
    .a(_al_u1839_o),
    .b(\PWM1/FreCnt [24]),
    .c(\PWM1/FreCnt [6]),
    .d(\PWM1/FreCntr [25]),
    .e(\PWM1/FreCntr [7]),
    .o(_al_u1840_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1841 (
    .a(\PWM1/FreCnt [0]),
    .b(\PWM1/FreCnt [11]),
    .c(\PWM1/FreCntr [1]),
    .d(\PWM1/FreCntr [12]),
    .o(_al_u1841_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u1842 (
    .a(_al_u1841_o),
    .b(\PWM1/FreCnt [2]),
    .c(\PWM1/FreCntr [3]),
    .o(_al_u1842_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u1843 (
    .a(\PWM1/FreCnt [15]),
    .b(\PWM1/FreCnt [19]),
    .c(\PWM1/FreCntr [16]),
    .d(\PWM1/FreCntr [20]),
    .o(_al_u1843_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*C)*~(D*~B))"),
    .INIT(32'h88aa080a))
    _al_u1844 (
    .a(_al_u1843_o),
    .b(\PWM1/FreCnt [25]),
    .c(\PWM1/FreCnt [3]),
    .d(\PWM1/FreCntr [26]),
    .e(\PWM1/FreCntr [4]),
    .o(_al_u1844_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u1845 (
    .a(\PWM1/FreCnt [7]),
    .b(\PWM1/FreCnt [8]),
    .c(\PWM1/FreCntr [8]),
    .d(\PWM1/FreCntr [9]),
    .o(_al_u1845_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*C)*~(~D*B))"),
    .INIT(32'haa220a02))
    _al_u1846 (
    .a(_al_u1845_o),
    .b(\PWM1/FreCnt [21]),
    .c(\PWM1/FreCnt [25]),
    .d(\PWM1/FreCntr [22]),
    .e(\PWM1/FreCntr [26]),
    .o(_al_u1846_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    _al_u1847 (
    .a(_al_u1838_o),
    .b(_al_u1840_o),
    .c(_al_u1842_o),
    .d(_al_u1844_o),
    .e(_al_u1846_o),
    .o(_al_u1847_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1848 (
    .a(_al_u1847_o),
    .b(pwm_state_read[1]),
    .o(\PWM1/u14_sel_is_1_o ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1849 (
    .a(\PWM2/n0_lutinv ),
    .b(pwm_state_read[2]),
    .o(\PWM2/n24 ));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u185 (
    .a(pwm_state_read[12]),
    .b(pwm_start_stop[28]),
    .o(\PWMC/n11 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1850 (
    .a(pnumcnt2[18]),
    .b(pnumcnt2[19]),
    .c(pnumcnt2[1]),
    .d(pnumcnt2[20]),
    .o(_al_u1850_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u1851 (
    .a(_al_u1850_o),
    .b(pnumcnt2[21]),
    .c(pnumcnt2[22]),
    .d(pnumcnt2[23]),
    .e(pnumcnt2[2]),
    .o(_al_u1851_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u1852 (
    .a(_al_u1851_o),
    .b(pnumcnt2[6]),
    .c(pnumcnt2[7]),
    .d(pnumcnt2[8]),
    .e(pnumcnt2[9]),
    .o(_al_u1852_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1853 (
    .a(pnumcnt2[10]),
    .b(pnumcnt2[11]),
    .c(pnumcnt2[12]),
    .d(pnumcnt2[13]),
    .o(_al_u1853_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u1854 (
    .a(_al_u1853_o),
    .b(pnumcnt2[14]),
    .c(pnumcnt2[15]),
    .d(pnumcnt2[16]),
    .e(pnumcnt2[17]),
    .o(_al_u1854_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u1855 (
    .a(pnumcnt2[3]),
    .b(pnumcnt2[4]),
    .c(pnumcnt2[5]),
    .o(_al_u1855_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u1856 (
    .a(_al_u1852_o),
    .b(_al_u1854_o),
    .c(_al_u1855_o),
    .d(pnumcnt2[0]),
    .o(\PWM2/n25_neg_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1857 (
    .a(\PWM2/n24 ),
    .b(\PWM2/n25_neg_lutinv ),
    .c(\PWM2/n26 [9]),
    .d(\PWM2/pnumr [9]),
    .o(_al_u1857_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1858 (
    .a(_al_u1857_o),
    .b(\PWM2/n24 ),
    .c(pnumcnt2[9]),
    .d(\PWM2/pnumr [9]),
    .e(pwm_start_stop[18]),
    .o(\PWM2/n31 [9]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1859 (
    .a(\PWM2/n24 ),
    .b(\PWM2/n25_neg_lutinv ),
    .c(\PWM2/n26 [8]),
    .d(\PWM2/pnumr [8]),
    .o(_al_u1859_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u186 (
    .a(pwm_state_read[13]),
    .b(pwm_start_stop[29]),
    .o(\PWMD/n11 ));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1860 (
    .a(_al_u1859_o),
    .b(\PWM2/n24 ),
    .c(pnumcnt2[8]),
    .d(\PWM2/pnumr [8]),
    .e(pwm_start_stop[18]),
    .o(\PWM2/n31 [8]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1861 (
    .a(\PWM2/n24 ),
    .b(\PWM2/n25_neg_lutinv ),
    .c(\PWM2/n26 [7]),
    .d(\PWM2/pnumr [7]),
    .o(_al_u1861_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1862 (
    .a(_al_u1861_o),
    .b(\PWM2/n24 ),
    .c(pnumcnt2[7]),
    .d(\PWM2/pnumr [7]),
    .e(pwm_start_stop[18]),
    .o(\PWM2/n31 [7]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1863 (
    .a(\PWM2/n24 ),
    .b(\PWM2/n25_neg_lutinv ),
    .c(\PWM2/n26 [6]),
    .d(\PWM2/pnumr [6]),
    .o(_al_u1863_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1864 (
    .a(_al_u1863_o),
    .b(\PWM2/n24 ),
    .c(pnumcnt2[6]),
    .d(\PWM2/pnumr [6]),
    .e(pwm_start_stop[18]),
    .o(\PWM2/n31 [6]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1865 (
    .a(\PWM2/n24 ),
    .b(\PWM2/n25_neg_lutinv ),
    .c(\PWM2/n26 [5]),
    .d(\PWM2/pnumr [5]),
    .o(_al_u1865_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1866 (
    .a(_al_u1865_o),
    .b(\PWM2/n24 ),
    .c(pnumcnt2[5]),
    .d(\PWM2/pnumr [5]),
    .e(pwm_start_stop[18]),
    .o(\PWM2/n31 [5]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1867 (
    .a(\PWM2/n24 ),
    .b(\PWM2/n25_neg_lutinv ),
    .c(\PWM2/n26 [4]),
    .d(\PWM2/pnumr [4]),
    .o(_al_u1867_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1868 (
    .a(_al_u1867_o),
    .b(\PWM2/n24 ),
    .c(pnumcnt2[4]),
    .d(\PWM2/pnumr [4]),
    .e(pwm_start_stop[18]),
    .o(\PWM2/n31 [4]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1869 (
    .a(\PWM2/n24 ),
    .b(\PWM2/n25_neg_lutinv ),
    .c(\PWM2/n26 [3]),
    .d(\PWM2/pnumr [3]),
    .o(_al_u1869_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u187 (
    .a(pwm_state_read[14]),
    .b(pwm_start_stop[30]),
    .o(\PWME/n11 ));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1870 (
    .a(_al_u1869_o),
    .b(\PWM2/n24 ),
    .c(pnumcnt2[3]),
    .d(\PWM2/pnumr [3]),
    .e(pwm_start_stop[18]),
    .o(\PWM2/n31 [3]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1871 (
    .a(\PWM2/n24 ),
    .b(\PWM2/n25_neg_lutinv ),
    .c(\PWM2/n26 [23]),
    .d(\PWM2/pnumr [23]),
    .o(_al_u1871_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1872 (
    .a(_al_u1871_o),
    .b(\PWM2/n24 ),
    .c(pnumcnt2[23]),
    .d(\PWM2/pnumr [23]),
    .e(pwm_start_stop[18]),
    .o(\PWM2/n31 [23]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1873 (
    .a(\PWM2/n24 ),
    .b(\PWM2/n25_neg_lutinv ),
    .c(\PWM2/n26 [22]),
    .d(\PWM2/pnumr [22]),
    .o(_al_u1873_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1874 (
    .a(_al_u1873_o),
    .b(\PWM2/n24 ),
    .c(pnumcnt2[22]),
    .d(\PWM2/pnumr [22]),
    .e(pwm_start_stop[18]),
    .o(\PWM2/n31 [22]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1875 (
    .a(\PWM2/n24 ),
    .b(\PWM2/n25_neg_lutinv ),
    .c(\PWM2/n26 [21]),
    .d(\PWM2/pnumr [21]),
    .o(_al_u1875_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1876 (
    .a(_al_u1875_o),
    .b(\PWM2/n24 ),
    .c(pnumcnt2[21]),
    .d(\PWM2/pnumr [21]),
    .e(pwm_start_stop[18]),
    .o(\PWM2/n31 [21]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1877 (
    .a(\PWM2/n24 ),
    .b(\PWM2/n25_neg_lutinv ),
    .c(\PWM2/n26 [20]),
    .d(\PWM2/pnumr [20]),
    .o(_al_u1877_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1878 (
    .a(_al_u1877_o),
    .b(\PWM2/n24 ),
    .c(pnumcnt2[20]),
    .d(\PWM2/pnumr [20]),
    .e(pwm_start_stop[18]),
    .o(\PWM2/n31 [20]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1879 (
    .a(\PWM2/n24 ),
    .b(\PWM2/n25_neg_lutinv ),
    .c(\PWM2/n26 [2]),
    .d(\PWM2/pnumr [2]),
    .o(_al_u1879_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u188 (
    .a(pwm_state_read[15]),
    .b(pwm_start_stop[31]),
    .o(\PWMF/n11 ));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1880 (
    .a(_al_u1879_o),
    .b(\PWM2/n24 ),
    .c(pnumcnt2[2]),
    .d(\PWM2/pnumr [2]),
    .e(pwm_start_stop[18]),
    .o(\PWM2/n31 [2]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1881 (
    .a(\PWM2/n24 ),
    .b(\PWM2/n25_neg_lutinv ),
    .c(\PWM2/n26 [19]),
    .d(\PWM2/pnumr [19]),
    .o(_al_u1881_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1882 (
    .a(_al_u1881_o),
    .b(\PWM2/n24 ),
    .c(pnumcnt2[19]),
    .d(\PWM2/pnumr [19]),
    .e(pwm_start_stop[18]),
    .o(\PWM2/n31 [19]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1883 (
    .a(\PWM2/n24 ),
    .b(\PWM2/n25_neg_lutinv ),
    .c(\PWM2/n26 [18]),
    .d(\PWM2/pnumr [18]),
    .o(_al_u1883_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1884 (
    .a(_al_u1883_o),
    .b(\PWM2/n24 ),
    .c(pnumcnt2[18]),
    .d(\PWM2/pnumr [18]),
    .e(pwm_start_stop[18]),
    .o(\PWM2/n31 [18]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1885 (
    .a(\PWM2/n24 ),
    .b(\PWM2/n25_neg_lutinv ),
    .c(\PWM2/n26 [17]),
    .d(\PWM2/pnumr [17]),
    .o(_al_u1885_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1886 (
    .a(_al_u1885_o),
    .b(\PWM2/n24 ),
    .c(pnumcnt2[17]),
    .d(\PWM2/pnumr [17]),
    .e(pwm_start_stop[18]),
    .o(\PWM2/n31 [17]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1887 (
    .a(\PWM2/n24 ),
    .b(\PWM2/n25_neg_lutinv ),
    .c(\PWM2/n26 [16]),
    .d(\PWM2/pnumr [16]),
    .o(_al_u1887_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1888 (
    .a(_al_u1887_o),
    .b(\PWM2/n24 ),
    .c(pnumcnt2[16]),
    .d(\PWM2/pnumr [16]),
    .e(pwm_start_stop[18]),
    .o(\PWM2/n31 [16]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1889 (
    .a(\PWM2/n24 ),
    .b(\PWM2/n25_neg_lutinv ),
    .c(\PWM2/n26 [15]),
    .d(\PWM2/pnumr [15]),
    .o(_al_u1889_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u189 (
    .a(\PWM0/pnumr [9]),
    .b(pnum0[32]),
    .c(pnum0[9]),
    .d(pwm_start_stop[16]),
    .o(\PWM0/n23 [9]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1890 (
    .a(_al_u1889_o),
    .b(\PWM2/n24 ),
    .c(pnumcnt2[15]),
    .d(\PWM2/pnumr [15]),
    .e(pwm_start_stop[18]),
    .o(\PWM2/n31 [15]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1891 (
    .a(\PWM2/n24 ),
    .b(\PWM2/n25_neg_lutinv ),
    .c(\PWM2/n26 [14]),
    .d(\PWM2/pnumr [14]),
    .o(_al_u1891_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1892 (
    .a(_al_u1891_o),
    .b(\PWM2/n24 ),
    .c(pnumcnt2[14]),
    .d(\PWM2/pnumr [14]),
    .e(pwm_start_stop[18]),
    .o(\PWM2/n31 [14]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1893 (
    .a(\PWM2/n24 ),
    .b(\PWM2/n25_neg_lutinv ),
    .c(\PWM2/n26 [13]),
    .d(\PWM2/pnumr [13]),
    .o(_al_u1893_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1894 (
    .a(_al_u1893_o),
    .b(\PWM2/n24 ),
    .c(pnumcnt2[13]),
    .d(\PWM2/pnumr [13]),
    .e(pwm_start_stop[18]),
    .o(\PWM2/n31 [13]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1895 (
    .a(\PWM2/n24 ),
    .b(\PWM2/n25_neg_lutinv ),
    .c(\PWM2/n26 [12]),
    .d(\PWM2/pnumr [12]),
    .o(_al_u1895_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1896 (
    .a(_al_u1895_o),
    .b(\PWM2/n24 ),
    .c(pnumcnt2[12]),
    .d(\PWM2/pnumr [12]),
    .e(pwm_start_stop[18]),
    .o(\PWM2/n31 [12]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1897 (
    .a(\PWM2/n24 ),
    .b(\PWM2/n25_neg_lutinv ),
    .c(\PWM2/n26 [11]),
    .d(\PWM2/pnumr [11]),
    .o(_al_u1897_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1898 (
    .a(_al_u1897_o),
    .b(\PWM2/n24 ),
    .c(pnumcnt2[11]),
    .d(\PWM2/pnumr [11]),
    .e(pwm_start_stop[18]),
    .o(\PWM2/n31 [11]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1899 (
    .a(\PWM2/n24 ),
    .b(\PWM2/n25_neg_lutinv ),
    .c(\PWM2/n26 [10]),
    .d(\PWM2/pnumr [10]),
    .o(_al_u1899_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u190 (
    .a(\PWM0/pnumr [8]),
    .b(pnum0[32]),
    .c(pnum0[8]),
    .d(pwm_start_stop[16]),
    .o(\PWM0/n23 [8]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1900 (
    .a(_al_u1899_o),
    .b(\PWM2/n24 ),
    .c(pnumcnt2[10]),
    .d(\PWM2/pnumr [10]),
    .e(pwm_start_stop[18]),
    .o(\PWM2/n31 [10]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1901 (
    .a(\PWM2/n24 ),
    .b(\PWM2/n25_neg_lutinv ),
    .c(\PWM2/n26 [1]),
    .d(\PWM2/pnumr [1]),
    .o(_al_u1901_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1902 (
    .a(_al_u1901_o),
    .b(\PWM2/n24 ),
    .c(pnumcnt2[1]),
    .d(\PWM2/pnumr [1]),
    .e(pwm_start_stop[18]),
    .o(\PWM2/n31 [1]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1903 (
    .a(\PWM2/n24 ),
    .b(\PWM2/n25_neg_lutinv ),
    .c(\PWM2/n26 [0]),
    .d(\PWM2/pnumr [0]),
    .o(_al_u1903_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1904 (
    .a(_al_u1903_o),
    .b(\PWM2/n24 ),
    .c(pnumcnt2[0]),
    .d(\PWM2/pnumr [0]),
    .e(pwm_start_stop[18]),
    .o(\PWM2/n31 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u1905 (
    .a(\PWM2/FreCnt [19]),
    .b(\PWM2/FreCnt [8]),
    .c(\PWM2/FreCntr [20]),
    .d(\PWM2/FreCntr [9]),
    .o(_al_u1905_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*~C)*~(D*~B))"),
    .INIT(32'h80a088aa))
    _al_u1906 (
    .a(_al_u1905_o),
    .b(\PWM2/FreCnt [17]),
    .c(\PWM2/FreCnt [25]),
    .d(\PWM2/FreCntr [18]),
    .e(\PWM2/FreCntr [26]),
    .o(_al_u1906_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u1907 (
    .a(\PWM2/FreCnt [21]),
    .b(\PWM2/FreCnt [5]),
    .c(\PWM2/FreCntr [22]),
    .d(\PWM2/FreCntr [6]),
    .o(_al_u1907_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(~D*C))"),
    .INIT(16'h8808))
    _al_u1908 (
    .a(_al_u1906_o),
    .b(_al_u1907_o),
    .c(\PWM2/FreCnt [10]),
    .d(\PWM2/FreCntr [11]),
    .o(_al_u1908_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u1909 (
    .a(\PWM2/FreCnt [3]),
    .b(\PWM2/FreCnt [7]),
    .c(\PWM2/FreCntr [4]),
    .d(\PWM2/FreCntr [8]),
    .o(_al_u1909_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u191 (
    .a(\PWM0/pnumr [7]),
    .b(pnum0[32]),
    .c(pnum0[7]),
    .d(pwm_start_stop[16]),
    .o(\PWM0/n23 [7]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*C)*~(D*~B))"),
    .INIT(32'h88aa080a))
    _al_u1910 (
    .a(_al_u1909_o),
    .b(\PWM2/FreCnt [10]),
    .c(\PWM2/FreCnt [25]),
    .d(\PWM2/FreCntr [11]),
    .e(\PWM2/FreCntr [26]),
    .o(_al_u1910_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u1911 (
    .a(\PWM2/FreCnt [1]),
    .b(\PWM2/FreCnt [5]),
    .c(\PWM2/FreCntr [2]),
    .d(\PWM2/FreCntr [6]),
    .o(_al_u1911_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u1912 (
    .a(_al_u1908_o),
    .b(_al_u1910_o),
    .c(_al_u1911_o),
    .d(\PWM2/FreCnt [16]),
    .e(\PWM2/FreCntr [17]),
    .o(_al_u1912_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1913 (
    .a(\PWM2/FreCnt [15]),
    .b(\PWM2/FreCntr [16]),
    .o(_al_u1913_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(E*~C)*~(D@B))"),
    .INIT(32'h40104411))
    _al_u1914 (
    .a(_al_u1913_o),
    .b(\PWM2/FreCnt [20]),
    .c(\PWM2/FreCnt [23]),
    .d(\PWM2/FreCntr [21]),
    .e(\PWM2/FreCntr [24]),
    .o(_al_u1914_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D@C)*~(E@B))"),
    .INIT(32'h80082002))
    _al_u1915 (
    .a(_al_u1914_o),
    .b(\PWM2/FreCnt [13]),
    .c(\PWM2/FreCnt [9]),
    .d(\PWM2/FreCntr [10]),
    .e(\PWM2/FreCntr [14]),
    .o(_al_u1915_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u1916 (
    .a(\PWM2/FreCnt [1]),
    .b(\PWM2/FreCnt [23]),
    .c(\PWM2/FreCntr [2]),
    .d(\PWM2/FreCntr [24]),
    .o(_al_u1916_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*~C)*~(~D*B))"),
    .INIT(32'ha020aa22))
    _al_u1917 (
    .a(_al_u1916_o),
    .b(\PWM2/FreCnt [15]),
    .c(\PWM2/FreCnt [21]),
    .d(\PWM2/FreCntr [16]),
    .e(\PWM2/FreCntr [22]),
    .o(_al_u1917_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u1918 (
    .a(\PWM2/FreCnt [7]),
    .b(\PWM2/FreCnt [8]),
    .c(\PWM2/FreCntr [8]),
    .d(\PWM2/FreCntr [9]),
    .o(_al_u1918_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u1919 (
    .a(_al_u1915_o),
    .b(_al_u1917_o),
    .c(_al_u1918_o),
    .d(\PWM2/FreCnt [12]),
    .e(\PWM2/FreCntr [13]),
    .o(_al_u1919_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u192 (
    .a(\PWM0/pnumr [6]),
    .b(pnum0[32]),
    .c(pnum0[6]),
    .d(pwm_start_stop[16]),
    .o(\PWM0/n23 [6]));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1920 (
    .a(\PWM2/FreCnt [0]),
    .b(\PWM2/FreCnt [18]),
    .c(\PWM2/FreCntr [1]),
    .d(\PWM2/FreCntr [19]),
    .o(_al_u1920_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u1921 (
    .a(_al_u1920_o),
    .b(\PWM2/FreCnt [4]),
    .c(\PWM2/FreCntr [5]),
    .o(_al_u1921_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1922 (
    .a(\PWM2/FreCnt [24]),
    .b(\PWM2/FreCnt [6]),
    .c(\PWM2/FreCntr [25]),
    .d(\PWM2/FreCntr [7]),
    .o(_al_u1922_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1923 (
    .a(_al_u1922_o),
    .b(\PWM2/FreCnt [14]),
    .c(\PWM2/FreCnt [2]),
    .d(\PWM2/FreCntr [15]),
    .e(\PWM2/FreCntr [3]),
    .o(_al_u1923_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u1924 (
    .a(\PWM2/FreCnt [17]),
    .b(\PWM2/FreCnt [3]),
    .c(\PWM2/FreCntr [18]),
    .d(\PWM2/FreCntr [4]),
    .o(_al_u1924_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*C)*~(D*~B))"),
    .INIT(32'h88aa080a))
    _al_u1925 (
    .a(_al_u1924_o),
    .b(\PWM2/FreCnt [11]),
    .c(\PWM2/FreCnt [19]),
    .d(\PWM2/FreCntr [12]),
    .e(\PWM2/FreCntr [20]),
    .o(_al_u1925_o));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(E@B)*~(~D*A))"),
    .INIT(32'h0c040301))
    _al_u1926 (
    .a(\PWM2/FreCnt [11]),
    .b(\PWM2/FreCnt [22]),
    .c(\PWM2/FreCnt [26]),
    .d(\PWM2/FreCntr [12]),
    .e(\PWM2/FreCntr [23]),
    .o(_al_u1926_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1927 (
    .a(_al_u1921_o),
    .b(_al_u1923_o),
    .c(_al_u1925_o),
    .d(_al_u1926_o),
    .o(_al_u1927_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*A))"),
    .INIT(16'h7f00))
    _al_u1928 (
    .a(_al_u1912_o),
    .b(_al_u1919_o),
    .c(_al_u1927_o),
    .d(pwm_state_read[2]),
    .o(\PWM2/u14_sel_is_1_o ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1929 (
    .a(\PWM3/n0_lutinv ),
    .b(pwm_state_read[3]),
    .o(\PWM3/n24 ));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u193 (
    .a(\PWM0/pnumr [5]),
    .b(pnum0[32]),
    .c(pnum0[5]),
    .d(pwm_start_stop[16]),
    .o(\PWM0/n23 [5]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1930 (
    .a(pnumcnt3[18]),
    .b(pnumcnt3[19]),
    .c(pnumcnt3[1]),
    .d(pnumcnt3[20]),
    .o(_al_u1930_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u1931 (
    .a(_al_u1930_o),
    .b(pnumcnt3[21]),
    .c(pnumcnt3[22]),
    .d(pnumcnt3[23]),
    .e(pnumcnt3[2]),
    .o(_al_u1931_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u1932 (
    .a(_al_u1931_o),
    .b(pnumcnt3[6]),
    .c(pnumcnt3[7]),
    .d(pnumcnt3[8]),
    .e(pnumcnt3[9]),
    .o(_al_u1932_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u1933 (
    .a(pnumcnt3[10]),
    .b(pnumcnt3[11]),
    .c(pnumcnt3[12]),
    .d(pnumcnt3[13]),
    .o(_al_u1933_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u1934 (
    .a(_al_u1933_o),
    .b(pnumcnt3[14]),
    .c(pnumcnt3[15]),
    .d(pnumcnt3[16]),
    .e(pnumcnt3[17]),
    .o(_al_u1934_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u1935 (
    .a(pnumcnt3[3]),
    .b(pnumcnt3[4]),
    .c(pnumcnt3[5]),
    .o(_al_u1935_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u1936 (
    .a(_al_u1932_o),
    .b(_al_u1934_o),
    .c(_al_u1935_o),
    .d(pnumcnt3[0]),
    .o(\PWM3/n25_neg_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1937 (
    .a(\PWM3/n24 ),
    .b(\PWM3/n25_neg_lutinv ),
    .c(\PWM3/n26 [9]),
    .d(\PWM3/pnumr [9]),
    .o(_al_u1937_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1938 (
    .a(_al_u1937_o),
    .b(\PWM3/n24 ),
    .c(pnumcnt3[9]),
    .d(\PWM3/pnumr [9]),
    .e(pwm_start_stop[19]),
    .o(\PWM3/n31 [9]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1939 (
    .a(\PWM3/n24 ),
    .b(\PWM3/n25_neg_lutinv ),
    .c(\PWM3/n26 [8]),
    .d(\PWM3/pnumr [8]),
    .o(_al_u1939_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u194 (
    .a(\PWM0/pnumr [4]),
    .b(pnum0[32]),
    .c(pnum0[4]),
    .d(pwm_start_stop[16]),
    .o(\PWM0/n23 [4]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1940 (
    .a(_al_u1939_o),
    .b(\PWM3/n24 ),
    .c(pnumcnt3[8]),
    .d(\PWM3/pnumr [8]),
    .e(pwm_start_stop[19]),
    .o(\PWM3/n31 [8]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1941 (
    .a(\PWM3/n24 ),
    .b(\PWM3/n25_neg_lutinv ),
    .c(\PWM3/n26 [7]),
    .d(\PWM3/pnumr [7]),
    .o(_al_u1941_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1942 (
    .a(_al_u1941_o),
    .b(\PWM3/n24 ),
    .c(pnumcnt3[7]),
    .d(\PWM3/pnumr [7]),
    .e(pwm_start_stop[19]),
    .o(\PWM3/n31 [7]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1943 (
    .a(\PWM3/n24 ),
    .b(\PWM3/n25_neg_lutinv ),
    .c(\PWM3/n26 [6]),
    .d(\PWM3/pnumr [6]),
    .o(_al_u1943_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1944 (
    .a(_al_u1943_o),
    .b(\PWM3/n24 ),
    .c(pnumcnt3[6]),
    .d(\PWM3/pnumr [6]),
    .e(pwm_start_stop[19]),
    .o(\PWM3/n31 [6]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1945 (
    .a(\PWM3/n24 ),
    .b(\PWM3/n25_neg_lutinv ),
    .c(\PWM3/n26 [5]),
    .d(\PWM3/pnumr [5]),
    .o(_al_u1945_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1946 (
    .a(_al_u1945_o),
    .b(\PWM3/n24 ),
    .c(pnumcnt3[5]),
    .d(\PWM3/pnumr [5]),
    .e(pwm_start_stop[19]),
    .o(\PWM3/n31 [5]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1947 (
    .a(\PWM3/n24 ),
    .b(\PWM3/n25_neg_lutinv ),
    .c(\PWM3/n26 [4]),
    .d(\PWM3/pnumr [4]),
    .o(_al_u1947_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1948 (
    .a(_al_u1947_o),
    .b(\PWM3/n24 ),
    .c(pnumcnt3[4]),
    .d(\PWM3/pnumr [4]),
    .e(pwm_start_stop[19]),
    .o(\PWM3/n31 [4]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1949 (
    .a(\PWM3/n24 ),
    .b(\PWM3/n25_neg_lutinv ),
    .c(\PWM3/n26 [3]),
    .d(\PWM3/pnumr [3]),
    .o(_al_u1949_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u195 (
    .a(\PWM0/pnumr [31]),
    .b(pnum0[31]),
    .c(pnum0[32]),
    .d(pwm_start_stop[16]),
    .o(\PWM0/n23 [31]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1950 (
    .a(_al_u1949_o),
    .b(\PWM3/n24 ),
    .c(pnumcnt3[3]),
    .d(\PWM3/pnumr [3]),
    .e(pwm_start_stop[19]),
    .o(\PWM3/n31 [3]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1951 (
    .a(\PWM3/n24 ),
    .b(\PWM3/n25_neg_lutinv ),
    .c(\PWM3/n26 [23]),
    .d(\PWM3/pnumr [23]),
    .o(_al_u1951_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1952 (
    .a(_al_u1951_o),
    .b(\PWM3/n24 ),
    .c(pnumcnt3[23]),
    .d(\PWM3/pnumr [23]),
    .e(pwm_start_stop[19]),
    .o(\PWM3/n31 [23]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1953 (
    .a(\PWM3/n24 ),
    .b(\PWM3/n25_neg_lutinv ),
    .c(\PWM3/n26 [22]),
    .d(\PWM3/pnumr [22]),
    .o(_al_u1953_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1954 (
    .a(_al_u1953_o),
    .b(\PWM3/n24 ),
    .c(pnumcnt3[22]),
    .d(\PWM3/pnumr [22]),
    .e(pwm_start_stop[19]),
    .o(\PWM3/n31 [22]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1955 (
    .a(\PWM3/n24 ),
    .b(\PWM3/n25_neg_lutinv ),
    .c(\PWM3/n26 [21]),
    .d(\PWM3/pnumr [21]),
    .o(_al_u1955_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1956 (
    .a(_al_u1955_o),
    .b(\PWM3/n24 ),
    .c(pnumcnt3[21]),
    .d(\PWM3/pnumr [21]),
    .e(pwm_start_stop[19]),
    .o(\PWM3/n31 [21]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1957 (
    .a(\PWM3/n24 ),
    .b(\PWM3/n25_neg_lutinv ),
    .c(\PWM3/n26 [20]),
    .d(\PWM3/pnumr [20]),
    .o(_al_u1957_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1958 (
    .a(_al_u1957_o),
    .b(\PWM3/n24 ),
    .c(pnumcnt3[20]),
    .d(\PWM3/pnumr [20]),
    .e(pwm_start_stop[19]),
    .o(\PWM3/n31 [20]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1959 (
    .a(\PWM3/n24 ),
    .b(\PWM3/n25_neg_lutinv ),
    .c(\PWM3/n26 [2]),
    .d(\PWM3/pnumr [2]),
    .o(_al_u1959_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u196 (
    .a(\PWM0/pnumr [30]),
    .b(pnum0[30]),
    .c(pnum0[32]),
    .d(pwm_start_stop[16]),
    .o(\PWM0/n23 [30]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1960 (
    .a(_al_u1959_o),
    .b(\PWM3/n24 ),
    .c(pnumcnt3[2]),
    .d(\PWM3/pnumr [2]),
    .e(pwm_start_stop[19]),
    .o(\PWM3/n31 [2]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1961 (
    .a(\PWM3/n24 ),
    .b(\PWM3/n25_neg_lutinv ),
    .c(\PWM3/n26 [19]),
    .d(\PWM3/pnumr [19]),
    .o(_al_u1961_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1962 (
    .a(_al_u1961_o),
    .b(\PWM3/n24 ),
    .c(pnumcnt3[19]),
    .d(\PWM3/pnumr [19]),
    .e(pwm_start_stop[19]),
    .o(\PWM3/n31 [19]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1963 (
    .a(\PWM3/n24 ),
    .b(\PWM3/n25_neg_lutinv ),
    .c(\PWM3/n26 [18]),
    .d(\PWM3/pnumr [18]),
    .o(_al_u1963_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1964 (
    .a(_al_u1963_o),
    .b(\PWM3/n24 ),
    .c(pnumcnt3[18]),
    .d(\PWM3/pnumr [18]),
    .e(pwm_start_stop[19]),
    .o(\PWM3/n31 [18]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1965 (
    .a(\PWM3/n24 ),
    .b(\PWM3/n25_neg_lutinv ),
    .c(\PWM3/n26 [17]),
    .d(\PWM3/pnumr [17]),
    .o(_al_u1965_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1966 (
    .a(_al_u1965_o),
    .b(\PWM3/n24 ),
    .c(pnumcnt3[17]),
    .d(\PWM3/pnumr [17]),
    .e(pwm_start_stop[19]),
    .o(\PWM3/n31 [17]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1967 (
    .a(\PWM3/n24 ),
    .b(\PWM3/n25_neg_lutinv ),
    .c(\PWM3/n26 [16]),
    .d(\PWM3/pnumr [16]),
    .o(_al_u1967_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1968 (
    .a(_al_u1967_o),
    .b(\PWM3/n24 ),
    .c(pnumcnt3[16]),
    .d(\PWM3/pnumr [16]),
    .e(pwm_start_stop[19]),
    .o(\PWM3/n31 [16]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1969 (
    .a(\PWM3/n24 ),
    .b(\PWM3/n25_neg_lutinv ),
    .c(\PWM3/n26 [15]),
    .d(\PWM3/pnumr [15]),
    .o(_al_u1969_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u197 (
    .a(\PWM0/pnumr [3]),
    .b(pnum0[3]),
    .c(pnum0[32]),
    .d(pwm_start_stop[16]),
    .o(\PWM0/n23 [3]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1970 (
    .a(_al_u1969_o),
    .b(\PWM3/n24 ),
    .c(pnumcnt3[15]),
    .d(\PWM3/pnumr [15]),
    .e(pwm_start_stop[19]),
    .o(\PWM3/n31 [15]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1971 (
    .a(\PWM3/n24 ),
    .b(\PWM3/n25_neg_lutinv ),
    .c(\PWM3/n26 [14]),
    .d(\PWM3/pnumr [14]),
    .o(_al_u1971_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1972 (
    .a(_al_u1971_o),
    .b(\PWM3/n24 ),
    .c(pnumcnt3[14]),
    .d(\PWM3/pnumr [14]),
    .e(pwm_start_stop[19]),
    .o(\PWM3/n31 [14]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1973 (
    .a(\PWM3/n24 ),
    .b(\PWM3/n25_neg_lutinv ),
    .c(\PWM3/n26 [13]),
    .d(\PWM3/pnumr [13]),
    .o(_al_u1973_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1974 (
    .a(_al_u1973_o),
    .b(\PWM3/n24 ),
    .c(pnumcnt3[13]),
    .d(\PWM3/pnumr [13]),
    .e(pwm_start_stop[19]),
    .o(\PWM3/n31 [13]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1975 (
    .a(\PWM3/n24 ),
    .b(\PWM3/n25_neg_lutinv ),
    .c(\PWM3/n26 [12]),
    .d(\PWM3/pnumr [12]),
    .o(_al_u1975_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1976 (
    .a(_al_u1975_o),
    .b(\PWM3/n24 ),
    .c(pnumcnt3[12]),
    .d(\PWM3/pnumr [12]),
    .e(pwm_start_stop[19]),
    .o(\PWM3/n31 [12]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1977 (
    .a(\PWM3/n24 ),
    .b(\PWM3/n25_neg_lutinv ),
    .c(\PWM3/n26 [11]),
    .d(\PWM3/pnumr [11]),
    .o(_al_u1977_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1978 (
    .a(_al_u1977_o),
    .b(\PWM3/n24 ),
    .c(pnumcnt3[11]),
    .d(\PWM3/pnumr [11]),
    .e(pwm_start_stop[19]),
    .o(\PWM3/n31 [11]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1979 (
    .a(\PWM3/n24 ),
    .b(\PWM3/n25_neg_lutinv ),
    .c(\PWM3/n26 [10]),
    .d(\PWM3/pnumr [10]),
    .o(_al_u1979_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u198 (
    .a(\PWM0/pnumr [29]),
    .b(pnum0[29]),
    .c(pnum0[32]),
    .d(pwm_start_stop[16]),
    .o(\PWM0/n23 [29]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1980 (
    .a(_al_u1979_o),
    .b(\PWM3/n24 ),
    .c(pnumcnt3[10]),
    .d(\PWM3/pnumr [10]),
    .e(pwm_start_stop[19]),
    .o(\PWM3/n31 [10]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1981 (
    .a(\PWM3/n24 ),
    .b(\PWM3/n25_neg_lutinv ),
    .c(\PWM3/n26 [1]),
    .d(\PWM3/pnumr [1]),
    .o(_al_u1981_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1982 (
    .a(_al_u1981_o),
    .b(\PWM3/n24 ),
    .c(pnumcnt3[1]),
    .d(\PWM3/pnumr [1]),
    .e(pwm_start_stop[19]),
    .o(\PWM3/n31 [1]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u1983 (
    .a(\PWM3/n24 ),
    .b(\PWM3/n25_neg_lutinv ),
    .c(\PWM3/n26 [0]),
    .d(\PWM3/pnumr [0]),
    .o(_al_u1983_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u1984 (
    .a(_al_u1983_o),
    .b(\PWM3/n24 ),
    .c(pnumcnt3[0]),
    .d(\PWM3/pnumr [0]),
    .e(pwm_start_stop[19]),
    .o(\PWM3/n31 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1985 (
    .a(\PWM3/FreCnt [0]),
    .b(\PWM3/FreCnt [22]),
    .c(\PWM3/FreCntr [1]),
    .d(\PWM3/FreCntr [23]),
    .o(_al_u1985_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u1986 (
    .a(_al_u1985_o),
    .b(\PWM3/FreCnt [2]),
    .c(\PWM3/FreCntr [3]),
    .o(_al_u1986_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u1987 (
    .a(\PWM3/FreCnt [14]),
    .b(\PWM3/FreCnt [24]),
    .c(\PWM3/FreCntr [15]),
    .d(\PWM3/FreCntr [25]),
    .o(_al_u1987_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u1988 (
    .a(_al_u1987_o),
    .b(\PWM3/FreCnt [4]),
    .c(\PWM3/FreCnt [5]),
    .d(\PWM3/FreCntr [5]),
    .e(\PWM3/FreCntr [6]),
    .o(_al_u1988_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u1989 (
    .a(\PWM3/FreCnt [1]),
    .b(\PWM3/FreCnt [3]),
    .c(\PWM3/FreCntr [2]),
    .d(\PWM3/FreCntr [4]),
    .o(_al_u1989_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u199 (
    .a(\PWM0/pnumr [28]),
    .b(pnum0[28]),
    .c(pnum0[32]),
    .d(pwm_start_stop[16]),
    .o(\PWM0/n23 [28]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*C)*~(D*~B))"),
    .INIT(32'h88aa080a))
    _al_u1990 (
    .a(_al_u1989_o),
    .b(\PWM3/FreCnt [12]),
    .c(\PWM3/FreCnt [25]),
    .d(\PWM3/FreCntr [13]),
    .e(\PWM3/FreCntr [26]),
    .o(_al_u1990_o));
  AL_MAP_LUT5 #(
    .EQN("(~B*~(E@C)*~(~D*A))"),
    .INIT(32'h30100301))
    _al_u1991 (
    .a(\PWM3/FreCnt [21]),
    .b(\PWM3/FreCnt [26]),
    .c(\PWM3/FreCnt [8]),
    .d(\PWM3/FreCntr [22]),
    .e(\PWM3/FreCntr [9]),
    .o(_al_u1991_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1992 (
    .a(_al_u1986_o),
    .b(_al_u1988_o),
    .c(_al_u1990_o),
    .d(_al_u1991_o),
    .o(_al_u1992_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C@A))"),
    .INIT(16'ha521))
    _al_u1993 (
    .a(\PWM3/FreCnt [6]),
    .b(\PWM3/FreCnt [7]),
    .c(\PWM3/FreCntr [7]),
    .d(\PWM3/FreCntr [8]),
    .o(_al_u1993_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u1994 (
    .a(\PWM3/FreCnt [13]),
    .b(\PWM3/FreCnt [7]),
    .c(\PWM3/FreCntr [14]),
    .d(\PWM3/FreCntr [8]),
    .o(_al_u1994_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D@C))"),
    .INIT(16'h8008))
    _al_u1995 (
    .a(_al_u1993_o),
    .b(_al_u1994_o),
    .c(\PWM3/FreCnt [10]),
    .d(\PWM3/FreCntr [11]),
    .o(_al_u1995_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1996 (
    .a(\PWM3/FreCnt [12]),
    .b(\PWM3/FreCntr [13]),
    .o(_al_u1996_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(~D*C)*~(E@B))"),
    .INIT(32'h44041101))
    _al_u1997 (
    .a(_al_u1996_o),
    .b(\PWM3/FreCnt [20]),
    .c(\PWM3/FreCnt [9]),
    .d(\PWM3/FreCntr [10]),
    .e(\PWM3/FreCntr [21]),
    .o(_al_u1997_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1998 (
    .a(\PWM3/FreCnt [9]),
    .b(\PWM3/FreCntr [10]),
    .o(_al_u1998_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(E@C)*~(D*~B))"),
    .INIT(32'h40500405))
    _al_u1999 (
    .a(_al_u1998_o),
    .b(\PWM3/FreCnt [16]),
    .c(\PWM3/FreCnt [18]),
    .d(\PWM3/FreCntr [17]),
    .e(\PWM3/FreCntr [19]),
    .o(_al_u1999_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u200 (
    .a(\PWM0/pnumr [27]),
    .b(pnum0[27]),
    .c(pnum0[32]),
    .d(pwm_start_stop[16]),
    .o(\PWM0/n23 [27]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u2000 (
    .a(_al_u1995_o),
    .b(_al_u1997_o),
    .c(_al_u1999_o),
    .o(_al_u2000_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u2001 (
    .a(\PWM3/FreCnt [15]),
    .b(\PWM3/FreCnt [21]),
    .c(\PWM3/FreCntr [16]),
    .d(\PWM3/FreCntr [22]),
    .o(_al_u2001_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*~C)*~(D*~B))"),
    .INIT(32'h80a088aa))
    _al_u2002 (
    .a(_al_u2001_o),
    .b(\PWM3/FreCnt [13]),
    .c(\PWM3/FreCnt [19]),
    .d(\PWM3/FreCntr [14]),
    .e(\PWM3/FreCntr [20]),
    .o(_al_u2002_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u2003 (
    .a(\PWM3/FreCnt [25]),
    .b(\PWM3/FreCnt [3]),
    .c(\PWM3/FreCntr [26]),
    .d(\PWM3/FreCntr [4]),
    .o(_al_u2003_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D@C))"),
    .INIT(16'h8008))
    _al_u2004 (
    .a(_al_u2002_o),
    .b(_al_u2003_o),
    .c(\PWM3/FreCnt [11]),
    .d(\PWM3/FreCntr [12]),
    .o(_al_u2004_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2005 (
    .a(\PWM3/FreCnt [16]),
    .b(\PWM3/FreCntr [17]),
    .o(_al_u2005_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(~E*C)*~(D@B))"),
    .INIT(32'h44110401))
    _al_u2006 (
    .a(_al_u2005_o),
    .b(\PWM3/FreCnt [17]),
    .c(\PWM3/FreCnt [19]),
    .d(\PWM3/FreCntr [18]),
    .e(\PWM3/FreCntr [20]),
    .o(_al_u2006_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2007 (
    .a(\PWM3/FreCnt [1]),
    .b(\PWM3/FreCntr [2]),
    .o(_al_u2007_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(E@C)*~(D*~B))"),
    .INIT(32'h40500405))
    _al_u2008 (
    .a(_al_u2007_o),
    .b(\PWM3/FreCnt [15]),
    .c(\PWM3/FreCnt [23]),
    .d(\PWM3/FreCntr [16]),
    .e(\PWM3/FreCntr [24]),
    .o(_al_u2008_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    _al_u2009 (
    .a(_al_u1992_o),
    .b(_al_u2000_o),
    .c(_al_u2004_o),
    .d(_al_u2006_o),
    .e(_al_u2008_o),
    .o(_al_u2009_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u201 (
    .a(\PWM0/pnumr [26]),
    .b(pnum0[26]),
    .c(pnum0[32]),
    .d(pwm_start_stop[16]),
    .o(\PWM0/n23 [26]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2010 (
    .a(_al_u2009_o),
    .b(pwm_state_read[3]),
    .o(\PWM3/u14_sel_is_1_o ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2011 (
    .a(\PWM4/n0_lutinv ),
    .b(pwm_state_read[4]),
    .o(\PWM4/n24 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u2012 (
    .a(pnumcnt4[18]),
    .b(pnumcnt4[19]),
    .c(pnumcnt4[1]),
    .d(pnumcnt4[20]),
    .o(_al_u2012_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u2013 (
    .a(_al_u2012_o),
    .b(pnumcnt4[21]),
    .c(pnumcnt4[22]),
    .d(pnumcnt4[23]),
    .e(pnumcnt4[2]),
    .o(_al_u2013_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u2014 (
    .a(_al_u2013_o),
    .b(pnumcnt4[6]),
    .c(pnumcnt4[7]),
    .d(pnumcnt4[8]),
    .e(pnumcnt4[9]),
    .o(_al_u2014_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u2015 (
    .a(pnumcnt4[10]),
    .b(pnumcnt4[11]),
    .c(pnumcnt4[12]),
    .d(pnumcnt4[13]),
    .o(_al_u2015_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u2016 (
    .a(_al_u2015_o),
    .b(pnumcnt4[14]),
    .c(pnumcnt4[15]),
    .d(pnumcnt4[16]),
    .e(pnumcnt4[17]),
    .o(_al_u2016_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u2017 (
    .a(pnumcnt4[3]),
    .b(pnumcnt4[4]),
    .c(pnumcnt4[5]),
    .o(_al_u2017_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u2018 (
    .a(_al_u2014_o),
    .b(_al_u2016_o),
    .c(_al_u2017_o),
    .d(pnumcnt4[0]),
    .o(\PWM4/n25_neg_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2019 (
    .a(\PWM4/n24 ),
    .b(\PWM4/n25_neg_lutinv ),
    .c(\PWM4/n26 [9]),
    .d(\PWM4/pnumr [9]),
    .o(_al_u2019_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u202 (
    .a(\PWM0/pnumr [25]),
    .b(pnum0[25]),
    .c(pnum0[32]),
    .d(pwm_start_stop[16]),
    .o(\PWM0/n23 [25]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2020 (
    .a(_al_u2019_o),
    .b(\PWM4/n24 ),
    .c(pnumcnt4[9]),
    .d(\PWM4/pnumr [9]),
    .e(pwm_start_stop[20]),
    .o(\PWM4/n31 [9]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2021 (
    .a(\PWM4/n24 ),
    .b(\PWM4/n25_neg_lutinv ),
    .c(\PWM4/n26 [8]),
    .d(\PWM4/pnumr [8]),
    .o(_al_u2021_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2022 (
    .a(_al_u2021_o),
    .b(\PWM4/n24 ),
    .c(pnumcnt4[8]),
    .d(\PWM4/pnumr [8]),
    .e(pwm_start_stop[20]),
    .o(\PWM4/n31 [8]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2023 (
    .a(\PWM4/n24 ),
    .b(\PWM4/n25_neg_lutinv ),
    .c(\PWM4/n26 [7]),
    .d(\PWM4/pnumr [7]),
    .o(_al_u2023_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2024 (
    .a(_al_u2023_o),
    .b(\PWM4/n24 ),
    .c(pnumcnt4[7]),
    .d(\PWM4/pnumr [7]),
    .e(pwm_start_stop[20]),
    .o(\PWM4/n31 [7]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2025 (
    .a(\PWM4/n24 ),
    .b(\PWM4/n25_neg_lutinv ),
    .c(\PWM4/n26 [6]),
    .d(\PWM4/pnumr [6]),
    .o(_al_u2025_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2026 (
    .a(_al_u2025_o),
    .b(\PWM4/n24 ),
    .c(pnumcnt4[6]),
    .d(\PWM4/pnumr [6]),
    .e(pwm_start_stop[20]),
    .o(\PWM4/n31 [6]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2027 (
    .a(\PWM4/n24 ),
    .b(\PWM4/n25_neg_lutinv ),
    .c(\PWM4/n26 [5]),
    .d(\PWM4/pnumr [5]),
    .o(_al_u2027_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2028 (
    .a(_al_u2027_o),
    .b(\PWM4/n24 ),
    .c(pnumcnt4[5]),
    .d(\PWM4/pnumr [5]),
    .e(pwm_start_stop[20]),
    .o(\PWM4/n31 [5]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2029 (
    .a(\PWM4/n24 ),
    .b(\PWM4/n25_neg_lutinv ),
    .c(\PWM4/n26 [4]),
    .d(\PWM4/pnumr [4]),
    .o(_al_u2029_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u203 (
    .a(\PWM0/pnumr [24]),
    .b(pnum0[24]),
    .c(pnum0[32]),
    .d(pwm_start_stop[16]),
    .o(\PWM0/n23 [24]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2030 (
    .a(_al_u2029_o),
    .b(\PWM4/n24 ),
    .c(pnumcnt4[4]),
    .d(\PWM4/pnumr [4]),
    .e(pwm_start_stop[20]),
    .o(\PWM4/n31 [4]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2031 (
    .a(\PWM4/n24 ),
    .b(\PWM4/n25_neg_lutinv ),
    .c(\PWM4/n26 [3]),
    .d(\PWM4/pnumr [3]),
    .o(_al_u2031_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2032 (
    .a(_al_u2031_o),
    .b(\PWM4/n24 ),
    .c(pnumcnt4[3]),
    .d(\PWM4/pnumr [3]),
    .e(pwm_start_stop[20]),
    .o(\PWM4/n31 [3]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2033 (
    .a(\PWM4/n24 ),
    .b(\PWM4/n25_neg_lutinv ),
    .c(\PWM4/n26 [23]),
    .d(\PWM4/pnumr [23]),
    .o(_al_u2033_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2034 (
    .a(_al_u2033_o),
    .b(\PWM4/n24 ),
    .c(pnumcnt4[23]),
    .d(\PWM4/pnumr [23]),
    .e(pwm_start_stop[20]),
    .o(\PWM4/n31 [23]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2035 (
    .a(\PWM4/n24 ),
    .b(\PWM4/n25_neg_lutinv ),
    .c(\PWM4/n26 [22]),
    .d(\PWM4/pnumr [22]),
    .o(_al_u2035_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2036 (
    .a(_al_u2035_o),
    .b(\PWM4/n24 ),
    .c(pnumcnt4[22]),
    .d(\PWM4/pnumr [22]),
    .e(pwm_start_stop[20]),
    .o(\PWM4/n31 [22]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2037 (
    .a(\PWM4/n24 ),
    .b(\PWM4/n25_neg_lutinv ),
    .c(\PWM4/n26 [21]),
    .d(\PWM4/pnumr [21]),
    .o(_al_u2037_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2038 (
    .a(_al_u2037_o),
    .b(\PWM4/n24 ),
    .c(pnumcnt4[21]),
    .d(\PWM4/pnumr [21]),
    .e(pwm_start_stop[20]),
    .o(\PWM4/n31 [21]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2039 (
    .a(\PWM4/n24 ),
    .b(\PWM4/n25_neg_lutinv ),
    .c(\PWM4/n26 [20]),
    .d(\PWM4/pnumr [20]),
    .o(_al_u2039_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u204 (
    .a(\PWM0/pnumr [23]),
    .b(pnum0[23]),
    .c(pnum0[32]),
    .d(pwm_start_stop[16]),
    .o(\PWM0/n23 [23]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2040 (
    .a(_al_u2039_o),
    .b(\PWM4/n24 ),
    .c(pnumcnt4[20]),
    .d(\PWM4/pnumr [20]),
    .e(pwm_start_stop[20]),
    .o(\PWM4/n31 [20]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2041 (
    .a(\PWM4/n24 ),
    .b(\PWM4/n25_neg_lutinv ),
    .c(\PWM4/n26 [2]),
    .d(\PWM4/pnumr [2]),
    .o(_al_u2041_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2042 (
    .a(_al_u2041_o),
    .b(\PWM4/n24 ),
    .c(pnumcnt4[2]),
    .d(\PWM4/pnumr [2]),
    .e(pwm_start_stop[20]),
    .o(\PWM4/n31 [2]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2043 (
    .a(\PWM4/n24 ),
    .b(\PWM4/n25_neg_lutinv ),
    .c(\PWM4/n26 [19]),
    .d(\PWM4/pnumr [19]),
    .o(_al_u2043_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2044 (
    .a(_al_u2043_o),
    .b(\PWM4/n24 ),
    .c(pnumcnt4[19]),
    .d(\PWM4/pnumr [19]),
    .e(pwm_start_stop[20]),
    .o(\PWM4/n31 [19]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2045 (
    .a(\PWM4/n24 ),
    .b(\PWM4/n25_neg_lutinv ),
    .c(\PWM4/n26 [18]),
    .d(\PWM4/pnumr [18]),
    .o(_al_u2045_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2046 (
    .a(_al_u2045_o),
    .b(\PWM4/n24 ),
    .c(pnumcnt4[18]),
    .d(\PWM4/pnumr [18]),
    .e(pwm_start_stop[20]),
    .o(\PWM4/n31 [18]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2047 (
    .a(\PWM4/n24 ),
    .b(\PWM4/n25_neg_lutinv ),
    .c(\PWM4/n26 [17]),
    .d(\PWM4/pnumr [17]),
    .o(_al_u2047_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2048 (
    .a(_al_u2047_o),
    .b(\PWM4/n24 ),
    .c(pnumcnt4[17]),
    .d(\PWM4/pnumr [17]),
    .e(pwm_start_stop[20]),
    .o(\PWM4/n31 [17]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2049 (
    .a(\PWM4/n24 ),
    .b(\PWM4/n25_neg_lutinv ),
    .c(\PWM4/n26 [16]),
    .d(\PWM4/pnumr [16]),
    .o(_al_u2049_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u205 (
    .a(\PWM0/pnumr [22]),
    .b(pnum0[22]),
    .c(pnum0[32]),
    .d(pwm_start_stop[16]),
    .o(\PWM0/n23 [22]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2050 (
    .a(_al_u2049_o),
    .b(\PWM4/n24 ),
    .c(pnumcnt4[16]),
    .d(\PWM4/pnumr [16]),
    .e(pwm_start_stop[20]),
    .o(\PWM4/n31 [16]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2051 (
    .a(\PWM4/n24 ),
    .b(\PWM4/n25_neg_lutinv ),
    .c(\PWM4/n26 [15]),
    .d(\PWM4/pnumr [15]),
    .o(_al_u2051_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2052 (
    .a(_al_u2051_o),
    .b(\PWM4/n24 ),
    .c(pnumcnt4[15]),
    .d(\PWM4/pnumr [15]),
    .e(pwm_start_stop[20]),
    .o(\PWM4/n31 [15]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2053 (
    .a(\PWM4/n24 ),
    .b(\PWM4/n25_neg_lutinv ),
    .c(\PWM4/n26 [14]),
    .d(\PWM4/pnumr [14]),
    .o(_al_u2053_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2054 (
    .a(_al_u2053_o),
    .b(\PWM4/n24 ),
    .c(pnumcnt4[14]),
    .d(\PWM4/pnumr [14]),
    .e(pwm_start_stop[20]),
    .o(\PWM4/n31 [14]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2055 (
    .a(\PWM4/n24 ),
    .b(\PWM4/n25_neg_lutinv ),
    .c(\PWM4/n26 [13]),
    .d(\PWM4/pnumr [13]),
    .o(_al_u2055_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2056 (
    .a(_al_u2055_o),
    .b(\PWM4/n24 ),
    .c(pnumcnt4[13]),
    .d(\PWM4/pnumr [13]),
    .e(pwm_start_stop[20]),
    .o(\PWM4/n31 [13]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2057 (
    .a(\PWM4/n24 ),
    .b(\PWM4/n25_neg_lutinv ),
    .c(\PWM4/n26 [12]),
    .d(\PWM4/pnumr [12]),
    .o(_al_u2057_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2058 (
    .a(_al_u2057_o),
    .b(\PWM4/n24 ),
    .c(pnumcnt4[12]),
    .d(\PWM4/pnumr [12]),
    .e(pwm_start_stop[20]),
    .o(\PWM4/n31 [12]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2059 (
    .a(\PWM4/n24 ),
    .b(\PWM4/n25_neg_lutinv ),
    .c(\PWM4/n26 [11]),
    .d(\PWM4/pnumr [11]),
    .o(_al_u2059_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u206 (
    .a(\PWM0/pnumr [21]),
    .b(pnum0[21]),
    .c(pnum0[32]),
    .d(pwm_start_stop[16]),
    .o(\PWM0/n23 [21]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2060 (
    .a(_al_u2059_o),
    .b(\PWM4/n24 ),
    .c(pnumcnt4[11]),
    .d(\PWM4/pnumr [11]),
    .e(pwm_start_stop[20]),
    .o(\PWM4/n31 [11]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2061 (
    .a(\PWM4/n24 ),
    .b(\PWM4/n25_neg_lutinv ),
    .c(\PWM4/n26 [10]),
    .d(\PWM4/pnumr [10]),
    .o(_al_u2061_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2062 (
    .a(_al_u2061_o),
    .b(\PWM4/n24 ),
    .c(pnumcnt4[10]),
    .d(\PWM4/pnumr [10]),
    .e(pwm_start_stop[20]),
    .o(\PWM4/n31 [10]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2063 (
    .a(\PWM4/n24 ),
    .b(\PWM4/n25_neg_lutinv ),
    .c(\PWM4/n26 [1]),
    .d(\PWM4/pnumr [1]),
    .o(_al_u2063_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2064 (
    .a(_al_u2063_o),
    .b(\PWM4/n24 ),
    .c(pnumcnt4[1]),
    .d(\PWM4/pnumr [1]),
    .e(pwm_start_stop[20]),
    .o(\PWM4/n31 [1]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2065 (
    .a(\PWM4/n24 ),
    .b(\PWM4/n25_neg_lutinv ),
    .c(\PWM4/n26 [0]),
    .d(\PWM4/pnumr [0]),
    .o(_al_u2065_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2066 (
    .a(_al_u2065_o),
    .b(\PWM4/n24 ),
    .c(pnumcnt4[0]),
    .d(\PWM4/pnumr [0]),
    .e(pwm_start_stop[20]),
    .o(\PWM4/n31 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(~D*A))"),
    .INIT(16'hf351))
    _al_u2067 (
    .a(\PWM4/FreCnt [1]),
    .b(\PWM4/FreCnt [12]),
    .c(\PWM4/FreCntr [13]),
    .d(\PWM4/FreCntr [2]),
    .o(_al_u2067_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*C)*~(~D*B))"),
    .INIT(32'haa220a02))
    _al_u2068 (
    .a(_al_u2067_o),
    .b(\PWM4/FreCnt [25]),
    .c(\PWM4/FreCnt [5]),
    .d(\PWM4/FreCntr [26]),
    .e(\PWM4/FreCntr [6]),
    .o(_al_u2068_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u2069 (
    .a(\PWM4/FreCnt [17]),
    .b(\PWM4/FreCnt [19]),
    .c(\PWM4/FreCntr [18]),
    .d(\PWM4/FreCntr [20]),
    .o(_al_u2069_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u207 (
    .a(\PWM0/pnumr [20]),
    .b(pnum0[20]),
    .c(pnum0[32]),
    .d(pwm_start_stop[16]),
    .o(\PWM0/n23 [20]));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D@C))"),
    .INIT(16'h8008))
    _al_u2070 (
    .a(_al_u2068_o),
    .b(_al_u2069_o),
    .c(\PWM4/FreCnt [16]),
    .d(\PWM4/FreCntr [17]),
    .o(_al_u2070_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u2071 (
    .a(\PWM4/FreCnt [0]),
    .b(\PWM4/FreCnt [8]),
    .c(\PWM4/FreCntr [1]),
    .d(\PWM4/FreCntr [9]),
    .o(_al_u2071_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*~C)*~(D*~B))"),
    .INIT(32'h80a088aa))
    _al_u2072 (
    .a(_al_u2071_o),
    .b(\PWM4/FreCnt [5]),
    .c(\PWM4/FreCnt [7]),
    .d(\PWM4/FreCntr [6]),
    .e(\PWM4/FreCntr [8]),
    .o(_al_u2072_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u2073 (
    .a(\PWM4/FreCnt [15]),
    .b(\PWM4/FreCnt [19]),
    .c(\PWM4/FreCntr [16]),
    .d(\PWM4/FreCntr [20]),
    .o(_al_u2073_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*~C)*~(D*~B))"),
    .INIT(32'h80a088aa))
    _al_u2074 (
    .a(_al_u2073_o),
    .b(\PWM4/FreCnt [12]),
    .c(\PWM4/FreCnt [8]),
    .d(\PWM4/FreCntr [13]),
    .e(\PWM4/FreCntr [9]),
    .o(_al_u2074_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u2075 (
    .a(_al_u2070_o),
    .b(_al_u2072_o),
    .c(_al_u2074_o),
    .o(_al_u2075_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u2076 (
    .a(\PWM4/FreCnt [14]),
    .b(\PWM4/FreCnt [4]),
    .c(\PWM4/FreCntr [15]),
    .d(\PWM4/FreCntr [5]),
    .o(_al_u2076_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u2077 (
    .a(_al_u2076_o),
    .b(\PWM4/FreCnt [20]),
    .c(\PWM4/FreCntr [21]),
    .o(_al_u2077_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u2078 (
    .a(\PWM4/FreCnt [18]),
    .b(\PWM4/FreCnt [2]),
    .c(\PWM4/FreCntr [19]),
    .d(\PWM4/FreCntr [3]),
    .o(_al_u2078_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u2079 (
    .a(_al_u2078_o),
    .b(\PWM4/FreCnt [21]),
    .c(\PWM4/FreCnt [22]),
    .d(\PWM4/FreCntr [22]),
    .e(\PWM4/FreCntr [23]),
    .o(_al_u2079_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u208 (
    .a(\PWM0/pnumr [2]),
    .b(pnum0[2]),
    .c(pnum0[32]),
    .d(pwm_start_stop[16]),
    .o(\PWM0/n23 [2]));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u2080 (
    .a(\PWM4/FreCnt [1]),
    .b(\PWM4/FreCnt [23]),
    .c(\PWM4/FreCntr [2]),
    .d(\PWM4/FreCntr [24]),
    .o(_al_u2080_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*~C)*~(~D*B))"),
    .INIT(32'ha020aa22))
    _al_u2081 (
    .a(_al_u2080_o),
    .b(\PWM4/FreCnt [17]),
    .c(\PWM4/FreCnt [3]),
    .d(\PWM4/FreCntr [18]),
    .e(\PWM4/FreCntr [4]),
    .o(_al_u2081_o));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(E*~B)*~(D@A))"),
    .INIT(32'h08040a05))
    _al_u2082 (
    .a(\PWM4/FreCnt [10]),
    .b(\PWM4/FreCnt [25]),
    .c(\PWM4/FreCnt [26]),
    .d(\PWM4/FreCntr [11]),
    .e(\PWM4/FreCntr [26]),
    .o(_al_u2082_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u2083 (
    .a(_al_u2077_o),
    .b(_al_u2079_o),
    .c(_al_u2081_o),
    .d(_al_u2082_o),
    .o(_al_u2083_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u2084 (
    .a(\PWM4/FreCnt [15]),
    .b(\PWM4/FreCnt [7]),
    .c(\PWM4/FreCntr [16]),
    .d(\PWM4/FreCntr [8]),
    .o(_al_u2084_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*C)*~(D*~B))"),
    .INIT(32'h88aa080a))
    _al_u2085 (
    .a(_al_u2084_o),
    .b(\PWM4/FreCnt [13]),
    .c(\PWM4/FreCnt [3]),
    .d(\PWM4/FreCntr [14]),
    .e(\PWM4/FreCntr [4]),
    .o(_al_u2085_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*~C)*~(D@B))"),
    .INIT(32'h80208822))
    _al_u2086 (
    .a(_al_u2085_o),
    .b(\PWM4/FreCnt [11]),
    .c(\PWM4/FreCnt [23]),
    .d(\PWM4/FreCntr [12]),
    .e(\PWM4/FreCntr [24]),
    .o(_al_u2086_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2087 (
    .a(\PWM4/FreCnt [13]),
    .b(\PWM4/FreCntr [14]),
    .o(_al_u2087_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(~E*C)*~(D@B))"),
    .INIT(32'h44110401))
    _al_u2088 (
    .a(_al_u2087_o),
    .b(\PWM4/FreCnt [24]),
    .c(\PWM4/FreCnt [6]),
    .d(\PWM4/FreCntr [25]),
    .e(\PWM4/FreCntr [7]),
    .o(_al_u2088_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2089 (
    .a(\PWM4/FreCnt [6]),
    .b(\PWM4/FreCntr [7]),
    .o(_al_u2089_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u209 (
    .a(\PWM0/pnumr [19]),
    .b(pnum0[19]),
    .c(pnum0[32]),
    .d(pwm_start_stop[16]),
    .o(\PWM0/n23 [19]));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(E@C)*~(D*~B))"),
    .INIT(32'h40500405))
    _al_u2090 (
    .a(_al_u2089_o),
    .b(\PWM4/FreCnt [0]),
    .c(\PWM4/FreCnt [9]),
    .d(\PWM4/FreCntr [1]),
    .e(\PWM4/FreCntr [10]),
    .o(_al_u2090_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    _al_u2091 (
    .a(_al_u2075_o),
    .b(_al_u2083_o),
    .c(_al_u2086_o),
    .d(_al_u2088_o),
    .e(_al_u2090_o),
    .o(_al_u2091_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2092 (
    .a(_al_u2091_o),
    .b(pwm_state_read[4]),
    .o(\PWM4/u14_sel_is_1_o ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2093 (
    .a(\PWM5/n0_lutinv ),
    .b(pwm_state_read[5]),
    .o(\PWM5/n24 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u2094 (
    .a(pnumcnt5[18]),
    .b(pnumcnt5[19]),
    .c(pnumcnt5[1]),
    .d(pnumcnt5[20]),
    .o(_al_u2094_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u2095 (
    .a(_al_u2094_o),
    .b(pnumcnt5[21]),
    .c(pnumcnt5[22]),
    .d(pnumcnt5[23]),
    .e(pnumcnt5[2]),
    .o(_al_u2095_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u2096 (
    .a(_al_u2095_o),
    .b(pnumcnt5[6]),
    .c(pnumcnt5[7]),
    .d(pnumcnt5[8]),
    .e(pnumcnt5[9]),
    .o(_al_u2096_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u2097 (
    .a(pnumcnt5[10]),
    .b(pnumcnt5[11]),
    .c(pnumcnt5[12]),
    .d(pnumcnt5[13]),
    .o(_al_u2097_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u2098 (
    .a(_al_u2097_o),
    .b(pnumcnt5[14]),
    .c(pnumcnt5[15]),
    .d(pnumcnt5[16]),
    .e(pnumcnt5[17]),
    .o(_al_u2098_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u2099 (
    .a(pnumcnt5[3]),
    .b(pnumcnt5[4]),
    .c(pnumcnt5[5]),
    .o(_al_u2099_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u210 (
    .a(\PWM0/pnumr [18]),
    .b(pnum0[18]),
    .c(pnum0[32]),
    .d(pwm_start_stop[16]),
    .o(\PWM0/n23 [18]));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u2100 (
    .a(_al_u2096_o),
    .b(_al_u2098_o),
    .c(_al_u2099_o),
    .d(pnumcnt5[0]),
    .o(\PWM5/n25_neg_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2101 (
    .a(\PWM5/n24 ),
    .b(\PWM5/n25_neg_lutinv ),
    .c(\PWM5/n26 [9]),
    .d(\PWM5/pnumr [9]),
    .o(_al_u2101_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2102 (
    .a(_al_u2101_o),
    .b(\PWM5/n24 ),
    .c(pnumcnt5[9]),
    .d(\PWM5/pnumr [9]),
    .e(pwm_start_stop[21]),
    .o(\PWM5/n31 [9]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2103 (
    .a(\PWM5/n24 ),
    .b(\PWM5/n25_neg_lutinv ),
    .c(\PWM5/n26 [8]),
    .d(\PWM5/pnumr [8]),
    .o(_al_u2103_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2104 (
    .a(_al_u2103_o),
    .b(\PWM5/n24 ),
    .c(pnumcnt5[8]),
    .d(\PWM5/pnumr [8]),
    .e(pwm_start_stop[21]),
    .o(\PWM5/n31 [8]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2105 (
    .a(\PWM5/n24 ),
    .b(\PWM5/n25_neg_lutinv ),
    .c(\PWM5/n26 [7]),
    .d(\PWM5/pnumr [7]),
    .o(_al_u2105_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2106 (
    .a(_al_u2105_o),
    .b(\PWM5/n24 ),
    .c(pnumcnt5[7]),
    .d(\PWM5/pnumr [7]),
    .e(pwm_start_stop[21]),
    .o(\PWM5/n31 [7]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2107 (
    .a(\PWM5/n24 ),
    .b(\PWM5/n25_neg_lutinv ),
    .c(\PWM5/n26 [6]),
    .d(\PWM5/pnumr [6]),
    .o(_al_u2107_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2108 (
    .a(_al_u2107_o),
    .b(\PWM5/n24 ),
    .c(pnumcnt5[6]),
    .d(\PWM5/pnumr [6]),
    .e(pwm_start_stop[21]),
    .o(\PWM5/n31 [6]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2109 (
    .a(\PWM5/n24 ),
    .b(\PWM5/n25_neg_lutinv ),
    .c(\PWM5/n26 [5]),
    .d(\PWM5/pnumr [5]),
    .o(_al_u2109_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u211 (
    .a(\PWM0/pnumr [17]),
    .b(pnum0[17]),
    .c(pnum0[32]),
    .d(pwm_start_stop[16]),
    .o(\PWM0/n23 [17]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2110 (
    .a(_al_u2109_o),
    .b(\PWM5/n24 ),
    .c(pnumcnt5[5]),
    .d(\PWM5/pnumr [5]),
    .e(pwm_start_stop[21]),
    .o(\PWM5/n31 [5]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2111 (
    .a(\PWM5/n24 ),
    .b(\PWM5/n25_neg_lutinv ),
    .c(\PWM5/n26 [4]),
    .d(\PWM5/pnumr [4]),
    .o(_al_u2111_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2112 (
    .a(_al_u2111_o),
    .b(\PWM5/n24 ),
    .c(pnumcnt5[4]),
    .d(\PWM5/pnumr [4]),
    .e(pwm_start_stop[21]),
    .o(\PWM5/n31 [4]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2113 (
    .a(\PWM5/n24 ),
    .b(\PWM5/n25_neg_lutinv ),
    .c(\PWM5/n26 [3]),
    .d(\PWM5/pnumr [3]),
    .o(_al_u2113_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2114 (
    .a(_al_u2113_o),
    .b(\PWM5/n24 ),
    .c(pnumcnt5[3]),
    .d(\PWM5/pnumr [3]),
    .e(pwm_start_stop[21]),
    .o(\PWM5/n31 [3]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2115 (
    .a(\PWM5/n24 ),
    .b(\PWM5/n25_neg_lutinv ),
    .c(\PWM5/n26 [23]),
    .d(\PWM5/pnumr [23]),
    .o(_al_u2115_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2116 (
    .a(_al_u2115_o),
    .b(\PWM5/n24 ),
    .c(pnumcnt5[23]),
    .d(\PWM5/pnumr [23]),
    .e(pwm_start_stop[21]),
    .o(\PWM5/n31 [23]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2117 (
    .a(\PWM5/n24 ),
    .b(\PWM5/n25_neg_lutinv ),
    .c(\PWM5/n26 [22]),
    .d(\PWM5/pnumr [22]),
    .o(_al_u2117_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2118 (
    .a(_al_u2117_o),
    .b(\PWM5/n24 ),
    .c(pnumcnt5[22]),
    .d(\PWM5/pnumr [22]),
    .e(pwm_start_stop[21]),
    .o(\PWM5/n31 [22]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2119 (
    .a(\PWM5/n24 ),
    .b(\PWM5/n25_neg_lutinv ),
    .c(\PWM5/n26 [21]),
    .d(\PWM5/pnumr [21]),
    .o(_al_u2119_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u212 (
    .a(\PWM0/pnumr [16]),
    .b(pnum0[16]),
    .c(pnum0[32]),
    .d(pwm_start_stop[16]),
    .o(\PWM0/n23 [16]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2120 (
    .a(_al_u2119_o),
    .b(\PWM5/n24 ),
    .c(pnumcnt5[21]),
    .d(\PWM5/pnumr [21]),
    .e(pwm_start_stop[21]),
    .o(\PWM5/n31 [21]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2121 (
    .a(\PWM5/n24 ),
    .b(\PWM5/n25_neg_lutinv ),
    .c(\PWM5/n26 [20]),
    .d(\PWM5/pnumr [20]),
    .o(_al_u2121_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2122 (
    .a(_al_u2121_o),
    .b(\PWM5/n24 ),
    .c(pnumcnt5[20]),
    .d(\PWM5/pnumr [20]),
    .e(pwm_start_stop[21]),
    .o(\PWM5/n31 [20]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2123 (
    .a(\PWM5/n24 ),
    .b(\PWM5/n25_neg_lutinv ),
    .c(\PWM5/n26 [2]),
    .d(\PWM5/pnumr [2]),
    .o(_al_u2123_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2124 (
    .a(_al_u2123_o),
    .b(\PWM5/n24 ),
    .c(pnumcnt5[2]),
    .d(\PWM5/pnumr [2]),
    .e(pwm_start_stop[21]),
    .o(\PWM5/n31 [2]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2125 (
    .a(\PWM5/n24 ),
    .b(\PWM5/n25_neg_lutinv ),
    .c(\PWM5/n26 [19]),
    .d(\PWM5/pnumr [19]),
    .o(_al_u2125_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2126 (
    .a(_al_u2125_o),
    .b(\PWM5/n24 ),
    .c(pnumcnt5[19]),
    .d(\PWM5/pnumr [19]),
    .e(pwm_start_stop[21]),
    .o(\PWM5/n31 [19]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2127 (
    .a(\PWM5/n24 ),
    .b(\PWM5/n25_neg_lutinv ),
    .c(\PWM5/n26 [18]),
    .d(\PWM5/pnumr [18]),
    .o(_al_u2127_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2128 (
    .a(_al_u2127_o),
    .b(\PWM5/n24 ),
    .c(pnumcnt5[18]),
    .d(\PWM5/pnumr [18]),
    .e(pwm_start_stop[21]),
    .o(\PWM5/n31 [18]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2129 (
    .a(\PWM5/n24 ),
    .b(\PWM5/n25_neg_lutinv ),
    .c(\PWM5/n26 [17]),
    .d(\PWM5/pnumr [17]),
    .o(_al_u2129_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u213 (
    .a(\PWM0/pnumr [15]),
    .b(pnum0[15]),
    .c(pnum0[32]),
    .d(pwm_start_stop[16]),
    .o(\PWM0/n23 [15]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2130 (
    .a(_al_u2129_o),
    .b(\PWM5/n24 ),
    .c(pnumcnt5[17]),
    .d(\PWM5/pnumr [17]),
    .e(pwm_start_stop[21]),
    .o(\PWM5/n31 [17]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2131 (
    .a(\PWM5/n24 ),
    .b(\PWM5/n25_neg_lutinv ),
    .c(\PWM5/n26 [16]),
    .d(\PWM5/pnumr [16]),
    .o(_al_u2131_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2132 (
    .a(_al_u2131_o),
    .b(\PWM5/n24 ),
    .c(pnumcnt5[16]),
    .d(\PWM5/pnumr [16]),
    .e(pwm_start_stop[21]),
    .o(\PWM5/n31 [16]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2133 (
    .a(\PWM5/n24 ),
    .b(\PWM5/n25_neg_lutinv ),
    .c(\PWM5/n26 [15]),
    .d(\PWM5/pnumr [15]),
    .o(_al_u2133_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2134 (
    .a(_al_u2133_o),
    .b(\PWM5/n24 ),
    .c(pnumcnt5[15]),
    .d(\PWM5/pnumr [15]),
    .e(pwm_start_stop[21]),
    .o(\PWM5/n31 [15]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2135 (
    .a(\PWM5/n24 ),
    .b(\PWM5/n25_neg_lutinv ),
    .c(\PWM5/n26 [14]),
    .d(\PWM5/pnumr [14]),
    .o(_al_u2135_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2136 (
    .a(_al_u2135_o),
    .b(\PWM5/n24 ),
    .c(pnumcnt5[14]),
    .d(\PWM5/pnumr [14]),
    .e(pwm_start_stop[21]),
    .o(\PWM5/n31 [14]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2137 (
    .a(\PWM5/n24 ),
    .b(\PWM5/n25_neg_lutinv ),
    .c(\PWM5/n26 [13]),
    .d(\PWM5/pnumr [13]),
    .o(_al_u2137_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2138 (
    .a(_al_u2137_o),
    .b(\PWM5/n24 ),
    .c(pnumcnt5[13]),
    .d(\PWM5/pnumr [13]),
    .e(pwm_start_stop[21]),
    .o(\PWM5/n31 [13]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2139 (
    .a(\PWM5/n24 ),
    .b(\PWM5/n25_neg_lutinv ),
    .c(\PWM5/n26 [12]),
    .d(\PWM5/pnumr [12]),
    .o(_al_u2139_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u214 (
    .a(\PWM0/pnumr [14]),
    .b(pnum0[14]),
    .c(pnum0[32]),
    .d(pwm_start_stop[16]),
    .o(\PWM0/n23 [14]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2140 (
    .a(_al_u2139_o),
    .b(\PWM5/n24 ),
    .c(pnumcnt5[12]),
    .d(\PWM5/pnumr [12]),
    .e(pwm_start_stop[21]),
    .o(\PWM5/n31 [12]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2141 (
    .a(\PWM5/n24 ),
    .b(\PWM5/n25_neg_lutinv ),
    .c(\PWM5/n26 [11]),
    .d(\PWM5/pnumr [11]),
    .o(_al_u2141_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2142 (
    .a(_al_u2141_o),
    .b(\PWM5/n24 ),
    .c(pnumcnt5[11]),
    .d(\PWM5/pnumr [11]),
    .e(pwm_start_stop[21]),
    .o(\PWM5/n31 [11]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2143 (
    .a(\PWM5/n24 ),
    .b(\PWM5/n25_neg_lutinv ),
    .c(\PWM5/n26 [10]),
    .d(\PWM5/pnumr [10]),
    .o(_al_u2143_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2144 (
    .a(_al_u2143_o),
    .b(\PWM5/n24 ),
    .c(pnumcnt5[10]),
    .d(\PWM5/pnumr [10]),
    .e(pwm_start_stop[21]),
    .o(\PWM5/n31 [10]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2145 (
    .a(\PWM5/n24 ),
    .b(\PWM5/n25_neg_lutinv ),
    .c(\PWM5/n26 [1]),
    .d(\PWM5/pnumr [1]),
    .o(_al_u2145_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2146 (
    .a(_al_u2145_o),
    .b(\PWM5/n24 ),
    .c(pnumcnt5[1]),
    .d(\PWM5/pnumr [1]),
    .e(pwm_start_stop[21]),
    .o(\PWM5/n31 [1]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2147 (
    .a(\PWM5/n24 ),
    .b(\PWM5/n25_neg_lutinv ),
    .c(\PWM5/n26 [0]),
    .d(\PWM5/pnumr [0]),
    .o(_al_u2147_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2148 (
    .a(_al_u2147_o),
    .b(\PWM5/n24 ),
    .c(pnumcnt5[0]),
    .d(\PWM5/pnumr [0]),
    .e(pwm_start_stop[21]),
    .o(\PWM5/n31 [0]));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(~D*B)*~(E@A))"),
    .INIT(32'h0a020501))
    _al_u2149 (
    .a(\PWM5/FreCnt [2]),
    .b(\PWM5/FreCnt [22]),
    .c(\PWM5/FreCnt [26]),
    .d(\PWM5/FreCntr [23]),
    .e(\PWM5/FreCntr [3]),
    .o(_al_u2149_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u215 (
    .a(\PWM0/pnumr [13]),
    .b(pnum0[13]),
    .c(pnum0[32]),
    .d(pwm_start_stop[16]),
    .o(\PWM0/n23 [13]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u2150 (
    .a(_al_u2149_o),
    .b(\PWM5/FreCnt [24]),
    .c(\PWM5/FreCnt [4]),
    .d(\PWM5/FreCntr [25]),
    .e(\PWM5/FreCntr [5]),
    .o(_al_u2150_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u2151 (
    .a(\PWM5/FreCnt [11]),
    .b(\PWM5/FreCnt [6]),
    .c(\PWM5/FreCntr [12]),
    .d(\PWM5/FreCntr [7]),
    .o(_al_u2151_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u2152 (
    .a(_al_u2151_o),
    .b(\PWM5/FreCnt [0]),
    .c(\PWM5/FreCntr [1]),
    .o(_al_u2152_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u2153 (
    .a(\PWM5/FreCnt [7]),
    .b(\PWM5/FreCnt [8]),
    .c(\PWM5/FreCntr [8]),
    .d(\PWM5/FreCntr [9]),
    .o(_al_u2153_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*C)*~(~D*B))"),
    .INIT(32'haa220a02))
    _al_u2154 (
    .a(_al_u2153_o),
    .b(\PWM5/FreCnt [17]),
    .c(\PWM5/FreCnt [21]),
    .d(\PWM5/FreCntr [18]),
    .e(\PWM5/FreCntr [22]),
    .o(_al_u2154_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2155 (
    .a(\PWM5/FreCnt [19]),
    .b(\PWM5/FreCntr [20]),
    .o(_al_u2155_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(E*~C)*~(D@B))"),
    .INIT(32'h40104411))
    _al_u2156 (
    .a(_al_u2155_o),
    .b(\PWM5/FreCnt [14]),
    .c(\PWM5/FreCnt [22]),
    .d(\PWM5/FreCntr [15]),
    .e(\PWM5/FreCntr [23]),
    .o(_al_u2156_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u2157 (
    .a(_al_u2150_o),
    .b(_al_u2152_o),
    .c(_al_u2154_o),
    .d(_al_u2156_o),
    .o(_al_u2157_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u2158 (
    .a(\PWM5/FreCnt [12]),
    .b(\PWM5/FreCnt [21]),
    .c(\PWM5/FreCntr [13]),
    .d(\PWM5/FreCntr [22]),
    .o(_al_u2158_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~D*C)*~(E*~B))"),
    .INIT(32'h8808aa0a))
    _al_u2159 (
    .a(_al_u2158_o),
    .b(\PWM5/FreCnt [1]),
    .c(\PWM5/FreCnt [15]),
    .d(\PWM5/FreCntr [16]),
    .e(\PWM5/FreCntr [2]),
    .o(_al_u2159_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u216 (
    .a(\PWM0/pnumr [12]),
    .b(pnum0[12]),
    .c(pnum0[32]),
    .d(pwm_start_stop[16]),
    .o(\PWM0/n23 [12]));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u2160 (
    .a(\PWM5/FreCnt [5]),
    .b(\PWM5/FreCnt [7]),
    .c(\PWM5/FreCntr [6]),
    .d(\PWM5/FreCntr [8]),
    .o(_al_u2160_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*C)*~(~D*B))"),
    .INIT(32'haa220a02))
    _al_u2161 (
    .a(_al_u2160_o),
    .b(\PWM5/FreCnt [13]),
    .c(\PWM5/FreCnt [23]),
    .d(\PWM5/FreCntr [14]),
    .e(\PWM5/FreCntr [24]),
    .o(_al_u2161_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u2162 (
    .a(\PWM5/FreCnt [16]),
    .b(\PWM5/FreCnt [18]),
    .c(\PWM5/FreCntr [17]),
    .d(\PWM5/FreCntr [19]),
    .o(_al_u2162_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D@C)*~(E@B))"),
    .INIT(32'h80082002))
    _al_u2163 (
    .a(_al_u2162_o),
    .b(\PWM5/FreCnt [20]),
    .c(\PWM5/FreCnt [9]),
    .d(\PWM5/FreCntr [10]),
    .e(\PWM5/FreCntr [21]),
    .o(_al_u2163_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u2164 (
    .a(_al_u2159_o),
    .b(_al_u2161_o),
    .c(_al_u2163_o),
    .o(_al_u2164_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u2165 (
    .a(\PWM5/FreCnt [10]),
    .b(\PWM5/FreCnt [12]),
    .c(\PWM5/FreCntr [11]),
    .d(\PWM5/FreCntr [13]),
    .o(_al_u2165_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*C)*~(D*~B))"),
    .INIT(32'h88aa080a))
    _al_u2166 (
    .a(_al_u2165_o),
    .b(\PWM5/FreCnt [25]),
    .c(\PWM5/FreCnt [3]),
    .d(\PWM5/FreCntr [26]),
    .e(\PWM5/FreCntr [4]),
    .o(_al_u2166_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u2167 (
    .a(\PWM5/FreCnt [10]),
    .b(\PWM5/FreCnt [5]),
    .c(\PWM5/FreCntr [11]),
    .d(\PWM5/FreCntr [6]),
    .o(_al_u2167_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(~D*C))"),
    .INIT(16'h8808))
    _al_u2168 (
    .a(_al_u2166_o),
    .b(_al_u2167_o),
    .c(\PWM5/FreCnt [8]),
    .d(\PWM5/FreCntr [9]),
    .o(_al_u2168_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u2169 (
    .a(\PWM5/FreCnt [15]),
    .b(\PWM5/FreCnt [19]),
    .c(\PWM5/FreCntr [16]),
    .d(\PWM5/FreCntr [20]),
    .o(_al_u2169_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u217 (
    .a(\PWM0/pnumr [11]),
    .b(pnum0[11]),
    .c(pnum0[32]),
    .d(pwm_start_stop[16]),
    .o(\PWM0/n23 [11]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*~C)*~(~D*B))"),
    .INIT(32'ha020aa22))
    _al_u2170 (
    .a(_al_u2169_o),
    .b(\PWM5/FreCnt [25]),
    .c(\PWM5/FreCnt [3]),
    .d(\PWM5/FreCntr [26]),
    .e(\PWM5/FreCntr [4]),
    .o(_al_u2170_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u2171 (
    .a(\PWM5/FreCnt [1]),
    .b(\PWM5/FreCnt [23]),
    .c(\PWM5/FreCntr [2]),
    .d(\PWM5/FreCntr [24]),
    .o(_al_u2171_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*~C)*~(D*~B))"),
    .INIT(32'h80a088aa))
    _al_u2172 (
    .a(_al_u2171_o),
    .b(\PWM5/FreCnt [13]),
    .c(\PWM5/FreCnt [17]),
    .d(\PWM5/FreCntr [14]),
    .e(\PWM5/FreCntr [18]),
    .o(_al_u2172_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    _al_u2173 (
    .a(_al_u2157_o),
    .b(_al_u2164_o),
    .c(_al_u2168_o),
    .d(_al_u2170_o),
    .e(_al_u2172_o),
    .o(_al_u2173_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2174 (
    .a(_al_u2173_o),
    .b(pwm_state_read[5]),
    .o(\PWM5/u14_sel_is_1_o ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2175 (
    .a(\PWM6/n0_lutinv ),
    .b(pwm_state_read[6]),
    .o(\PWM6/n24 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u2176 (
    .a(pnumcnt6[18]),
    .b(pnumcnt6[19]),
    .c(pnumcnt6[1]),
    .d(pnumcnt6[20]),
    .o(_al_u2176_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u2177 (
    .a(_al_u2176_o),
    .b(pnumcnt6[21]),
    .c(pnumcnt6[22]),
    .d(pnumcnt6[23]),
    .e(pnumcnt6[2]),
    .o(_al_u2177_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u2178 (
    .a(_al_u2177_o),
    .b(pnumcnt6[6]),
    .c(pnumcnt6[7]),
    .d(pnumcnt6[8]),
    .e(pnumcnt6[9]),
    .o(_al_u2178_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u2179 (
    .a(pnumcnt6[10]),
    .b(pnumcnt6[11]),
    .c(pnumcnt6[12]),
    .d(pnumcnt6[13]),
    .o(_al_u2179_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u218 (
    .a(\PWM0/pnumr [10]),
    .b(pnum0[10]),
    .c(pnum0[32]),
    .d(pwm_start_stop[16]),
    .o(\PWM0/n23 [10]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u2180 (
    .a(_al_u2179_o),
    .b(pnumcnt6[14]),
    .c(pnumcnt6[15]),
    .d(pnumcnt6[16]),
    .e(pnumcnt6[17]),
    .o(_al_u2180_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u2181 (
    .a(pnumcnt6[3]),
    .b(pnumcnt6[4]),
    .c(pnumcnt6[5]),
    .o(_al_u2181_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u2182 (
    .a(_al_u2178_o),
    .b(_al_u2180_o),
    .c(_al_u2181_o),
    .d(pnumcnt6[0]),
    .o(\PWM6/n25_neg_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2183 (
    .a(\PWM6/n24 ),
    .b(\PWM6/n25_neg_lutinv ),
    .c(\PWM6/n26 [9]),
    .d(\PWM6/pnumr [9]),
    .o(_al_u2183_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2184 (
    .a(_al_u2183_o),
    .b(\PWM6/n24 ),
    .c(pnumcnt6[9]),
    .d(\PWM6/pnumr [9]),
    .e(pwm_start_stop[22]),
    .o(\PWM6/n31 [9]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2185 (
    .a(\PWM6/n24 ),
    .b(\PWM6/n25_neg_lutinv ),
    .c(\PWM6/n26 [8]),
    .d(\PWM6/pnumr [8]),
    .o(_al_u2185_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2186 (
    .a(_al_u2185_o),
    .b(\PWM6/n24 ),
    .c(pnumcnt6[8]),
    .d(\PWM6/pnumr [8]),
    .e(pwm_start_stop[22]),
    .o(\PWM6/n31 [8]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2187 (
    .a(\PWM6/n24 ),
    .b(\PWM6/n25_neg_lutinv ),
    .c(\PWM6/n26 [7]),
    .d(\PWM6/pnumr [7]),
    .o(_al_u2187_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2188 (
    .a(_al_u2187_o),
    .b(\PWM6/n24 ),
    .c(pnumcnt6[7]),
    .d(\PWM6/pnumr [7]),
    .e(pwm_start_stop[22]),
    .o(\PWM6/n31 [7]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2189 (
    .a(\PWM6/n24 ),
    .b(\PWM6/n25_neg_lutinv ),
    .c(\PWM6/n26 [6]),
    .d(\PWM6/pnumr [6]),
    .o(_al_u2189_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u219 (
    .a(\PWM0/pnumr [1]),
    .b(pnum0[1]),
    .c(pnum0[32]),
    .d(pwm_start_stop[16]),
    .o(\PWM0/n23 [1]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2190 (
    .a(_al_u2189_o),
    .b(\PWM6/n24 ),
    .c(pnumcnt6[6]),
    .d(\PWM6/pnumr [6]),
    .e(pwm_start_stop[22]),
    .o(\PWM6/n31 [6]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2191 (
    .a(\PWM6/n24 ),
    .b(\PWM6/n25_neg_lutinv ),
    .c(\PWM6/n26 [5]),
    .d(\PWM6/pnumr [5]),
    .o(_al_u2191_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2192 (
    .a(_al_u2191_o),
    .b(\PWM6/n24 ),
    .c(pnumcnt6[5]),
    .d(\PWM6/pnumr [5]),
    .e(pwm_start_stop[22]),
    .o(\PWM6/n31 [5]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2193 (
    .a(\PWM6/n24 ),
    .b(\PWM6/n25_neg_lutinv ),
    .c(\PWM6/n26 [4]),
    .d(\PWM6/pnumr [4]),
    .o(_al_u2193_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2194 (
    .a(_al_u2193_o),
    .b(\PWM6/n24 ),
    .c(pnumcnt6[4]),
    .d(\PWM6/pnumr [4]),
    .e(pwm_start_stop[22]),
    .o(\PWM6/n31 [4]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2195 (
    .a(\PWM6/n24 ),
    .b(\PWM6/n25_neg_lutinv ),
    .c(\PWM6/n26 [3]),
    .d(\PWM6/pnumr [3]),
    .o(_al_u2195_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2196 (
    .a(_al_u2195_o),
    .b(\PWM6/n24 ),
    .c(pnumcnt6[3]),
    .d(\PWM6/pnumr [3]),
    .e(pwm_start_stop[22]),
    .o(\PWM6/n31 [3]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2197 (
    .a(\PWM6/n24 ),
    .b(\PWM6/n25_neg_lutinv ),
    .c(\PWM6/n26 [23]),
    .d(\PWM6/pnumr [23]),
    .o(_al_u2197_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2198 (
    .a(_al_u2197_o),
    .b(\PWM6/n24 ),
    .c(pnumcnt6[23]),
    .d(\PWM6/pnumr [23]),
    .e(pwm_start_stop[22]),
    .o(\PWM6/n31 [23]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2199 (
    .a(\PWM6/n24 ),
    .b(\PWM6/n25_neg_lutinv ),
    .c(\PWM6/n26 [22]),
    .d(\PWM6/pnumr [22]),
    .o(_al_u2199_o));
  EF2_PHY_SPAD #(
    //.LOCATION("P28"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u22 (
    .ipad(clkin),
    .ts(1'b1),
    .di(clkin_pad));  // CPLD_SOC_AHB_TOP.v(3)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u220 (
    .a(\PWM0/pnumr [0]),
    .b(pnum0[0]),
    .c(pnum0[32]),
    .d(pwm_start_stop[16]),
    .o(\PWM0/n23 [0]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2200 (
    .a(_al_u2199_o),
    .b(\PWM6/n24 ),
    .c(pnumcnt6[22]),
    .d(\PWM6/pnumr [22]),
    .e(pwm_start_stop[22]),
    .o(\PWM6/n31 [22]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2201 (
    .a(\PWM6/n24 ),
    .b(\PWM6/n25_neg_lutinv ),
    .c(\PWM6/n26 [21]),
    .d(\PWM6/pnumr [21]),
    .o(_al_u2201_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2202 (
    .a(_al_u2201_o),
    .b(\PWM6/n24 ),
    .c(pnumcnt6[21]),
    .d(\PWM6/pnumr [21]),
    .e(pwm_start_stop[22]),
    .o(\PWM6/n31 [21]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2203 (
    .a(\PWM6/n24 ),
    .b(\PWM6/n25_neg_lutinv ),
    .c(\PWM6/n26 [20]),
    .d(\PWM6/pnumr [20]),
    .o(_al_u2203_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2204 (
    .a(_al_u2203_o),
    .b(\PWM6/n24 ),
    .c(pnumcnt6[20]),
    .d(\PWM6/pnumr [20]),
    .e(pwm_start_stop[22]),
    .o(\PWM6/n31 [20]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2205 (
    .a(\PWM6/n24 ),
    .b(\PWM6/n25_neg_lutinv ),
    .c(\PWM6/n26 [2]),
    .d(\PWM6/pnumr [2]),
    .o(_al_u2205_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2206 (
    .a(_al_u2205_o),
    .b(\PWM6/n24 ),
    .c(pnumcnt6[2]),
    .d(\PWM6/pnumr [2]),
    .e(pwm_start_stop[22]),
    .o(\PWM6/n31 [2]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2207 (
    .a(\PWM6/n24 ),
    .b(\PWM6/n25_neg_lutinv ),
    .c(\PWM6/n26 [19]),
    .d(\PWM6/pnumr [19]),
    .o(_al_u2207_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2208 (
    .a(_al_u2207_o),
    .b(\PWM6/n24 ),
    .c(pnumcnt6[19]),
    .d(\PWM6/pnumr [19]),
    .e(pwm_start_stop[22]),
    .o(\PWM6/n31 [19]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2209 (
    .a(\PWM6/n24 ),
    .b(\PWM6/n25_neg_lutinv ),
    .c(\PWM6/n26 [18]),
    .d(\PWM6/pnumr [18]),
    .o(_al_u2209_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u221 (
    .a(\PWM1/pnumr [9]),
    .b(pnum1[32]),
    .c(pnum1[9]),
    .d(pwm_start_stop[17]),
    .o(\PWM1/n23 [9]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2210 (
    .a(_al_u2209_o),
    .b(\PWM6/n24 ),
    .c(pnumcnt6[18]),
    .d(\PWM6/pnumr [18]),
    .e(pwm_start_stop[22]),
    .o(\PWM6/n31 [18]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2211 (
    .a(\PWM6/n24 ),
    .b(\PWM6/n25_neg_lutinv ),
    .c(\PWM6/n26 [17]),
    .d(\PWM6/pnumr [17]),
    .o(_al_u2211_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2212 (
    .a(_al_u2211_o),
    .b(\PWM6/n24 ),
    .c(pnumcnt6[17]),
    .d(\PWM6/pnumr [17]),
    .e(pwm_start_stop[22]),
    .o(\PWM6/n31 [17]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2213 (
    .a(\PWM6/n24 ),
    .b(\PWM6/n25_neg_lutinv ),
    .c(\PWM6/n26 [16]),
    .d(\PWM6/pnumr [16]),
    .o(_al_u2213_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2214 (
    .a(_al_u2213_o),
    .b(\PWM6/n24 ),
    .c(pnumcnt6[16]),
    .d(\PWM6/pnumr [16]),
    .e(pwm_start_stop[22]),
    .o(\PWM6/n31 [16]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2215 (
    .a(\PWM6/n24 ),
    .b(\PWM6/n25_neg_lutinv ),
    .c(\PWM6/n26 [15]),
    .d(\PWM6/pnumr [15]),
    .o(_al_u2215_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2216 (
    .a(_al_u2215_o),
    .b(\PWM6/n24 ),
    .c(pnumcnt6[15]),
    .d(\PWM6/pnumr [15]),
    .e(pwm_start_stop[22]),
    .o(\PWM6/n31 [15]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2217 (
    .a(\PWM6/n24 ),
    .b(\PWM6/n25_neg_lutinv ),
    .c(\PWM6/n26 [14]),
    .d(\PWM6/pnumr [14]),
    .o(_al_u2217_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2218 (
    .a(_al_u2217_o),
    .b(\PWM6/n24 ),
    .c(pnumcnt6[14]),
    .d(\PWM6/pnumr [14]),
    .e(pwm_start_stop[22]),
    .o(\PWM6/n31 [14]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2219 (
    .a(\PWM6/n24 ),
    .b(\PWM6/n25_neg_lutinv ),
    .c(\PWM6/n26 [13]),
    .d(\PWM6/pnumr [13]),
    .o(_al_u2219_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u222 (
    .a(\PWM1/pnumr [8]),
    .b(pnum1[32]),
    .c(pnum1[8]),
    .d(pwm_start_stop[17]),
    .o(\PWM1/n23 [8]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2220 (
    .a(_al_u2219_o),
    .b(\PWM6/n24 ),
    .c(pnumcnt6[13]),
    .d(\PWM6/pnumr [13]),
    .e(pwm_start_stop[22]),
    .o(\PWM6/n31 [13]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2221 (
    .a(\PWM6/n24 ),
    .b(\PWM6/n25_neg_lutinv ),
    .c(\PWM6/n26 [12]),
    .d(\PWM6/pnumr [12]),
    .o(_al_u2221_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2222 (
    .a(_al_u2221_o),
    .b(\PWM6/n24 ),
    .c(pnumcnt6[12]),
    .d(\PWM6/pnumr [12]),
    .e(pwm_start_stop[22]),
    .o(\PWM6/n31 [12]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2223 (
    .a(\PWM6/n24 ),
    .b(\PWM6/n25_neg_lutinv ),
    .c(\PWM6/n26 [11]),
    .d(\PWM6/pnumr [11]),
    .o(_al_u2223_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2224 (
    .a(_al_u2223_o),
    .b(\PWM6/n24 ),
    .c(pnumcnt6[11]),
    .d(\PWM6/pnumr [11]),
    .e(pwm_start_stop[22]),
    .o(\PWM6/n31 [11]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2225 (
    .a(\PWM6/n24 ),
    .b(\PWM6/n25_neg_lutinv ),
    .c(\PWM6/n26 [10]),
    .d(\PWM6/pnumr [10]),
    .o(_al_u2225_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2226 (
    .a(_al_u2225_o),
    .b(\PWM6/n24 ),
    .c(pnumcnt6[10]),
    .d(\PWM6/pnumr [10]),
    .e(pwm_start_stop[22]),
    .o(\PWM6/n31 [10]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2227 (
    .a(\PWM6/n24 ),
    .b(\PWM6/n25_neg_lutinv ),
    .c(\PWM6/n26 [1]),
    .d(\PWM6/pnumr [1]),
    .o(_al_u2227_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2228 (
    .a(_al_u2227_o),
    .b(\PWM6/n24 ),
    .c(pnumcnt6[1]),
    .d(\PWM6/pnumr [1]),
    .e(pwm_start_stop[22]),
    .o(\PWM6/n31 [1]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2229 (
    .a(\PWM6/n24 ),
    .b(\PWM6/n25_neg_lutinv ),
    .c(\PWM6/n26 [0]),
    .d(\PWM6/pnumr [0]),
    .o(_al_u2229_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u223 (
    .a(\PWM1/pnumr [7]),
    .b(pnum1[32]),
    .c(pnum1[7]),
    .d(pwm_start_stop[17]),
    .o(\PWM1/n23 [7]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2230 (
    .a(_al_u2229_o),
    .b(\PWM6/n24 ),
    .c(pnumcnt6[0]),
    .d(\PWM6/pnumr [0]),
    .e(pwm_start_stop[22]),
    .o(\PWM6/n31 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u2231 (
    .a(\PWM6/FreCnt [10]),
    .b(\PWM6/FreCnt [19]),
    .c(\PWM6/FreCntr [11]),
    .d(\PWM6/FreCntr [20]),
    .o(_al_u2231_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*~C)*~(D*~B))"),
    .INIT(32'h80a088aa))
    _al_u2232 (
    .a(_al_u2231_o),
    .b(\PWM6/FreCnt [17]),
    .c(\PWM6/FreCnt [25]),
    .d(\PWM6/FreCntr [18]),
    .e(\PWM6/FreCntr [26]),
    .o(_al_u2232_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u2233 (
    .a(\PWM6/FreCnt [21]),
    .b(\PWM6/FreCnt [5]),
    .c(\PWM6/FreCntr [22]),
    .d(\PWM6/FreCntr [6]),
    .o(_al_u2233_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(~D*C))"),
    .INIT(16'h8808))
    _al_u2234 (
    .a(_al_u2232_o),
    .b(_al_u2233_o),
    .c(\PWM6/FreCnt [8]),
    .d(\PWM6/FreCntr [9]),
    .o(_al_u2234_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u2235 (
    .a(\PWM6/FreCnt [3]),
    .b(\PWM6/FreCnt [7]),
    .c(\PWM6/FreCntr [4]),
    .d(\PWM6/FreCntr [8]),
    .o(_al_u2235_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*C)*~(D*~B))"),
    .INIT(32'h88aa080a))
    _al_u2236 (
    .a(_al_u2235_o),
    .b(\PWM6/FreCnt [10]),
    .c(\PWM6/FreCnt [25]),
    .d(\PWM6/FreCntr [11]),
    .e(\PWM6/FreCntr [26]),
    .o(_al_u2236_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u2237 (
    .a(\PWM6/FreCnt [1]),
    .b(\PWM6/FreCnt [5]),
    .c(\PWM6/FreCntr [2]),
    .d(\PWM6/FreCntr [6]),
    .o(_al_u2237_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u2238 (
    .a(_al_u2234_o),
    .b(_al_u2236_o),
    .c(_al_u2237_o),
    .d(\PWM6/FreCnt [16]),
    .e(\PWM6/FreCntr [17]),
    .o(_al_u2238_o));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(~D*B)*~(E@A))"),
    .INIT(32'h0a020501))
    _al_u2239 (
    .a(\PWM6/FreCnt [2]),
    .b(\PWM6/FreCnt [22]),
    .c(\PWM6/FreCnt [26]),
    .d(\PWM6/FreCntr [23]),
    .e(\PWM6/FreCntr [3]),
    .o(_al_u2239_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u224 (
    .a(\PWM1/pnumr [6]),
    .b(pnum1[32]),
    .c(pnum1[6]),
    .d(pwm_start_stop[17]),
    .o(\PWM1/n23 [6]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u2240 (
    .a(_al_u2239_o),
    .b(\PWM6/FreCnt [24]),
    .c(\PWM6/FreCnt [6]),
    .d(\PWM6/FreCntr [25]),
    .e(\PWM6/FreCntr [7]),
    .o(_al_u2240_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u2241 (
    .a(\PWM6/FreCnt [0]),
    .b(\PWM6/FreCnt [18]),
    .c(\PWM6/FreCntr [1]),
    .d(\PWM6/FreCntr [19]),
    .o(_al_u2241_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u2242 (
    .a(_al_u2241_o),
    .b(\PWM6/FreCnt [4]),
    .c(\PWM6/FreCntr [5]),
    .o(_al_u2242_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u2243 (
    .a(\PWM6/FreCnt [7]),
    .b(\PWM6/FreCnt [8]),
    .c(\PWM6/FreCntr [8]),
    .d(\PWM6/FreCntr [9]),
    .o(_al_u2243_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*C)*~(~D*B))"),
    .INIT(32'haa220a02))
    _al_u2244 (
    .a(_al_u2243_o),
    .b(\PWM6/FreCnt [17]),
    .c(\PWM6/FreCnt [3]),
    .d(\PWM6/FreCntr [18]),
    .e(\PWM6/FreCntr [4]),
    .o(_al_u2244_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2245 (
    .a(\PWM6/FreCnt [19]),
    .b(\PWM6/FreCntr [20]),
    .o(_al_u2245_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(E*~C)*~(D@B))"),
    .INIT(32'h40104411))
    _al_u2246 (
    .a(_al_u2245_o),
    .b(\PWM6/FreCnt [11]),
    .c(\PWM6/FreCnt [22]),
    .d(\PWM6/FreCntr [12]),
    .e(\PWM6/FreCntr [23]),
    .o(_al_u2246_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u2247 (
    .a(_al_u2240_o),
    .b(_al_u2242_o),
    .c(_al_u2244_o),
    .d(_al_u2246_o),
    .o(_al_u2247_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u2248 (
    .a(\PWM6/FreCnt [13]),
    .b(\PWM6/FreCnt [14]),
    .c(\PWM6/FreCntr [14]),
    .d(\PWM6/FreCntr [15]),
    .o(_al_u2248_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D@C)*~(E@B))"),
    .INIT(32'h80082002))
    _al_u2249 (
    .a(_al_u2248_o),
    .b(\PWM6/FreCnt [20]),
    .c(\PWM6/FreCnt [9]),
    .d(\PWM6/FreCntr [10]),
    .e(\PWM6/FreCntr [21]),
    .o(_al_u2249_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u225 (
    .a(\PWM1/pnumr [5]),
    .b(pnum1[32]),
    .c(pnum1[5]),
    .d(pwm_start_stop[17]),
    .o(\PWM1/n23 [5]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2250 (
    .a(\PWM6/FreCnt [15]),
    .b(\PWM6/FreCntr [16]),
    .o(_al_u2250_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(E@C)*~(~D*B))"),
    .INIT(32'h50100501))
    _al_u2251 (
    .a(_al_u2250_o),
    .b(\PWM6/FreCnt [1]),
    .c(\PWM6/FreCnt [23]),
    .d(\PWM6/FreCntr [2]),
    .e(\PWM6/FreCntr [24]),
    .o(_al_u2251_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u2252 (
    .a(\PWM6/FreCnt [15]),
    .b(\PWM6/FreCnt [21]),
    .c(\PWM6/FreCntr [16]),
    .d(\PWM6/FreCntr [22]),
    .o(_al_u2252_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u2253 (
    .a(_al_u2249_o),
    .b(_al_u2251_o),
    .c(_al_u2252_o),
    .d(\PWM6/FreCnt [12]),
    .e(\PWM6/FreCntr [13]),
    .o(_al_u2253_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*A))"),
    .INIT(16'h7f00))
    _al_u2254 (
    .a(_al_u2238_o),
    .b(_al_u2247_o),
    .c(_al_u2253_o),
    .d(pwm_state_read[6]),
    .o(\PWM6/u14_sel_is_1_o ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2255 (
    .a(\PWM7/n0_lutinv ),
    .b(pwm_state_read[7]),
    .o(\PWM7/n24 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u2256 (
    .a(pnumcnt7[18]),
    .b(pnumcnt7[19]),
    .c(pnumcnt7[1]),
    .d(pnumcnt7[20]),
    .o(_al_u2256_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u2257 (
    .a(_al_u2256_o),
    .b(pnumcnt7[21]),
    .c(pnumcnt7[22]),
    .d(pnumcnt7[23]),
    .e(pnumcnt7[2]),
    .o(_al_u2257_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u2258 (
    .a(_al_u2257_o),
    .b(pnumcnt7[6]),
    .c(pnumcnt7[7]),
    .d(pnumcnt7[8]),
    .e(pnumcnt7[9]),
    .o(_al_u2258_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u2259 (
    .a(pnumcnt7[10]),
    .b(pnumcnt7[11]),
    .c(pnumcnt7[12]),
    .d(pnumcnt7[13]),
    .o(_al_u2259_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u226 (
    .a(\PWM1/pnumr [4]),
    .b(pnum1[32]),
    .c(pnum1[4]),
    .d(pwm_start_stop[17]),
    .o(\PWM1/n23 [4]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u2260 (
    .a(_al_u2259_o),
    .b(pnumcnt7[14]),
    .c(pnumcnt7[15]),
    .d(pnumcnt7[16]),
    .e(pnumcnt7[17]),
    .o(_al_u2260_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u2261 (
    .a(pnumcnt7[3]),
    .b(pnumcnt7[4]),
    .c(pnumcnt7[5]),
    .o(_al_u2261_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u2262 (
    .a(_al_u2258_o),
    .b(_al_u2260_o),
    .c(_al_u2261_o),
    .d(pnumcnt7[0]),
    .o(\PWM7/n25_neg_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2263 (
    .a(\PWM7/n24 ),
    .b(\PWM7/n25_neg_lutinv ),
    .c(\PWM7/n26 [9]),
    .d(\PWM7/pnumr [9]),
    .o(_al_u2263_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2264 (
    .a(_al_u2263_o),
    .b(\PWM7/n24 ),
    .c(pnumcnt7[9]),
    .d(\PWM7/pnumr [9]),
    .e(pwm_start_stop[23]),
    .o(\PWM7/n31 [9]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2265 (
    .a(\PWM7/n24 ),
    .b(\PWM7/n25_neg_lutinv ),
    .c(\PWM7/n26 [8]),
    .d(\PWM7/pnumr [8]),
    .o(_al_u2265_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2266 (
    .a(_al_u2265_o),
    .b(\PWM7/n24 ),
    .c(pnumcnt7[8]),
    .d(\PWM7/pnumr [8]),
    .e(pwm_start_stop[23]),
    .o(\PWM7/n31 [8]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2267 (
    .a(\PWM7/n24 ),
    .b(\PWM7/n25_neg_lutinv ),
    .c(\PWM7/n26 [7]),
    .d(\PWM7/pnumr [7]),
    .o(_al_u2267_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2268 (
    .a(_al_u2267_o),
    .b(\PWM7/n24 ),
    .c(pnumcnt7[7]),
    .d(\PWM7/pnumr [7]),
    .e(pwm_start_stop[23]),
    .o(\PWM7/n31 [7]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2269 (
    .a(\PWM7/n24 ),
    .b(\PWM7/n25_neg_lutinv ),
    .c(\PWM7/n26 [6]),
    .d(\PWM7/pnumr [6]),
    .o(_al_u2269_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u227 (
    .a(\PWM1/pnumr [31]),
    .b(pnum1[31]),
    .c(pnum1[32]),
    .d(pwm_start_stop[17]),
    .o(\PWM1/n23 [31]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2270 (
    .a(_al_u2269_o),
    .b(\PWM7/n24 ),
    .c(pnumcnt7[6]),
    .d(\PWM7/pnumr [6]),
    .e(pwm_start_stop[23]),
    .o(\PWM7/n31 [6]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2271 (
    .a(\PWM7/n24 ),
    .b(\PWM7/n25_neg_lutinv ),
    .c(\PWM7/n26 [5]),
    .d(\PWM7/pnumr [5]),
    .o(_al_u2271_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2272 (
    .a(_al_u2271_o),
    .b(\PWM7/n24 ),
    .c(pnumcnt7[5]),
    .d(\PWM7/pnumr [5]),
    .e(pwm_start_stop[23]),
    .o(\PWM7/n31 [5]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2273 (
    .a(\PWM7/n24 ),
    .b(\PWM7/n25_neg_lutinv ),
    .c(\PWM7/n26 [4]),
    .d(\PWM7/pnumr [4]),
    .o(_al_u2273_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2274 (
    .a(_al_u2273_o),
    .b(\PWM7/n24 ),
    .c(pnumcnt7[4]),
    .d(\PWM7/pnumr [4]),
    .e(pwm_start_stop[23]),
    .o(\PWM7/n31 [4]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2275 (
    .a(\PWM7/n24 ),
    .b(\PWM7/n25_neg_lutinv ),
    .c(\PWM7/n26 [3]),
    .d(\PWM7/pnumr [3]),
    .o(_al_u2275_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2276 (
    .a(_al_u2275_o),
    .b(\PWM7/n24 ),
    .c(pnumcnt7[3]),
    .d(\PWM7/pnumr [3]),
    .e(pwm_start_stop[23]),
    .o(\PWM7/n31 [3]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2277 (
    .a(\PWM7/n24 ),
    .b(\PWM7/n25_neg_lutinv ),
    .c(\PWM7/n26 [23]),
    .d(\PWM7/pnumr [23]),
    .o(_al_u2277_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2278 (
    .a(_al_u2277_o),
    .b(\PWM7/n24 ),
    .c(pnumcnt7[23]),
    .d(\PWM7/pnumr [23]),
    .e(pwm_start_stop[23]),
    .o(\PWM7/n31 [23]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2279 (
    .a(\PWM7/n24 ),
    .b(\PWM7/n25_neg_lutinv ),
    .c(\PWM7/n26 [22]),
    .d(\PWM7/pnumr [22]),
    .o(_al_u2279_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u228 (
    .a(\PWM1/pnumr [30]),
    .b(pnum1[30]),
    .c(pnum1[32]),
    .d(pwm_start_stop[17]),
    .o(\PWM1/n23 [30]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2280 (
    .a(_al_u2279_o),
    .b(\PWM7/n24 ),
    .c(pnumcnt7[22]),
    .d(\PWM7/pnumr [22]),
    .e(pwm_start_stop[23]),
    .o(\PWM7/n31 [22]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2281 (
    .a(\PWM7/n24 ),
    .b(\PWM7/n25_neg_lutinv ),
    .c(\PWM7/n26 [21]),
    .d(\PWM7/pnumr [21]),
    .o(_al_u2281_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2282 (
    .a(_al_u2281_o),
    .b(\PWM7/n24 ),
    .c(pnumcnt7[21]),
    .d(\PWM7/pnumr [21]),
    .e(pwm_start_stop[23]),
    .o(\PWM7/n31 [21]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2283 (
    .a(\PWM7/n24 ),
    .b(\PWM7/n25_neg_lutinv ),
    .c(\PWM7/n26 [20]),
    .d(\PWM7/pnumr [20]),
    .o(_al_u2283_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2284 (
    .a(_al_u2283_o),
    .b(\PWM7/n24 ),
    .c(pnumcnt7[20]),
    .d(\PWM7/pnumr [20]),
    .e(pwm_start_stop[23]),
    .o(\PWM7/n31 [20]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2285 (
    .a(\PWM7/n24 ),
    .b(\PWM7/n25_neg_lutinv ),
    .c(\PWM7/n26 [2]),
    .d(\PWM7/pnumr [2]),
    .o(_al_u2285_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2286 (
    .a(_al_u2285_o),
    .b(\PWM7/n24 ),
    .c(pnumcnt7[2]),
    .d(\PWM7/pnumr [2]),
    .e(pwm_start_stop[23]),
    .o(\PWM7/n31 [2]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2287 (
    .a(\PWM7/n24 ),
    .b(\PWM7/n25_neg_lutinv ),
    .c(\PWM7/n26 [19]),
    .d(\PWM7/pnumr [19]),
    .o(_al_u2287_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2288 (
    .a(_al_u2287_o),
    .b(\PWM7/n24 ),
    .c(pnumcnt7[19]),
    .d(\PWM7/pnumr [19]),
    .e(pwm_start_stop[23]),
    .o(\PWM7/n31 [19]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2289 (
    .a(\PWM7/n24 ),
    .b(\PWM7/n25_neg_lutinv ),
    .c(\PWM7/n26 [18]),
    .d(\PWM7/pnumr [18]),
    .o(_al_u2289_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u229 (
    .a(\PWM1/pnumr [3]),
    .b(pnum1[3]),
    .c(pnum1[32]),
    .d(pwm_start_stop[17]),
    .o(\PWM1/n23 [3]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2290 (
    .a(_al_u2289_o),
    .b(\PWM7/n24 ),
    .c(pnumcnt7[18]),
    .d(\PWM7/pnumr [18]),
    .e(pwm_start_stop[23]),
    .o(\PWM7/n31 [18]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2291 (
    .a(\PWM7/n24 ),
    .b(\PWM7/n25_neg_lutinv ),
    .c(\PWM7/n26 [17]),
    .d(\PWM7/pnumr [17]),
    .o(_al_u2291_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2292 (
    .a(_al_u2291_o),
    .b(\PWM7/n24 ),
    .c(pnumcnt7[17]),
    .d(\PWM7/pnumr [17]),
    .e(pwm_start_stop[23]),
    .o(\PWM7/n31 [17]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2293 (
    .a(\PWM7/n24 ),
    .b(\PWM7/n25_neg_lutinv ),
    .c(\PWM7/n26 [16]),
    .d(\PWM7/pnumr [16]),
    .o(_al_u2293_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2294 (
    .a(_al_u2293_o),
    .b(\PWM7/n24 ),
    .c(pnumcnt7[16]),
    .d(\PWM7/pnumr [16]),
    .e(pwm_start_stop[23]),
    .o(\PWM7/n31 [16]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2295 (
    .a(\PWM7/n24 ),
    .b(\PWM7/n25_neg_lutinv ),
    .c(\PWM7/n26 [15]),
    .d(\PWM7/pnumr [15]),
    .o(_al_u2295_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2296 (
    .a(_al_u2295_o),
    .b(\PWM7/n24 ),
    .c(pnumcnt7[15]),
    .d(\PWM7/pnumr [15]),
    .e(pwm_start_stop[23]),
    .o(\PWM7/n31 [15]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2297 (
    .a(\PWM7/n24 ),
    .b(\PWM7/n25_neg_lutinv ),
    .c(\PWM7/n26 [14]),
    .d(\PWM7/pnumr [14]),
    .o(_al_u2297_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2298 (
    .a(_al_u2297_o),
    .b(\PWM7/n24 ),
    .c(pnumcnt7[14]),
    .d(\PWM7/pnumr [14]),
    .e(pwm_start_stop[23]),
    .o(\PWM7/n31 [14]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2299 (
    .a(\PWM7/n24 ),
    .b(\PWM7/n25_neg_lutinv ),
    .c(\PWM7/n26 [13]),
    .d(\PWM7/pnumr [13]),
    .o(_al_u2299_o));
  EF2_PHY_PAD #(
    //.LOCATION("P142"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u23 (
    .do({open_n754,open_n755,open_n756,dir_pad[15]}),
    .opad(dir[15]));  // CPLD_SOC_AHB_TOP.v(7)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u230 (
    .a(\PWM1/pnumr [29]),
    .b(pnum1[29]),
    .c(pnum1[32]),
    .d(pwm_start_stop[17]),
    .o(\PWM1/n23 [29]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2300 (
    .a(_al_u2299_o),
    .b(\PWM7/n24 ),
    .c(pnumcnt7[13]),
    .d(\PWM7/pnumr [13]),
    .e(pwm_start_stop[23]),
    .o(\PWM7/n31 [13]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2301 (
    .a(\PWM7/n24 ),
    .b(\PWM7/n25_neg_lutinv ),
    .c(\PWM7/n26 [12]),
    .d(\PWM7/pnumr [12]),
    .o(_al_u2301_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2302 (
    .a(_al_u2301_o),
    .b(\PWM7/n24 ),
    .c(pnumcnt7[12]),
    .d(\PWM7/pnumr [12]),
    .e(pwm_start_stop[23]),
    .o(\PWM7/n31 [12]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2303 (
    .a(\PWM7/n24 ),
    .b(\PWM7/n25_neg_lutinv ),
    .c(\PWM7/n26 [11]),
    .d(\PWM7/pnumr [11]),
    .o(_al_u2303_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2304 (
    .a(_al_u2303_o),
    .b(\PWM7/n24 ),
    .c(pnumcnt7[11]),
    .d(\PWM7/pnumr [11]),
    .e(pwm_start_stop[23]),
    .o(\PWM7/n31 [11]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2305 (
    .a(\PWM7/n24 ),
    .b(\PWM7/n25_neg_lutinv ),
    .c(\PWM7/n26 [10]),
    .d(\PWM7/pnumr [10]),
    .o(_al_u2305_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2306 (
    .a(_al_u2305_o),
    .b(\PWM7/n24 ),
    .c(pnumcnt7[10]),
    .d(\PWM7/pnumr [10]),
    .e(pwm_start_stop[23]),
    .o(\PWM7/n31 [10]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2307 (
    .a(\PWM7/n24 ),
    .b(\PWM7/n25_neg_lutinv ),
    .c(\PWM7/n26 [1]),
    .d(\PWM7/pnumr [1]),
    .o(_al_u2307_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2308 (
    .a(_al_u2307_o),
    .b(\PWM7/n24 ),
    .c(pnumcnt7[1]),
    .d(\PWM7/pnumr [1]),
    .e(pwm_start_stop[23]),
    .o(\PWM7/n31 [1]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2309 (
    .a(\PWM7/n24 ),
    .b(\PWM7/n25_neg_lutinv ),
    .c(\PWM7/n26 [0]),
    .d(\PWM7/pnumr [0]),
    .o(_al_u2309_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u231 (
    .a(\PWM1/pnumr [28]),
    .b(pnum1[28]),
    .c(pnum1[32]),
    .d(pwm_start_stop[17]),
    .o(\PWM1/n23 [28]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2310 (
    .a(_al_u2309_o),
    .b(\PWM7/n24 ),
    .c(pnumcnt7[0]),
    .d(\PWM7/pnumr [0]),
    .e(pwm_start_stop[23]),
    .o(\PWM7/n31 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(D*~A))"),
    .INIT(16'h8acf))
    _al_u2311 (
    .a(\PWM7/FreCnt [1]),
    .b(\PWM7/FreCnt [15]),
    .c(\PWM7/FreCntr [16]),
    .d(\PWM7/FreCntr [2]),
    .o(_al_u2311_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u2312 (
    .a(_al_u2311_o),
    .b(\PWM7/FreCnt [4]),
    .c(\PWM7/FreCntr [5]),
    .o(_al_u2312_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u2313 (
    .a(\PWM7/FreCnt [15]),
    .b(\PWM7/FreCnt [3]),
    .c(\PWM7/FreCntr [16]),
    .d(\PWM7/FreCntr [4]),
    .o(_al_u2313_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D@C))"),
    .INIT(16'h8008))
    _al_u2314 (
    .a(_al_u2312_o),
    .b(_al_u2313_o),
    .c(\PWM7/FreCnt [14]),
    .d(\PWM7/FreCntr [15]),
    .o(_al_u2314_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u2315 (
    .a(\PWM7/FreCnt [10]),
    .b(\PWM7/FreCnt [19]),
    .c(\PWM7/FreCntr [11]),
    .d(\PWM7/FreCntr [20]),
    .o(_al_u2315_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*~C)*~(~D*B))"),
    .INIT(32'ha020aa22))
    _al_u2316 (
    .a(_al_u2315_o),
    .b(\PWM7/FreCnt [12]),
    .c(\PWM7/FreCnt [5]),
    .d(\PWM7/FreCntr [13]),
    .e(\PWM7/FreCntr [6]),
    .o(_al_u2316_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u2317 (
    .a(\PWM7/FreCnt [12]),
    .b(\PWM7/FreCnt [17]),
    .c(\PWM7/FreCntr [13]),
    .d(\PWM7/FreCntr [18]),
    .o(_al_u2317_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*C)*~(D*~B))"),
    .INIT(32'h88aa080a))
    _al_u2318 (
    .a(_al_u2317_o),
    .b(\PWM7/FreCnt [21]),
    .c(\PWM7/FreCnt [23]),
    .d(\PWM7/FreCntr [22]),
    .e(\PWM7/FreCntr [24]),
    .o(_al_u2318_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u2319 (
    .a(_al_u2314_o),
    .b(_al_u2316_o),
    .c(_al_u2318_o),
    .o(_al_u2319_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u232 (
    .a(\PWM1/pnumr [27]),
    .b(pnum1[27]),
    .c(pnum1[32]),
    .d(pwm_start_stop[17]),
    .o(\PWM1/n23 [27]));
  AL_MAP_LUT4 #(
    .EQN("(~(C@B)*~(D@A))"),
    .INIT(16'h8241))
    _al_u2320 (
    .a(\PWM7/FreCnt [24]),
    .b(\PWM7/FreCnt [9]),
    .c(\PWM7/FreCntr [10]),
    .d(\PWM7/FreCntr [25]),
    .o(_al_u2320_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u2321 (
    .a(_al_u2320_o),
    .b(\PWM7/FreCnt [22]),
    .c(\PWM7/FreCntr [23]),
    .o(_al_u2321_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u2322 (
    .a(\PWM7/FreCnt [20]),
    .b(\PWM7/FreCnt [6]),
    .c(\PWM7/FreCntr [21]),
    .d(\PWM7/FreCntr [7]),
    .o(_al_u2322_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u2323 (
    .a(_al_u2322_o),
    .b(\PWM7/FreCnt [18]),
    .c(\PWM7/FreCnt [25]),
    .d(\PWM7/FreCntr [19]),
    .e(\PWM7/FreCntr [26]),
    .o(_al_u2323_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u2324 (
    .a(\PWM7/FreCnt [17]),
    .b(\PWM7/FreCnt [23]),
    .c(\PWM7/FreCntr [18]),
    .d(\PWM7/FreCntr [24]),
    .o(_al_u2324_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*~C)*~(~D*B))"),
    .INIT(32'ha020aa22))
    _al_u2325 (
    .a(_al_u2324_o),
    .b(\PWM7/FreCnt [1]),
    .c(\PWM7/FreCnt [19]),
    .d(\PWM7/FreCntr [2]),
    .e(\PWM7/FreCntr [20]),
    .o(_al_u2325_o));
  AL_MAP_LUT5 #(
    .EQN("(~B*~(E@C)*~(~D*A))"),
    .INIT(32'h30100301))
    _al_u2326 (
    .a(\PWM7/FreCnt [13]),
    .b(\PWM7/FreCnt [26]),
    .c(\PWM7/FreCnt [8]),
    .d(\PWM7/FreCntr [14]),
    .e(\PWM7/FreCntr [9]),
    .o(_al_u2326_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u2327 (
    .a(_al_u2321_o),
    .b(_al_u2323_o),
    .c(_al_u2325_o),
    .d(_al_u2326_o),
    .o(_al_u2327_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u2328 (
    .a(\PWM7/FreCnt [2]),
    .b(\PWM7/FreCnt [5]),
    .c(\PWM7/FreCntr [3]),
    .d(\PWM7/FreCntr [6]),
    .o(_al_u2328_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*~C)*~(D*~B))"),
    .INIT(32'h80a088aa))
    _al_u2329 (
    .a(_al_u2328_o),
    .b(\PWM7/FreCnt [3]),
    .c(\PWM7/FreCnt [7]),
    .d(\PWM7/FreCntr [4]),
    .e(\PWM7/FreCntr [8]),
    .o(_al_u2329_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u233 (
    .a(\PWM1/pnumr [26]),
    .b(pnum1[26]),
    .c(pnum1[32]),
    .d(pwm_start_stop[17]),
    .o(\PWM1/n23 [26]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*~C)*~(D@B))"),
    .INIT(32'h80208822))
    _al_u2330 (
    .a(_al_u2329_o),
    .b(\PWM7/FreCnt [16]),
    .c(\PWM7/FreCnt [2]),
    .d(\PWM7/FreCntr [17]),
    .e(\PWM7/FreCntr [3]),
    .o(_al_u2330_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u2331 (
    .a(\PWM7/FreCnt [11]),
    .b(\PWM7/FreCnt [21]),
    .c(\PWM7/FreCntr [12]),
    .d(\PWM7/FreCntr [22]),
    .o(_al_u2331_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*~C)*~(D*~B))"),
    .INIT(32'h80a088aa))
    _al_u2332 (
    .a(_al_u2331_o),
    .b(\PWM7/FreCnt [10]),
    .c(\PWM7/FreCnt [13]),
    .d(\PWM7/FreCntr [11]),
    .e(\PWM7/FreCntr [14]),
    .o(_al_u2332_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2333 (
    .a(\PWM7/FreCnt [7]),
    .b(\PWM7/FreCntr [8]),
    .o(_al_u2333_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(E*~C)*~(D@B))"),
    .INIT(32'h40104411))
    _al_u2334 (
    .a(_al_u2333_o),
    .b(\PWM7/FreCnt [0]),
    .c(\PWM7/FreCnt [11]),
    .d(\PWM7/FreCntr [1]),
    .e(\PWM7/FreCntr [12]),
    .o(_al_u2334_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    _al_u2335 (
    .a(_al_u2319_o),
    .b(_al_u2327_o),
    .c(_al_u2330_o),
    .d(_al_u2332_o),
    .e(_al_u2334_o),
    .o(_al_u2335_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2336 (
    .a(_al_u2335_o),
    .b(pwm_state_read[7]),
    .o(\PWM7/u14_sel_is_1_o ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2337 (
    .a(\PWM8/n0_lutinv ),
    .b(pwm_state_read[8]),
    .o(\PWM8/n24 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u2338 (
    .a(pnumcnt8[18]),
    .b(pnumcnt8[19]),
    .c(pnumcnt8[1]),
    .d(pnumcnt8[20]),
    .o(_al_u2338_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u2339 (
    .a(_al_u2338_o),
    .b(pnumcnt8[21]),
    .c(pnumcnt8[22]),
    .d(pnumcnt8[23]),
    .e(pnumcnt8[2]),
    .o(_al_u2339_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u234 (
    .a(\PWM1/pnumr [25]),
    .b(pnum1[25]),
    .c(pnum1[32]),
    .d(pwm_start_stop[17]),
    .o(\PWM1/n23 [25]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u2340 (
    .a(_al_u2339_o),
    .b(pnumcnt8[6]),
    .c(pnumcnt8[7]),
    .d(pnumcnt8[8]),
    .e(pnumcnt8[9]),
    .o(_al_u2340_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u2341 (
    .a(pnumcnt8[10]),
    .b(pnumcnt8[11]),
    .c(pnumcnt8[12]),
    .d(pnumcnt8[13]),
    .o(_al_u2341_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u2342 (
    .a(_al_u2341_o),
    .b(pnumcnt8[14]),
    .c(pnumcnt8[15]),
    .d(pnumcnt8[16]),
    .e(pnumcnt8[17]),
    .o(_al_u2342_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u2343 (
    .a(pnumcnt8[3]),
    .b(pnumcnt8[4]),
    .c(pnumcnt8[5]),
    .o(_al_u2343_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u2344 (
    .a(_al_u2340_o),
    .b(_al_u2342_o),
    .c(_al_u2343_o),
    .d(pnumcnt8[0]),
    .o(\PWM8/n25_neg_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2345 (
    .a(\PWM8/n24 ),
    .b(\PWM8/n25_neg_lutinv ),
    .c(\PWM8/n26 [9]),
    .d(\PWM8/pnumr [9]),
    .o(_al_u2345_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2346 (
    .a(_al_u2345_o),
    .b(\PWM8/n24 ),
    .c(pnumcnt8[9]),
    .d(\PWM8/pnumr [9]),
    .e(pwm_start_stop[24]),
    .o(\PWM8/n31 [9]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2347 (
    .a(\PWM8/n24 ),
    .b(\PWM8/n25_neg_lutinv ),
    .c(\PWM8/n26 [8]),
    .d(\PWM8/pnumr [8]),
    .o(_al_u2347_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2348 (
    .a(_al_u2347_o),
    .b(\PWM8/n24 ),
    .c(pnumcnt8[8]),
    .d(\PWM8/pnumr [8]),
    .e(pwm_start_stop[24]),
    .o(\PWM8/n31 [8]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2349 (
    .a(\PWM8/n24 ),
    .b(\PWM8/n25_neg_lutinv ),
    .c(\PWM8/n26 [7]),
    .d(\PWM8/pnumr [7]),
    .o(_al_u2349_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u235 (
    .a(\PWM1/pnumr [24]),
    .b(pnum1[24]),
    .c(pnum1[32]),
    .d(pwm_start_stop[17]),
    .o(\PWM1/n23 [24]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2350 (
    .a(_al_u2349_o),
    .b(\PWM8/n24 ),
    .c(pnumcnt8[7]),
    .d(\PWM8/pnumr [7]),
    .e(pwm_start_stop[24]),
    .o(\PWM8/n31 [7]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2351 (
    .a(\PWM8/n24 ),
    .b(\PWM8/n25_neg_lutinv ),
    .c(\PWM8/n26 [6]),
    .d(\PWM8/pnumr [6]),
    .o(_al_u2351_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2352 (
    .a(_al_u2351_o),
    .b(\PWM8/n24 ),
    .c(pnumcnt8[6]),
    .d(\PWM8/pnumr [6]),
    .e(pwm_start_stop[24]),
    .o(\PWM8/n31 [6]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2353 (
    .a(\PWM8/n24 ),
    .b(\PWM8/n25_neg_lutinv ),
    .c(\PWM8/n26 [5]),
    .d(\PWM8/pnumr [5]),
    .o(_al_u2353_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2354 (
    .a(_al_u2353_o),
    .b(\PWM8/n24 ),
    .c(pnumcnt8[5]),
    .d(\PWM8/pnumr [5]),
    .e(pwm_start_stop[24]),
    .o(\PWM8/n31 [5]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2355 (
    .a(\PWM8/n24 ),
    .b(\PWM8/n25_neg_lutinv ),
    .c(\PWM8/n26 [4]),
    .d(\PWM8/pnumr [4]),
    .o(_al_u2355_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2356 (
    .a(_al_u2355_o),
    .b(\PWM8/n24 ),
    .c(pnumcnt8[4]),
    .d(\PWM8/pnumr [4]),
    .e(pwm_start_stop[24]),
    .o(\PWM8/n31 [4]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2357 (
    .a(\PWM8/n24 ),
    .b(\PWM8/n25_neg_lutinv ),
    .c(\PWM8/n26 [3]),
    .d(\PWM8/pnumr [3]),
    .o(_al_u2357_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2358 (
    .a(_al_u2357_o),
    .b(\PWM8/n24 ),
    .c(pnumcnt8[3]),
    .d(\PWM8/pnumr [3]),
    .e(pwm_start_stop[24]),
    .o(\PWM8/n31 [3]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2359 (
    .a(\PWM8/n24 ),
    .b(\PWM8/n25_neg_lutinv ),
    .c(\PWM8/n26 [23]),
    .d(\PWM8/pnumr [23]),
    .o(_al_u2359_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u236 (
    .a(\PWM1/pnumr [23]),
    .b(pnum1[23]),
    .c(pnum1[32]),
    .d(pwm_start_stop[17]),
    .o(\PWM1/n23 [23]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2360 (
    .a(_al_u2359_o),
    .b(\PWM8/n24 ),
    .c(pnumcnt8[23]),
    .d(\PWM8/pnumr [23]),
    .e(pwm_start_stop[24]),
    .o(\PWM8/n31 [23]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2361 (
    .a(\PWM8/n24 ),
    .b(\PWM8/n25_neg_lutinv ),
    .c(\PWM8/n26 [22]),
    .d(\PWM8/pnumr [22]),
    .o(_al_u2361_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2362 (
    .a(_al_u2361_o),
    .b(\PWM8/n24 ),
    .c(pnumcnt8[22]),
    .d(\PWM8/pnumr [22]),
    .e(pwm_start_stop[24]),
    .o(\PWM8/n31 [22]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2363 (
    .a(\PWM8/n24 ),
    .b(\PWM8/n25_neg_lutinv ),
    .c(\PWM8/n26 [21]),
    .d(\PWM8/pnumr [21]),
    .o(_al_u2363_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2364 (
    .a(_al_u2363_o),
    .b(\PWM8/n24 ),
    .c(pnumcnt8[21]),
    .d(\PWM8/pnumr [21]),
    .e(pwm_start_stop[24]),
    .o(\PWM8/n31 [21]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2365 (
    .a(\PWM8/n24 ),
    .b(\PWM8/n25_neg_lutinv ),
    .c(\PWM8/n26 [20]),
    .d(\PWM8/pnumr [20]),
    .o(_al_u2365_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2366 (
    .a(_al_u2365_o),
    .b(\PWM8/n24 ),
    .c(pnumcnt8[20]),
    .d(\PWM8/pnumr [20]),
    .e(pwm_start_stop[24]),
    .o(\PWM8/n31 [20]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2367 (
    .a(\PWM8/n24 ),
    .b(\PWM8/n25_neg_lutinv ),
    .c(\PWM8/n26 [2]),
    .d(\PWM8/pnumr [2]),
    .o(_al_u2367_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2368 (
    .a(_al_u2367_o),
    .b(\PWM8/n24 ),
    .c(pnumcnt8[2]),
    .d(\PWM8/pnumr [2]),
    .e(pwm_start_stop[24]),
    .o(\PWM8/n31 [2]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2369 (
    .a(\PWM8/n24 ),
    .b(\PWM8/n25_neg_lutinv ),
    .c(\PWM8/n26 [19]),
    .d(\PWM8/pnumr [19]),
    .o(_al_u2369_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u237 (
    .a(\PWM1/pnumr [22]),
    .b(pnum1[22]),
    .c(pnum1[32]),
    .d(pwm_start_stop[17]),
    .o(\PWM1/n23 [22]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2370 (
    .a(_al_u2369_o),
    .b(\PWM8/n24 ),
    .c(pnumcnt8[19]),
    .d(\PWM8/pnumr [19]),
    .e(pwm_start_stop[24]),
    .o(\PWM8/n31 [19]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2371 (
    .a(\PWM8/n24 ),
    .b(\PWM8/n25_neg_lutinv ),
    .c(\PWM8/n26 [18]),
    .d(\PWM8/pnumr [18]),
    .o(_al_u2371_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2372 (
    .a(_al_u2371_o),
    .b(\PWM8/n24 ),
    .c(pnumcnt8[18]),
    .d(\PWM8/pnumr [18]),
    .e(pwm_start_stop[24]),
    .o(\PWM8/n31 [18]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2373 (
    .a(\PWM8/n24 ),
    .b(\PWM8/n25_neg_lutinv ),
    .c(\PWM8/n26 [17]),
    .d(\PWM8/pnumr [17]),
    .o(_al_u2373_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2374 (
    .a(_al_u2373_o),
    .b(\PWM8/n24 ),
    .c(pnumcnt8[17]),
    .d(\PWM8/pnumr [17]),
    .e(pwm_start_stop[24]),
    .o(\PWM8/n31 [17]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2375 (
    .a(\PWM8/n24 ),
    .b(\PWM8/n25_neg_lutinv ),
    .c(\PWM8/n26 [16]),
    .d(\PWM8/pnumr [16]),
    .o(_al_u2375_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2376 (
    .a(_al_u2375_o),
    .b(\PWM8/n24 ),
    .c(pnumcnt8[16]),
    .d(\PWM8/pnumr [16]),
    .e(pwm_start_stop[24]),
    .o(\PWM8/n31 [16]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2377 (
    .a(\PWM8/n24 ),
    .b(\PWM8/n25_neg_lutinv ),
    .c(\PWM8/n26 [15]),
    .d(\PWM8/pnumr [15]),
    .o(_al_u2377_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2378 (
    .a(_al_u2377_o),
    .b(\PWM8/n24 ),
    .c(pnumcnt8[15]),
    .d(\PWM8/pnumr [15]),
    .e(pwm_start_stop[24]),
    .o(\PWM8/n31 [15]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2379 (
    .a(\PWM8/n24 ),
    .b(\PWM8/n25_neg_lutinv ),
    .c(\PWM8/n26 [14]),
    .d(\PWM8/pnumr [14]),
    .o(_al_u2379_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u238 (
    .a(\PWM1/pnumr [21]),
    .b(pnum1[21]),
    .c(pnum1[32]),
    .d(pwm_start_stop[17]),
    .o(\PWM1/n23 [21]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2380 (
    .a(_al_u2379_o),
    .b(\PWM8/n24 ),
    .c(pnumcnt8[14]),
    .d(\PWM8/pnumr [14]),
    .e(pwm_start_stop[24]),
    .o(\PWM8/n31 [14]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2381 (
    .a(\PWM8/n24 ),
    .b(\PWM8/n25_neg_lutinv ),
    .c(\PWM8/n26 [13]),
    .d(\PWM8/pnumr [13]),
    .o(_al_u2381_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2382 (
    .a(_al_u2381_o),
    .b(\PWM8/n24 ),
    .c(pnumcnt8[13]),
    .d(\PWM8/pnumr [13]),
    .e(pwm_start_stop[24]),
    .o(\PWM8/n31 [13]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2383 (
    .a(\PWM8/n24 ),
    .b(\PWM8/n25_neg_lutinv ),
    .c(\PWM8/n26 [12]),
    .d(\PWM8/pnumr [12]),
    .o(_al_u2383_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2384 (
    .a(_al_u2383_o),
    .b(\PWM8/n24 ),
    .c(pnumcnt8[12]),
    .d(\PWM8/pnumr [12]),
    .e(pwm_start_stop[24]),
    .o(\PWM8/n31 [12]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2385 (
    .a(\PWM8/n24 ),
    .b(\PWM8/n25_neg_lutinv ),
    .c(\PWM8/n26 [11]),
    .d(\PWM8/pnumr [11]),
    .o(_al_u2385_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2386 (
    .a(_al_u2385_o),
    .b(\PWM8/n24 ),
    .c(pnumcnt8[11]),
    .d(\PWM8/pnumr [11]),
    .e(pwm_start_stop[24]),
    .o(\PWM8/n31 [11]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2387 (
    .a(\PWM8/n24 ),
    .b(\PWM8/n25_neg_lutinv ),
    .c(\PWM8/n26 [10]),
    .d(\PWM8/pnumr [10]),
    .o(_al_u2387_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2388 (
    .a(_al_u2387_o),
    .b(\PWM8/n24 ),
    .c(pnumcnt8[10]),
    .d(\PWM8/pnumr [10]),
    .e(pwm_start_stop[24]),
    .o(\PWM8/n31 [10]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2389 (
    .a(\PWM8/n24 ),
    .b(\PWM8/n25_neg_lutinv ),
    .c(\PWM8/n26 [1]),
    .d(\PWM8/pnumr [1]),
    .o(_al_u2389_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u239 (
    .a(\PWM1/pnumr [20]),
    .b(pnum1[20]),
    .c(pnum1[32]),
    .d(pwm_start_stop[17]),
    .o(\PWM1/n23 [20]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2390 (
    .a(_al_u2389_o),
    .b(\PWM8/n24 ),
    .c(pnumcnt8[1]),
    .d(\PWM8/pnumr [1]),
    .e(pwm_start_stop[24]),
    .o(\PWM8/n31 [1]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2391 (
    .a(\PWM8/n24 ),
    .b(\PWM8/n25_neg_lutinv ),
    .c(\PWM8/n26 [0]),
    .d(\PWM8/pnumr [0]),
    .o(_al_u2391_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2392 (
    .a(_al_u2391_o),
    .b(\PWM8/n24 ),
    .c(pnumcnt8[0]),
    .d(\PWM8/pnumr [0]),
    .e(pwm_start_stop[24]),
    .o(\PWM8/n31 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u2393 (
    .a(\PWM8/FreCnt [22]),
    .b(\PWM8/FreCnt [8]),
    .c(\PWM8/FreCntr [23]),
    .d(\PWM8/FreCntr [9]),
    .o(_al_u2393_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*C)*~(D*~B))"),
    .INIT(32'h88aa080a))
    _al_u2394 (
    .a(_al_u2393_o),
    .b(\PWM8/FreCnt [10]),
    .c(\PWM8/FreCnt [17]),
    .d(\PWM8/FreCntr [11]),
    .e(\PWM8/FreCntr [18]),
    .o(_al_u2394_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*~C)*~(D@B))"),
    .INIT(32'h80208822))
    _al_u2395 (
    .a(_al_u2394_o),
    .b(\PWM8/FreCnt [11]),
    .c(\PWM8/FreCnt [22]),
    .d(\PWM8/FreCntr [12]),
    .e(\PWM8/FreCntr [23]),
    .o(_al_u2395_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u2396 (
    .a(\PWM8/FreCnt [1]),
    .b(\PWM8/FreCnt [5]),
    .c(\PWM8/FreCntr [2]),
    .d(\PWM8/FreCntr [6]),
    .o(_al_u2396_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C@B)*~(D@A))"),
    .INIT(16'h8241))
    _al_u2397 (
    .a(\PWM8/FreCnt [16]),
    .b(\PWM8/FreCnt [9]),
    .c(\PWM8/FreCntr [10]),
    .d(\PWM8/FreCntr [17]),
    .o(_al_u2397_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u2398 (
    .a(_al_u2395_o),
    .b(_al_u2396_o),
    .c(_al_u2397_o),
    .d(\PWM8/FreCnt [12]),
    .e(\PWM8/FreCntr [13]),
    .o(_al_u2398_o));
  AL_MAP_LUT5 #(
    .EQN("(~B*~(E@C)*~(~D*A))"),
    .INIT(32'h30100301))
    _al_u2399 (
    .a(\PWM8/FreCnt [23]),
    .b(\PWM8/FreCnt [26]),
    .c(\PWM8/FreCnt [4]),
    .d(\PWM8/FreCntr [24]),
    .e(\PWM8/FreCntr [5]),
    .o(_al_u2399_o));
  EF2_PHY_PAD #(
    //.LOCATION("P54"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u24 (
    .do({open_n777,open_n778,open_n779,dir_pad[14]}),
    .opad(dir[14]));  // CPLD_SOC_AHB_TOP.v(7)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u240 (
    .a(\PWM1/pnumr [2]),
    .b(pnum1[2]),
    .c(pnum1[32]),
    .d(pwm_start_stop[17]),
    .o(\PWM1/n23 [2]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D@C)*~(E@B))"),
    .INIT(32'h80082002))
    _al_u2400 (
    .a(_al_u2399_o),
    .b(\PWM8/FreCnt [2]),
    .c(\PWM8/FreCnt [24]),
    .d(\PWM8/FreCntr [25]),
    .e(\PWM8/FreCntr [3]),
    .o(_al_u2400_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u2401 (
    .a(\PWM8/FreCnt [18]),
    .b(\PWM8/FreCnt [6]),
    .c(\PWM8/FreCntr [19]),
    .d(\PWM8/FreCntr [7]),
    .o(_al_u2401_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u2402 (
    .a(_al_u2401_o),
    .b(\PWM8/FreCnt [0]),
    .c(\PWM8/FreCntr [1]),
    .o(_al_u2402_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u2403 (
    .a(\PWM8/FreCnt [21]),
    .b(\PWM8/FreCnt [7]),
    .c(\PWM8/FreCntr [22]),
    .d(\PWM8/FreCntr [8]),
    .o(_al_u2403_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*~C)*~(~D*B))"),
    .INIT(32'ha020aa22))
    _al_u2404 (
    .a(_al_u2403_o),
    .b(\PWM8/FreCnt [25]),
    .c(\PWM8/FreCnt [3]),
    .d(\PWM8/FreCntr [26]),
    .e(\PWM8/FreCntr [4]),
    .o(_al_u2404_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u2405 (
    .a(\PWM8/FreCnt [7]),
    .b(\PWM8/FreCnt [8]),
    .c(\PWM8/FreCntr [8]),
    .d(\PWM8/FreCntr [9]),
    .o(_al_u2405_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*C)*~(~D*B))"),
    .INIT(32'haa220a02))
    _al_u2406 (
    .a(_al_u2405_o),
    .b(\PWM8/FreCnt [21]),
    .c(\PWM8/FreCnt [3]),
    .d(\PWM8/FreCntr [22]),
    .e(\PWM8/FreCntr [4]),
    .o(_al_u2406_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u2407 (
    .a(_al_u2400_o),
    .b(_al_u2402_o),
    .c(_al_u2404_o),
    .d(_al_u2406_o),
    .o(_al_u2407_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u2408 (
    .a(\PWM8/FreCnt [14]),
    .b(\PWM8/FreCnt [20]),
    .c(\PWM8/FreCntr [15]),
    .d(\PWM8/FreCntr [21]),
    .o(_al_u2408_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u2409 (
    .a(\PWM8/FreCnt [15]),
    .b(\PWM8/FreCnt [23]),
    .c(\PWM8/FreCntr [16]),
    .d(\PWM8/FreCntr [24]),
    .o(_al_u2409_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u241 (
    .a(\PWM1/pnumr [19]),
    .b(pnum1[19]),
    .c(pnum1[32]),
    .d(pwm_start_stop[17]),
    .o(\PWM1/n23 [19]));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D@C))"),
    .INIT(16'h8008))
    _al_u2410 (
    .a(_al_u2408_o),
    .b(_al_u2409_o),
    .c(\PWM8/FreCnt [13]),
    .d(\PWM8/FreCntr [14]),
    .o(_al_u2410_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u2411 (
    .a(\PWM8/FreCnt [10]),
    .b(\PWM8/FreCnt [5]),
    .c(\PWM8/FreCntr [11]),
    .d(\PWM8/FreCntr [6]),
    .o(_al_u2411_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*~C)*~(D*~B))"),
    .INIT(32'h80a088aa))
    _al_u2412 (
    .a(_al_u2411_o),
    .b(\PWM8/FreCnt [15]),
    .c(\PWM8/FreCnt [25]),
    .d(\PWM8/FreCntr [16]),
    .e(\PWM8/FreCntr [26]),
    .o(_al_u2412_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2413 (
    .a(\PWM8/FreCnt [1]),
    .b(\PWM8/FreCntr [2]),
    .o(_al_u2413_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(E@C)*~(D*~B))"),
    .INIT(32'h40500405))
    _al_u2414 (
    .a(_al_u2413_o),
    .b(\PWM8/FreCnt [17]),
    .c(\PWM8/FreCnt [19]),
    .d(\PWM8/FreCntr [18]),
    .e(\PWM8/FreCntr [20]),
    .o(_al_u2414_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    _al_u2415 (
    .a(_al_u2398_o),
    .b(_al_u2407_o),
    .c(_al_u2410_o),
    .d(_al_u2412_o),
    .e(_al_u2414_o),
    .o(_al_u2415_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2416 (
    .a(_al_u2415_o),
    .b(pwm_state_read[8]),
    .o(\PWM8/u14_sel_is_1_o ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2417 (
    .a(\PWM9/n0_lutinv ),
    .b(pwm_state_read[9]),
    .o(\PWM9/n24 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u2418 (
    .a(pnumcnt9[18]),
    .b(pnumcnt9[19]),
    .c(pnumcnt9[1]),
    .d(pnumcnt9[20]),
    .o(_al_u2418_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u2419 (
    .a(_al_u2418_o),
    .b(pnumcnt9[21]),
    .c(pnumcnt9[22]),
    .d(pnumcnt9[23]),
    .e(pnumcnt9[2]),
    .o(_al_u2419_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u242 (
    .a(\PWM1/pnumr [18]),
    .b(pnum1[18]),
    .c(pnum1[32]),
    .d(pwm_start_stop[17]),
    .o(\PWM1/n23 [18]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u2420 (
    .a(_al_u2419_o),
    .b(pnumcnt9[6]),
    .c(pnumcnt9[7]),
    .d(pnumcnt9[8]),
    .e(pnumcnt9[9]),
    .o(_al_u2420_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u2421 (
    .a(pnumcnt9[10]),
    .b(pnumcnt9[11]),
    .c(pnumcnt9[12]),
    .d(pnumcnt9[13]),
    .o(_al_u2421_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u2422 (
    .a(_al_u2421_o),
    .b(pnumcnt9[14]),
    .c(pnumcnt9[15]),
    .d(pnumcnt9[16]),
    .e(pnumcnt9[17]),
    .o(_al_u2422_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u2423 (
    .a(pnumcnt9[3]),
    .b(pnumcnt9[4]),
    .c(pnumcnt9[5]),
    .o(_al_u2423_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u2424 (
    .a(_al_u2420_o),
    .b(_al_u2422_o),
    .c(_al_u2423_o),
    .d(pnumcnt9[0]),
    .o(\PWM9/n25_neg_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2425 (
    .a(\PWM9/n24 ),
    .b(\PWM9/n25_neg_lutinv ),
    .c(\PWM9/n26 [9]),
    .d(\PWM9/pnumr [9]),
    .o(_al_u2425_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2426 (
    .a(_al_u2425_o),
    .b(\PWM9/n24 ),
    .c(pnumcnt9[9]),
    .d(\PWM9/pnumr [9]),
    .e(pwm_start_stop[25]),
    .o(\PWM9/n31 [9]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2427 (
    .a(\PWM9/n24 ),
    .b(\PWM9/n25_neg_lutinv ),
    .c(\PWM9/n26 [8]),
    .d(\PWM9/pnumr [8]),
    .o(_al_u2427_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2428 (
    .a(_al_u2427_o),
    .b(\PWM9/n24 ),
    .c(pnumcnt9[8]),
    .d(\PWM9/pnumr [8]),
    .e(pwm_start_stop[25]),
    .o(\PWM9/n31 [8]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2429 (
    .a(\PWM9/n24 ),
    .b(\PWM9/n25_neg_lutinv ),
    .c(\PWM9/n26 [7]),
    .d(\PWM9/pnumr [7]),
    .o(_al_u2429_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u243 (
    .a(\PWM1/pnumr [17]),
    .b(pnum1[17]),
    .c(pnum1[32]),
    .d(pwm_start_stop[17]),
    .o(\PWM1/n23 [17]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2430 (
    .a(_al_u2429_o),
    .b(\PWM9/n24 ),
    .c(pnumcnt9[7]),
    .d(\PWM9/pnumr [7]),
    .e(pwm_start_stop[25]),
    .o(\PWM9/n31 [7]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2431 (
    .a(\PWM9/n24 ),
    .b(\PWM9/n25_neg_lutinv ),
    .c(\PWM9/n26 [6]),
    .d(\PWM9/pnumr [6]),
    .o(_al_u2431_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2432 (
    .a(_al_u2431_o),
    .b(\PWM9/n24 ),
    .c(pnumcnt9[6]),
    .d(\PWM9/pnumr [6]),
    .e(pwm_start_stop[25]),
    .o(\PWM9/n31 [6]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2433 (
    .a(\PWM9/n24 ),
    .b(\PWM9/n25_neg_lutinv ),
    .c(\PWM9/n26 [5]),
    .d(\PWM9/pnumr [5]),
    .o(_al_u2433_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2434 (
    .a(_al_u2433_o),
    .b(\PWM9/n24 ),
    .c(pnumcnt9[5]),
    .d(\PWM9/pnumr [5]),
    .e(pwm_start_stop[25]),
    .o(\PWM9/n31 [5]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2435 (
    .a(\PWM9/n24 ),
    .b(\PWM9/n25_neg_lutinv ),
    .c(\PWM9/n26 [4]),
    .d(\PWM9/pnumr [4]),
    .o(_al_u2435_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2436 (
    .a(_al_u2435_o),
    .b(\PWM9/n24 ),
    .c(pnumcnt9[4]),
    .d(\PWM9/pnumr [4]),
    .e(pwm_start_stop[25]),
    .o(\PWM9/n31 [4]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2437 (
    .a(\PWM9/n24 ),
    .b(\PWM9/n25_neg_lutinv ),
    .c(\PWM9/n26 [3]),
    .d(\PWM9/pnumr [3]),
    .o(_al_u2437_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2438 (
    .a(_al_u2437_o),
    .b(\PWM9/n24 ),
    .c(pnumcnt9[3]),
    .d(\PWM9/pnumr [3]),
    .e(pwm_start_stop[25]),
    .o(\PWM9/n31 [3]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2439 (
    .a(\PWM9/n24 ),
    .b(\PWM9/n25_neg_lutinv ),
    .c(\PWM9/n26 [23]),
    .d(\PWM9/pnumr [23]),
    .o(_al_u2439_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u244 (
    .a(\PWM1/pnumr [16]),
    .b(pnum1[16]),
    .c(pnum1[32]),
    .d(pwm_start_stop[17]),
    .o(\PWM1/n23 [16]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2440 (
    .a(_al_u2439_o),
    .b(\PWM9/n24 ),
    .c(pnumcnt9[23]),
    .d(\PWM9/pnumr [23]),
    .e(pwm_start_stop[25]),
    .o(\PWM9/n31 [23]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2441 (
    .a(\PWM9/n24 ),
    .b(\PWM9/n25_neg_lutinv ),
    .c(\PWM9/n26 [22]),
    .d(\PWM9/pnumr [22]),
    .o(_al_u2441_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2442 (
    .a(_al_u2441_o),
    .b(\PWM9/n24 ),
    .c(pnumcnt9[22]),
    .d(\PWM9/pnumr [22]),
    .e(pwm_start_stop[25]),
    .o(\PWM9/n31 [22]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2443 (
    .a(\PWM9/n24 ),
    .b(\PWM9/n25_neg_lutinv ),
    .c(\PWM9/n26 [21]),
    .d(\PWM9/pnumr [21]),
    .o(_al_u2443_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2444 (
    .a(_al_u2443_o),
    .b(\PWM9/n24 ),
    .c(pnumcnt9[21]),
    .d(\PWM9/pnumr [21]),
    .e(pwm_start_stop[25]),
    .o(\PWM9/n31 [21]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2445 (
    .a(\PWM9/n24 ),
    .b(\PWM9/n25_neg_lutinv ),
    .c(\PWM9/n26 [20]),
    .d(\PWM9/pnumr [20]),
    .o(_al_u2445_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2446 (
    .a(_al_u2445_o),
    .b(\PWM9/n24 ),
    .c(pnumcnt9[20]),
    .d(\PWM9/pnumr [20]),
    .e(pwm_start_stop[25]),
    .o(\PWM9/n31 [20]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2447 (
    .a(\PWM9/n24 ),
    .b(\PWM9/n25_neg_lutinv ),
    .c(\PWM9/n26 [2]),
    .d(\PWM9/pnumr [2]),
    .o(_al_u2447_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2448 (
    .a(_al_u2447_o),
    .b(\PWM9/n24 ),
    .c(pnumcnt9[2]),
    .d(\PWM9/pnumr [2]),
    .e(pwm_start_stop[25]),
    .o(\PWM9/n31 [2]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2449 (
    .a(\PWM9/n24 ),
    .b(\PWM9/n25_neg_lutinv ),
    .c(\PWM9/n26 [19]),
    .d(\PWM9/pnumr [19]),
    .o(_al_u2449_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u245 (
    .a(\PWM1/pnumr [15]),
    .b(pnum1[15]),
    .c(pnum1[32]),
    .d(pwm_start_stop[17]),
    .o(\PWM1/n23 [15]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2450 (
    .a(_al_u2449_o),
    .b(\PWM9/n24 ),
    .c(pnumcnt9[19]),
    .d(\PWM9/pnumr [19]),
    .e(pwm_start_stop[25]),
    .o(\PWM9/n31 [19]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2451 (
    .a(\PWM9/n24 ),
    .b(\PWM9/n25_neg_lutinv ),
    .c(\PWM9/n26 [18]),
    .d(\PWM9/pnumr [18]),
    .o(_al_u2451_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2452 (
    .a(_al_u2451_o),
    .b(\PWM9/n24 ),
    .c(pnumcnt9[18]),
    .d(\PWM9/pnumr [18]),
    .e(pwm_start_stop[25]),
    .o(\PWM9/n31 [18]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2453 (
    .a(\PWM9/n24 ),
    .b(\PWM9/n25_neg_lutinv ),
    .c(\PWM9/n26 [17]),
    .d(\PWM9/pnumr [17]),
    .o(_al_u2453_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2454 (
    .a(_al_u2453_o),
    .b(\PWM9/n24 ),
    .c(pnumcnt9[17]),
    .d(\PWM9/pnumr [17]),
    .e(pwm_start_stop[25]),
    .o(\PWM9/n31 [17]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2455 (
    .a(\PWM9/n24 ),
    .b(\PWM9/n25_neg_lutinv ),
    .c(\PWM9/n26 [16]),
    .d(\PWM9/pnumr [16]),
    .o(_al_u2455_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2456 (
    .a(_al_u2455_o),
    .b(\PWM9/n24 ),
    .c(pnumcnt9[16]),
    .d(\PWM9/pnumr [16]),
    .e(pwm_start_stop[25]),
    .o(\PWM9/n31 [16]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2457 (
    .a(\PWM9/n24 ),
    .b(\PWM9/n25_neg_lutinv ),
    .c(\PWM9/n26 [15]),
    .d(\PWM9/pnumr [15]),
    .o(_al_u2457_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2458 (
    .a(_al_u2457_o),
    .b(\PWM9/n24 ),
    .c(pnumcnt9[15]),
    .d(\PWM9/pnumr [15]),
    .e(pwm_start_stop[25]),
    .o(\PWM9/n31 [15]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2459 (
    .a(\PWM9/n24 ),
    .b(\PWM9/n25_neg_lutinv ),
    .c(\PWM9/n26 [14]),
    .d(\PWM9/pnumr [14]),
    .o(_al_u2459_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u246 (
    .a(\PWM1/pnumr [14]),
    .b(pnum1[14]),
    .c(pnum1[32]),
    .d(pwm_start_stop[17]),
    .o(\PWM1/n23 [14]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2460 (
    .a(_al_u2459_o),
    .b(\PWM9/n24 ),
    .c(pnumcnt9[14]),
    .d(\PWM9/pnumr [14]),
    .e(pwm_start_stop[25]),
    .o(\PWM9/n31 [14]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2461 (
    .a(\PWM9/n24 ),
    .b(\PWM9/n25_neg_lutinv ),
    .c(\PWM9/n26 [13]),
    .d(\PWM9/pnumr [13]),
    .o(_al_u2461_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2462 (
    .a(_al_u2461_o),
    .b(\PWM9/n24 ),
    .c(pnumcnt9[13]),
    .d(\PWM9/pnumr [13]),
    .e(pwm_start_stop[25]),
    .o(\PWM9/n31 [13]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2463 (
    .a(\PWM9/n24 ),
    .b(\PWM9/n25_neg_lutinv ),
    .c(\PWM9/n26 [12]),
    .d(\PWM9/pnumr [12]),
    .o(_al_u2463_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2464 (
    .a(_al_u2463_o),
    .b(\PWM9/n24 ),
    .c(pnumcnt9[12]),
    .d(\PWM9/pnumr [12]),
    .e(pwm_start_stop[25]),
    .o(\PWM9/n31 [12]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2465 (
    .a(\PWM9/n24 ),
    .b(\PWM9/n25_neg_lutinv ),
    .c(\PWM9/n26 [11]),
    .d(\PWM9/pnumr [11]),
    .o(_al_u2465_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2466 (
    .a(_al_u2465_o),
    .b(\PWM9/n24 ),
    .c(pnumcnt9[11]),
    .d(\PWM9/pnumr [11]),
    .e(pwm_start_stop[25]),
    .o(\PWM9/n31 [11]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2467 (
    .a(\PWM9/n24 ),
    .b(\PWM9/n25_neg_lutinv ),
    .c(\PWM9/n26 [10]),
    .d(\PWM9/pnumr [10]),
    .o(_al_u2467_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2468 (
    .a(_al_u2467_o),
    .b(\PWM9/n24 ),
    .c(pnumcnt9[10]),
    .d(\PWM9/pnumr [10]),
    .e(pwm_start_stop[25]),
    .o(\PWM9/n31 [10]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2469 (
    .a(\PWM9/n24 ),
    .b(\PWM9/n25_neg_lutinv ),
    .c(\PWM9/n26 [1]),
    .d(\PWM9/pnumr [1]),
    .o(_al_u2469_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u247 (
    .a(\PWM1/pnumr [13]),
    .b(pnum1[13]),
    .c(pnum1[32]),
    .d(pwm_start_stop[17]),
    .o(\PWM1/n23 [13]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2470 (
    .a(_al_u2469_o),
    .b(\PWM9/n24 ),
    .c(pnumcnt9[1]),
    .d(\PWM9/pnumr [1]),
    .e(pwm_start_stop[25]),
    .o(\PWM9/n31 [1]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2471 (
    .a(\PWM9/n24 ),
    .b(\PWM9/n25_neg_lutinv ),
    .c(\PWM9/n26 [0]),
    .d(\PWM9/pnumr [0]),
    .o(_al_u2471_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2472 (
    .a(_al_u2471_o),
    .b(\PWM9/n24 ),
    .c(pnumcnt9[0]),
    .d(\PWM9/pnumr [0]),
    .e(pwm_start_stop[25]),
    .o(\PWM9/n31 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u2473 (
    .a(\PWM9/FreCnt [10]),
    .b(\PWM9/FreCnt [3]),
    .c(\PWM9/FreCntr [11]),
    .d(\PWM9/FreCntr [4]),
    .o(_al_u2473_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*C)*~(D*~B))"),
    .INIT(32'h88aa080a))
    _al_u2474 (
    .a(_al_u2473_o),
    .b(\PWM9/FreCnt [1]),
    .c(\PWM9/FreCnt [5]),
    .d(\PWM9/FreCntr [2]),
    .e(\PWM9/FreCntr [6]),
    .o(_al_u2474_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*C)*~(D@B))"),
    .INIT(32'h88220802))
    _al_u2475 (
    .a(_al_u2474_o),
    .b(\PWM9/FreCnt [14]),
    .c(\PWM9/FreCnt [8]),
    .d(\PWM9/FreCntr [15]),
    .e(\PWM9/FreCntr [9]),
    .o(_al_u2475_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u2476 (
    .a(\PWM9/FreCnt [12]),
    .b(\PWM9/FreCnt [21]),
    .c(\PWM9/FreCntr [13]),
    .d(\PWM9/FreCntr [22]),
    .o(_al_u2476_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u2477 (
    .a(_al_u2476_o),
    .b(\PWM9/FreCnt [16]),
    .c(\PWM9/FreCntr [17]),
    .o(_al_u2477_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u2478 (
    .a(\PWM9/FreCnt [13]),
    .b(\PWM9/FreCnt [17]),
    .c(\PWM9/FreCntr [14]),
    .d(\PWM9/FreCntr [18]),
    .o(_al_u2478_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u2479 (
    .a(_al_u2475_o),
    .b(_al_u2477_o),
    .c(_al_u2478_o),
    .d(\PWM9/FreCnt [9]),
    .e(\PWM9/FreCntr [10]),
    .o(_al_u2479_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u248 (
    .a(\PWM1/pnumr [12]),
    .b(pnum1[12]),
    .c(pnum1[32]),
    .d(pwm_start_stop[17]),
    .o(\PWM1/n23 [12]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u2480 (
    .a(\PWM9/FreCnt [1]),
    .b(\PWM9/FreCnt [23]),
    .c(\PWM9/FreCntr [2]),
    .d(\PWM9/FreCntr [24]),
    .o(_al_u2480_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*~C)*~(~D*B))"),
    .INIT(32'ha020aa22))
    _al_u2481 (
    .a(_al_u2480_o),
    .b(\PWM9/FreCnt [12]),
    .c(\PWM9/FreCnt [5]),
    .d(\PWM9/FreCntr [13]),
    .e(\PWM9/FreCntr [6]),
    .o(_al_u2481_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u2482 (
    .a(\PWM9/FreCnt [13]),
    .b(\PWM9/FreCnt [7]),
    .c(\PWM9/FreCntr [14]),
    .d(\PWM9/FreCntr [8]),
    .o(_al_u2482_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*C)*~(D*~B))"),
    .INIT(32'h88aa080a))
    _al_u2483 (
    .a(_al_u2482_o),
    .b(\PWM9/FreCnt [18]),
    .c(\PWM9/FreCnt [23]),
    .d(\PWM9/FreCntr [19]),
    .e(\PWM9/FreCntr [24]),
    .o(_al_u2483_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2484 (
    .a(\PWM9/FreCnt [10]),
    .b(\PWM9/FreCntr [11]),
    .o(_al_u2484_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(E*~C)*~(D@B))"),
    .INIT(32'h40104411))
    _al_u2485 (
    .a(_al_u2484_o),
    .b(\PWM9/FreCnt [22]),
    .c(\PWM9/FreCnt [3]),
    .d(\PWM9/FreCntr [23]),
    .e(\PWM9/FreCntr [4]),
    .o(_al_u2485_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2486 (
    .a(\PWM9/FreCnt [18]),
    .b(\PWM9/FreCntr [19]),
    .o(_al_u2486_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(E@C)*~(~D*B))"),
    .INIT(32'h50100501))
    _al_u2487 (
    .a(_al_u2486_o),
    .b(\PWM9/FreCnt [15]),
    .c(\PWM9/FreCnt [20]),
    .d(\PWM9/FreCntr [16]),
    .e(\PWM9/FreCntr [21]),
    .o(_al_u2487_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    _al_u2488 (
    .a(_al_u2479_o),
    .b(_al_u2481_o),
    .c(_al_u2483_o),
    .d(_al_u2485_o),
    .e(_al_u2487_o),
    .o(_al_u2488_o));
  AL_MAP_LUT5 #(
    .EQN("(~B*~(E@C)*~(D*~A))"),
    .INIT(32'h20300203))
    _al_u2489 (
    .a(\PWM9/FreCnt [19]),
    .b(\PWM9/FreCnt [26]),
    .c(\PWM9/FreCnt [4]),
    .d(\PWM9/FreCntr [20]),
    .e(\PWM9/FreCntr [5]),
    .o(_al_u2489_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u249 (
    .a(\PWM1/pnumr [11]),
    .b(pnum1[11]),
    .c(pnum1[32]),
    .d(pwm_start_stop[17]),
    .o(\PWM1/n23 [11]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u2490 (
    .a(_al_u2489_o),
    .b(\PWM9/FreCnt [24]),
    .c(\PWM9/FreCnt [6]),
    .d(\PWM9/FreCntr [25]),
    .e(\PWM9/FreCntr [7]),
    .o(_al_u2490_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u2491 (
    .a(\PWM9/FreCnt [0]),
    .b(\PWM9/FreCnt [11]),
    .c(\PWM9/FreCntr [1]),
    .d(\PWM9/FreCntr [12]),
    .o(_al_u2491_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u2492 (
    .a(_al_u2491_o),
    .b(\PWM9/FreCnt [2]),
    .c(\PWM9/FreCntr [3]),
    .o(_al_u2492_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u2493 (
    .a(\PWM9/FreCnt [7]),
    .b(\PWM9/FreCnt [8]),
    .c(\PWM9/FreCntr [8]),
    .d(\PWM9/FreCntr [9]),
    .o(_al_u2493_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*C)*~(~D*B))"),
    .INIT(32'haa220a02))
    _al_u2494 (
    .a(_al_u2493_o),
    .b(\PWM9/FreCnt [17]),
    .c(\PWM9/FreCnt [21]),
    .d(\PWM9/FreCntr [18]),
    .e(\PWM9/FreCntr [22]),
    .o(_al_u2494_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2495 (
    .a(\PWM9/FreCnt [15]),
    .b(\PWM9/FreCntr [16]),
    .o(_al_u2495_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(E@C)*~(~D*B))"),
    .INIT(32'h50100501))
    _al_u2496 (
    .a(_al_u2495_o),
    .b(\PWM9/FreCnt [19]),
    .c(\PWM9/FreCnt [25]),
    .d(\PWM9/FreCntr [20]),
    .e(\PWM9/FreCntr [26]),
    .o(_al_u2496_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    _al_u2497 (
    .a(_al_u2488_o),
    .b(_al_u2490_o),
    .c(_al_u2492_o),
    .d(_al_u2494_o),
    .e(_al_u2496_o),
    .o(_al_u2497_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2498 (
    .a(_al_u2497_o),
    .b(pwm_state_read[9]),
    .o(\PWM9/u14_sel_is_1_o ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2499 (
    .a(\PWMA/n0_lutinv ),
    .b(pwm_state_read[10]),
    .o(\PWMA/n24 ));
  EF2_PHY_PAD #(
    //.LOCATION("P48"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u25 (
    .do({open_n800,open_n801,open_n802,dir_pad[13]}),
    .opad(dir[13]));  // CPLD_SOC_AHB_TOP.v(7)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u250 (
    .a(\PWM1/pnumr [10]),
    .b(pnum1[10]),
    .c(pnum1[32]),
    .d(pwm_start_stop[17]),
    .o(\PWM1/n23 [10]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u2500 (
    .a(pnumcntA[18]),
    .b(pnumcntA[19]),
    .c(pnumcntA[1]),
    .d(pnumcntA[20]),
    .o(_al_u2500_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u2501 (
    .a(_al_u2500_o),
    .b(pnumcntA[21]),
    .c(pnumcntA[22]),
    .d(pnumcntA[23]),
    .e(pnumcntA[2]),
    .o(_al_u2501_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u2502 (
    .a(_al_u2501_o),
    .b(pnumcntA[6]),
    .c(pnumcntA[7]),
    .d(pnumcntA[8]),
    .e(pnumcntA[9]),
    .o(_al_u2502_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u2503 (
    .a(pnumcntA[10]),
    .b(pnumcntA[11]),
    .c(pnumcntA[12]),
    .d(pnumcntA[13]),
    .o(_al_u2503_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u2504 (
    .a(_al_u2503_o),
    .b(pnumcntA[14]),
    .c(pnumcntA[15]),
    .d(pnumcntA[16]),
    .e(pnumcntA[17]),
    .o(_al_u2504_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u2505 (
    .a(pnumcntA[3]),
    .b(pnumcntA[4]),
    .c(pnumcntA[5]),
    .o(_al_u2505_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u2506 (
    .a(_al_u2502_o),
    .b(_al_u2504_o),
    .c(_al_u2505_o),
    .d(pnumcntA[0]),
    .o(\PWMA/n25_neg_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2507 (
    .a(\PWMA/n24 ),
    .b(\PWMA/n25_neg_lutinv ),
    .c(\PWMA/n26 [9]),
    .d(\PWMA/pnumr [9]),
    .o(_al_u2507_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2508 (
    .a(_al_u2507_o),
    .b(\PWMA/n24 ),
    .c(pnumcntA[9]),
    .d(\PWMA/pnumr [9]),
    .e(pwm_start_stop[26]),
    .o(\PWMA/n31 [9]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2509 (
    .a(\PWMA/n24 ),
    .b(\PWMA/n25_neg_lutinv ),
    .c(\PWMA/n26 [8]),
    .d(\PWMA/pnumr [8]),
    .o(_al_u2509_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u251 (
    .a(\PWM1/pnumr [1]),
    .b(pnum1[1]),
    .c(pnum1[32]),
    .d(pwm_start_stop[17]),
    .o(\PWM1/n23 [1]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2510 (
    .a(_al_u2509_o),
    .b(\PWMA/n24 ),
    .c(pnumcntA[8]),
    .d(\PWMA/pnumr [8]),
    .e(pwm_start_stop[26]),
    .o(\PWMA/n31 [8]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2511 (
    .a(\PWMA/n24 ),
    .b(\PWMA/n25_neg_lutinv ),
    .c(\PWMA/n26 [7]),
    .d(\PWMA/pnumr [7]),
    .o(_al_u2511_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2512 (
    .a(_al_u2511_o),
    .b(\PWMA/n24 ),
    .c(pnumcntA[7]),
    .d(\PWMA/pnumr [7]),
    .e(pwm_start_stop[26]),
    .o(\PWMA/n31 [7]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2513 (
    .a(\PWMA/n24 ),
    .b(\PWMA/n25_neg_lutinv ),
    .c(\PWMA/n26 [6]),
    .d(\PWMA/pnumr [6]),
    .o(_al_u2513_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2514 (
    .a(_al_u2513_o),
    .b(\PWMA/n24 ),
    .c(pnumcntA[6]),
    .d(\PWMA/pnumr [6]),
    .e(pwm_start_stop[26]),
    .o(\PWMA/n31 [6]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2515 (
    .a(\PWMA/n24 ),
    .b(\PWMA/n25_neg_lutinv ),
    .c(\PWMA/n26 [5]),
    .d(\PWMA/pnumr [5]),
    .o(_al_u2515_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2516 (
    .a(_al_u2515_o),
    .b(\PWMA/n24 ),
    .c(pnumcntA[5]),
    .d(\PWMA/pnumr [5]),
    .e(pwm_start_stop[26]),
    .o(\PWMA/n31 [5]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2517 (
    .a(\PWMA/n24 ),
    .b(\PWMA/n25_neg_lutinv ),
    .c(\PWMA/n26 [4]),
    .d(\PWMA/pnumr [4]),
    .o(_al_u2517_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2518 (
    .a(_al_u2517_o),
    .b(\PWMA/n24 ),
    .c(pnumcntA[4]),
    .d(\PWMA/pnumr [4]),
    .e(pwm_start_stop[26]),
    .o(\PWMA/n31 [4]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2519 (
    .a(\PWMA/n24 ),
    .b(\PWMA/n25_neg_lutinv ),
    .c(\PWMA/n26 [3]),
    .d(\PWMA/pnumr [3]),
    .o(_al_u2519_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u252 (
    .a(\PWM1/pnumr [0]),
    .b(pnum1[0]),
    .c(pnum1[32]),
    .d(pwm_start_stop[17]),
    .o(\PWM1/n23 [0]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2520 (
    .a(_al_u2519_o),
    .b(\PWMA/n24 ),
    .c(pnumcntA[3]),
    .d(\PWMA/pnumr [3]),
    .e(pwm_start_stop[26]),
    .o(\PWMA/n31 [3]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2521 (
    .a(\PWMA/n24 ),
    .b(\PWMA/n25_neg_lutinv ),
    .c(\PWMA/n26 [23]),
    .d(\PWMA/pnumr [23]),
    .o(_al_u2521_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2522 (
    .a(_al_u2521_o),
    .b(\PWMA/n24 ),
    .c(pnumcntA[23]),
    .d(\PWMA/pnumr [23]),
    .e(pwm_start_stop[26]),
    .o(\PWMA/n31 [23]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2523 (
    .a(\PWMA/n24 ),
    .b(\PWMA/n25_neg_lutinv ),
    .c(\PWMA/n26 [22]),
    .d(\PWMA/pnumr [22]),
    .o(_al_u2523_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2524 (
    .a(_al_u2523_o),
    .b(\PWMA/n24 ),
    .c(pnumcntA[22]),
    .d(\PWMA/pnumr [22]),
    .e(pwm_start_stop[26]),
    .o(\PWMA/n31 [22]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2525 (
    .a(\PWMA/n24 ),
    .b(\PWMA/n25_neg_lutinv ),
    .c(\PWMA/n26 [21]),
    .d(\PWMA/pnumr [21]),
    .o(_al_u2525_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2526 (
    .a(_al_u2525_o),
    .b(\PWMA/n24 ),
    .c(pnumcntA[21]),
    .d(\PWMA/pnumr [21]),
    .e(pwm_start_stop[26]),
    .o(\PWMA/n31 [21]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2527 (
    .a(\PWMA/n24 ),
    .b(\PWMA/n25_neg_lutinv ),
    .c(\PWMA/n26 [20]),
    .d(\PWMA/pnumr [20]),
    .o(_al_u2527_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2528 (
    .a(_al_u2527_o),
    .b(\PWMA/n24 ),
    .c(pnumcntA[20]),
    .d(\PWMA/pnumr [20]),
    .e(pwm_start_stop[26]),
    .o(\PWMA/n31 [20]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2529 (
    .a(\PWMA/n24 ),
    .b(\PWMA/n25_neg_lutinv ),
    .c(\PWMA/n26 [2]),
    .d(\PWMA/pnumr [2]),
    .o(_al_u2529_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u253 (
    .a(\PWM2/pnumr [9]),
    .b(pnum2[32]),
    .c(pnum2[9]),
    .d(pwm_start_stop[18]),
    .o(\PWM2/n23 [9]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2530 (
    .a(_al_u2529_o),
    .b(\PWMA/n24 ),
    .c(pnumcntA[2]),
    .d(\PWMA/pnumr [2]),
    .e(pwm_start_stop[26]),
    .o(\PWMA/n31 [2]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2531 (
    .a(\PWMA/n24 ),
    .b(\PWMA/n25_neg_lutinv ),
    .c(\PWMA/n26 [19]),
    .d(\PWMA/pnumr [19]),
    .o(_al_u2531_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2532 (
    .a(_al_u2531_o),
    .b(\PWMA/n24 ),
    .c(pnumcntA[19]),
    .d(\PWMA/pnumr [19]),
    .e(pwm_start_stop[26]),
    .o(\PWMA/n31 [19]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2533 (
    .a(\PWMA/n24 ),
    .b(\PWMA/n25_neg_lutinv ),
    .c(\PWMA/n26 [18]),
    .d(\PWMA/pnumr [18]),
    .o(_al_u2533_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2534 (
    .a(_al_u2533_o),
    .b(\PWMA/n24 ),
    .c(pnumcntA[18]),
    .d(\PWMA/pnumr [18]),
    .e(pwm_start_stop[26]),
    .o(\PWMA/n31 [18]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2535 (
    .a(\PWMA/n24 ),
    .b(\PWMA/n25_neg_lutinv ),
    .c(\PWMA/n26 [17]),
    .d(\PWMA/pnumr [17]),
    .o(_al_u2535_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2536 (
    .a(_al_u2535_o),
    .b(\PWMA/n24 ),
    .c(pnumcntA[17]),
    .d(\PWMA/pnumr [17]),
    .e(pwm_start_stop[26]),
    .o(\PWMA/n31 [17]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2537 (
    .a(\PWMA/n24 ),
    .b(\PWMA/n25_neg_lutinv ),
    .c(\PWMA/n26 [16]),
    .d(\PWMA/pnumr [16]),
    .o(_al_u2537_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2538 (
    .a(_al_u2537_o),
    .b(\PWMA/n24 ),
    .c(pnumcntA[16]),
    .d(\PWMA/pnumr [16]),
    .e(pwm_start_stop[26]),
    .o(\PWMA/n31 [16]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2539 (
    .a(\PWMA/n24 ),
    .b(\PWMA/n25_neg_lutinv ),
    .c(\PWMA/n26 [15]),
    .d(\PWMA/pnumr [15]),
    .o(_al_u2539_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u254 (
    .a(\PWM2/pnumr [8]),
    .b(pnum2[32]),
    .c(pnum2[8]),
    .d(pwm_start_stop[18]),
    .o(\PWM2/n23 [8]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2540 (
    .a(_al_u2539_o),
    .b(\PWMA/n24 ),
    .c(pnumcntA[15]),
    .d(\PWMA/pnumr [15]),
    .e(pwm_start_stop[26]),
    .o(\PWMA/n31 [15]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2541 (
    .a(\PWMA/n24 ),
    .b(\PWMA/n25_neg_lutinv ),
    .c(\PWMA/n26 [14]),
    .d(\PWMA/pnumr [14]),
    .o(_al_u2541_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2542 (
    .a(_al_u2541_o),
    .b(\PWMA/n24 ),
    .c(pnumcntA[14]),
    .d(\PWMA/pnumr [14]),
    .e(pwm_start_stop[26]),
    .o(\PWMA/n31 [14]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2543 (
    .a(\PWMA/n24 ),
    .b(\PWMA/n25_neg_lutinv ),
    .c(\PWMA/n26 [13]),
    .d(\PWMA/pnumr [13]),
    .o(_al_u2543_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2544 (
    .a(_al_u2543_o),
    .b(\PWMA/n24 ),
    .c(pnumcntA[13]),
    .d(\PWMA/pnumr [13]),
    .e(pwm_start_stop[26]),
    .o(\PWMA/n31 [13]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2545 (
    .a(\PWMA/n24 ),
    .b(\PWMA/n25_neg_lutinv ),
    .c(\PWMA/n26 [12]),
    .d(\PWMA/pnumr [12]),
    .o(_al_u2545_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2546 (
    .a(_al_u2545_o),
    .b(\PWMA/n24 ),
    .c(pnumcntA[12]),
    .d(\PWMA/pnumr [12]),
    .e(pwm_start_stop[26]),
    .o(\PWMA/n31 [12]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2547 (
    .a(\PWMA/n24 ),
    .b(\PWMA/n25_neg_lutinv ),
    .c(\PWMA/n26 [11]),
    .d(\PWMA/pnumr [11]),
    .o(_al_u2547_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2548 (
    .a(_al_u2547_o),
    .b(\PWMA/n24 ),
    .c(pnumcntA[11]),
    .d(\PWMA/pnumr [11]),
    .e(pwm_start_stop[26]),
    .o(\PWMA/n31 [11]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2549 (
    .a(\PWMA/n24 ),
    .b(\PWMA/n25_neg_lutinv ),
    .c(\PWMA/n26 [10]),
    .d(\PWMA/pnumr [10]),
    .o(_al_u2549_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u255 (
    .a(\PWM2/pnumr [7]),
    .b(pnum2[32]),
    .c(pnum2[7]),
    .d(pwm_start_stop[18]),
    .o(\PWM2/n23 [7]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2550 (
    .a(_al_u2549_o),
    .b(\PWMA/n24 ),
    .c(pnumcntA[10]),
    .d(\PWMA/pnumr [10]),
    .e(pwm_start_stop[26]),
    .o(\PWMA/n31 [10]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2551 (
    .a(\PWMA/n24 ),
    .b(\PWMA/n25_neg_lutinv ),
    .c(\PWMA/n26 [1]),
    .d(\PWMA/pnumr [1]),
    .o(_al_u2551_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2552 (
    .a(_al_u2551_o),
    .b(\PWMA/n24 ),
    .c(pnumcntA[1]),
    .d(\PWMA/pnumr [1]),
    .e(pwm_start_stop[26]),
    .o(\PWMA/n31 [1]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2553 (
    .a(\PWMA/n24 ),
    .b(\PWMA/n25_neg_lutinv ),
    .c(\PWMA/n26 [0]),
    .d(\PWMA/pnumr [0]),
    .o(_al_u2553_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2554 (
    .a(_al_u2553_o),
    .b(\PWMA/n24 ),
    .c(pnumcntA[0]),
    .d(\PWMA/pnumr [0]),
    .e(pwm_start_stop[26]),
    .o(\PWMA/n31 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u2555 (
    .a(\PWMA/FreCnt [10]),
    .b(\PWMA/FreCnt [15]),
    .c(\PWMA/FreCntr [11]),
    .d(\PWMA/FreCntr [16]),
    .o(_al_u2555_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*~C)*~(~E*B))"),
    .INIT(32'ha0aa2022))
    _al_u2556 (
    .a(_al_u2555_o),
    .b(\PWMA/FreCnt [7]),
    .c(\PWMA/FreCnt [9]),
    .d(\PWMA/FreCntr [10]),
    .e(\PWMA/FreCntr [8]),
    .o(_al_u2556_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*C)*~(D@B))"),
    .INIT(32'h88220802))
    _al_u2557 (
    .a(_al_u2556_o),
    .b(\PWMA/FreCnt [2]),
    .c(\PWMA/FreCnt [8]),
    .d(\PWMA/FreCntr [3]),
    .e(\PWMA/FreCntr [9]),
    .o(_al_u2557_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2558 (
    .a(\PWMA/FreCnt [9]),
    .b(\PWMA/FreCntr [10]),
    .o(_al_u2558_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(~E*C)*~(D@B))"),
    .INIT(32'h44110401))
    _al_u2559 (
    .a(_al_u2558_o),
    .b(\PWMA/FreCnt [24]),
    .c(\PWMA/FreCnt [3]),
    .d(\PWMA/FreCntr [25]),
    .e(\PWMA/FreCntr [4]),
    .o(_al_u2559_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u256 (
    .a(\PWM2/pnumr [6]),
    .b(pnum2[32]),
    .c(pnum2[6]),
    .d(pwm_start_stop[18]),
    .o(\PWM2/n23 [6]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u2560 (
    .a(\PWMA/FreCnt [23]),
    .b(\PWMA/FreCnt [3]),
    .c(\PWMA/FreCntr [24]),
    .d(\PWMA/FreCntr [4]),
    .o(_al_u2560_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u2561 (
    .a(_al_u2557_o),
    .b(_al_u2559_o),
    .c(_al_u2560_o),
    .d(\PWMA/FreCnt [1]),
    .e(\PWMA/FreCntr [2]),
    .o(_al_u2561_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u2562 (
    .a(\PWMA/FreCnt [15]),
    .b(\PWMA/FreCnt [5]),
    .c(\PWMA/FreCntr [16]),
    .d(\PWMA/FreCntr [6]),
    .o(_al_u2562_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*C)*~(~D*B))"),
    .INIT(32'haa220a02))
    _al_u2563 (
    .a(_al_u2562_o),
    .b(\PWMA/FreCnt [12]),
    .c(\PWMA/FreCnt [19]),
    .d(\PWMA/FreCntr [13]),
    .e(\PWMA/FreCntr [20]),
    .o(_al_u2563_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u2564 (
    .a(_al_u2563_o),
    .b(\PWMA/FreCnt [0]),
    .c(\PWMA/FreCnt [4]),
    .d(\PWMA/FreCntr [1]),
    .e(\PWMA/FreCntr [5]),
    .o(_al_u2564_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u2565 (
    .a(\PWMA/FreCnt [17]),
    .b(\PWMA/FreCnt [19]),
    .c(\PWMA/FreCntr [18]),
    .d(\PWMA/FreCntr [20]),
    .o(_al_u2565_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*C)*~(D*~B))"),
    .INIT(32'h88aa080a))
    _al_u2566 (
    .a(_al_u2565_o),
    .b(\PWMA/FreCnt [12]),
    .c(\PWMA/FreCnt [23]),
    .d(\PWMA/FreCntr [13]),
    .e(\PWMA/FreCntr [24]),
    .o(_al_u2566_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u2567 (
    .a(\PWMA/FreCnt [10]),
    .b(\PWMA/FreCnt [5]),
    .c(\PWMA/FreCntr [11]),
    .d(\PWMA/FreCntr [6]),
    .o(_al_u2567_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u2568 (
    .a(_al_u2564_o),
    .b(_al_u2566_o),
    .c(_al_u2567_o),
    .d(\PWMA/FreCnt [16]),
    .e(\PWMA/FreCntr [17]),
    .o(_al_u2568_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u2569 (
    .a(\PWMA/FreCnt [14]),
    .b(\PWMA/FreCnt [21]),
    .c(\PWMA/FreCntr [15]),
    .d(\PWMA/FreCntr [22]),
    .o(_al_u2569_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u257 (
    .a(\PWM2/pnumr [5]),
    .b(pnum2[32]),
    .c(pnum2[5]),
    .d(pwm_start_stop[18]),
    .o(\PWM2/n23 [5]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u2570 (
    .a(_al_u2569_o),
    .b(\PWMA/FreCnt [20]),
    .c(\PWMA/FreCntr [21]),
    .o(_al_u2570_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u2571 (
    .a(\PWMA/FreCnt [11]),
    .b(\PWMA/FreCnt [6]),
    .c(\PWMA/FreCntr [12]),
    .d(\PWMA/FreCntr [7]),
    .o(_al_u2571_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u2572 (
    .a(_al_u2571_o),
    .b(\PWMA/FreCnt [18]),
    .c(\PWMA/FreCnt [22]),
    .d(\PWMA/FreCntr [19]),
    .e(\PWMA/FreCntr [23]),
    .o(_al_u2572_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u2573 (
    .a(\PWMA/FreCnt [17]),
    .b(\PWMA/FreCnt [8]),
    .c(\PWMA/FreCntr [18]),
    .d(\PWMA/FreCntr [9]),
    .o(_al_u2573_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*~C)*~(D*~B))"),
    .INIT(32'h80a088aa))
    _al_u2574 (
    .a(_al_u2573_o),
    .b(\PWMA/FreCnt [13]),
    .c(\PWMA/FreCnt [7]),
    .d(\PWMA/FreCntr [14]),
    .e(\PWMA/FreCntr [8]),
    .o(_al_u2574_o));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(E@B)*~(~D*A))"),
    .INIT(32'h0c040301))
    _al_u2575 (
    .a(\PWMA/FreCnt [13]),
    .b(\PWMA/FreCnt [25]),
    .c(\PWMA/FreCnt [26]),
    .d(\PWMA/FreCntr [14]),
    .e(\PWMA/FreCntr [26]),
    .o(_al_u2575_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u2576 (
    .a(_al_u2570_o),
    .b(_al_u2572_o),
    .c(_al_u2574_o),
    .d(_al_u2575_o),
    .o(_al_u2576_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*A))"),
    .INIT(16'h7f00))
    _al_u2577 (
    .a(_al_u2561_o),
    .b(_al_u2568_o),
    .c(_al_u2576_o),
    .d(pwm_state_read[10]),
    .o(\PWMA/u14_sel_is_1_o ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2578 (
    .a(\PWMB/n0_lutinv ),
    .b(pwm_state_read[11]),
    .o(\PWMB/n24 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u2579 (
    .a(pnumcntB[18]),
    .b(pnumcntB[19]),
    .c(pnumcntB[1]),
    .d(pnumcntB[20]),
    .o(_al_u2579_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u258 (
    .a(\PWM2/pnumr [4]),
    .b(pnum2[32]),
    .c(pnum2[4]),
    .d(pwm_start_stop[18]),
    .o(\PWM2/n23 [4]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u2580 (
    .a(_al_u2579_o),
    .b(pnumcntB[21]),
    .c(pnumcntB[22]),
    .d(pnumcntB[23]),
    .e(pnumcntB[2]),
    .o(_al_u2580_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u2581 (
    .a(_al_u2580_o),
    .b(pnumcntB[6]),
    .c(pnumcntB[7]),
    .d(pnumcntB[8]),
    .e(pnumcntB[9]),
    .o(_al_u2581_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u2582 (
    .a(pnumcntB[10]),
    .b(pnumcntB[11]),
    .c(pnumcntB[12]),
    .d(pnumcntB[13]),
    .o(_al_u2582_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u2583 (
    .a(_al_u2582_o),
    .b(pnumcntB[14]),
    .c(pnumcntB[15]),
    .d(pnumcntB[16]),
    .e(pnumcntB[17]),
    .o(_al_u2583_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u2584 (
    .a(pnumcntB[3]),
    .b(pnumcntB[4]),
    .c(pnumcntB[5]),
    .o(_al_u2584_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u2585 (
    .a(_al_u2581_o),
    .b(_al_u2583_o),
    .c(_al_u2584_o),
    .d(pnumcntB[0]),
    .o(\PWMB/n25_neg_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2586 (
    .a(\PWMB/n24 ),
    .b(\PWMB/n25_neg_lutinv ),
    .c(\PWMB/n26 [9]),
    .d(\PWMB/pnumr [9]),
    .o(_al_u2586_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2587 (
    .a(_al_u2586_o),
    .b(\PWMB/n24 ),
    .c(pnumcntB[9]),
    .d(\PWMB/pnumr [9]),
    .e(pwm_start_stop[27]),
    .o(\PWMB/n31 [9]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2588 (
    .a(\PWMB/n24 ),
    .b(\PWMB/n25_neg_lutinv ),
    .c(\PWMB/n26 [8]),
    .d(\PWMB/pnumr [8]),
    .o(_al_u2588_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2589 (
    .a(_al_u2588_o),
    .b(\PWMB/n24 ),
    .c(pnumcntB[8]),
    .d(\PWMB/pnumr [8]),
    .e(pwm_start_stop[27]),
    .o(\PWMB/n31 [8]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u259 (
    .a(\PWM2/pnumr [31]),
    .b(pnum2[31]),
    .c(pnum2[32]),
    .d(pwm_start_stop[18]),
    .o(\PWM2/n23 [31]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2590 (
    .a(\PWMB/n24 ),
    .b(\PWMB/n25_neg_lutinv ),
    .c(\PWMB/n26 [7]),
    .d(\PWMB/pnumr [7]),
    .o(_al_u2590_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2591 (
    .a(_al_u2590_o),
    .b(\PWMB/n24 ),
    .c(pnumcntB[7]),
    .d(\PWMB/pnumr [7]),
    .e(pwm_start_stop[27]),
    .o(\PWMB/n31 [7]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2592 (
    .a(\PWMB/n24 ),
    .b(\PWMB/n25_neg_lutinv ),
    .c(\PWMB/n26 [6]),
    .d(\PWMB/pnumr [6]),
    .o(_al_u2592_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2593 (
    .a(_al_u2592_o),
    .b(\PWMB/n24 ),
    .c(pnumcntB[6]),
    .d(\PWMB/pnumr [6]),
    .e(pwm_start_stop[27]),
    .o(\PWMB/n31 [6]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2594 (
    .a(\PWMB/n24 ),
    .b(\PWMB/n25_neg_lutinv ),
    .c(\PWMB/n26 [5]),
    .d(\PWMB/pnumr [5]),
    .o(_al_u2594_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2595 (
    .a(_al_u2594_o),
    .b(\PWMB/n24 ),
    .c(pnumcntB[5]),
    .d(\PWMB/pnumr [5]),
    .e(pwm_start_stop[27]),
    .o(\PWMB/n31 [5]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2596 (
    .a(\PWMB/n24 ),
    .b(\PWMB/n25_neg_lutinv ),
    .c(\PWMB/n26 [4]),
    .d(\PWMB/pnumr [4]),
    .o(_al_u2596_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2597 (
    .a(_al_u2596_o),
    .b(\PWMB/n24 ),
    .c(pnumcntB[4]),
    .d(\PWMB/pnumr [4]),
    .e(pwm_start_stop[27]),
    .o(\PWMB/n31 [4]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2598 (
    .a(\PWMB/n24 ),
    .b(\PWMB/n25_neg_lutinv ),
    .c(\PWMB/n26 [3]),
    .d(\PWMB/pnumr [3]),
    .o(_al_u2598_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2599 (
    .a(_al_u2598_o),
    .b(\PWMB/n24 ),
    .c(pnumcntB[3]),
    .d(\PWMB/pnumr [3]),
    .e(pwm_start_stop[27]),
    .o(\PWMB/n31 [3]));
  EF2_PHY_PAD #(
    //.LOCATION("P45"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u26 (
    .do({open_n823,open_n824,open_n825,dir_pad[12]}),
    .opad(dir[12]));  // CPLD_SOC_AHB_TOP.v(7)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u260 (
    .a(\PWM2/pnumr [30]),
    .b(pnum2[30]),
    .c(pnum2[32]),
    .d(pwm_start_stop[18]),
    .o(\PWM2/n23 [30]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2600 (
    .a(\PWMB/n24 ),
    .b(\PWMB/n25_neg_lutinv ),
    .c(\PWMB/n26 [23]),
    .d(\PWMB/pnumr [23]),
    .o(_al_u2600_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2601 (
    .a(_al_u2600_o),
    .b(\PWMB/n24 ),
    .c(pnumcntB[23]),
    .d(\PWMB/pnumr [23]),
    .e(pwm_start_stop[27]),
    .o(\PWMB/n31 [23]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2602 (
    .a(\PWMB/n24 ),
    .b(\PWMB/n25_neg_lutinv ),
    .c(\PWMB/n26 [22]),
    .d(\PWMB/pnumr [22]),
    .o(_al_u2602_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2603 (
    .a(_al_u2602_o),
    .b(\PWMB/n24 ),
    .c(pnumcntB[22]),
    .d(\PWMB/pnumr [22]),
    .e(pwm_start_stop[27]),
    .o(\PWMB/n31 [22]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2604 (
    .a(\PWMB/n24 ),
    .b(\PWMB/n25_neg_lutinv ),
    .c(\PWMB/n26 [21]),
    .d(\PWMB/pnumr [21]),
    .o(_al_u2604_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2605 (
    .a(_al_u2604_o),
    .b(\PWMB/n24 ),
    .c(pnumcntB[21]),
    .d(\PWMB/pnumr [21]),
    .e(pwm_start_stop[27]),
    .o(\PWMB/n31 [21]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2606 (
    .a(\PWMB/n24 ),
    .b(\PWMB/n25_neg_lutinv ),
    .c(\PWMB/n26 [20]),
    .d(\PWMB/pnumr [20]),
    .o(_al_u2606_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2607 (
    .a(_al_u2606_o),
    .b(\PWMB/n24 ),
    .c(pnumcntB[20]),
    .d(\PWMB/pnumr [20]),
    .e(pwm_start_stop[27]),
    .o(\PWMB/n31 [20]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2608 (
    .a(\PWMB/n24 ),
    .b(\PWMB/n25_neg_lutinv ),
    .c(\PWMB/n26 [2]),
    .d(\PWMB/pnumr [2]),
    .o(_al_u2608_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2609 (
    .a(_al_u2608_o),
    .b(\PWMB/n24 ),
    .c(pnumcntB[2]),
    .d(\PWMB/pnumr [2]),
    .e(pwm_start_stop[27]),
    .o(\PWMB/n31 [2]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u261 (
    .a(\PWM2/pnumr [3]),
    .b(pnum2[3]),
    .c(pnum2[32]),
    .d(pwm_start_stop[18]),
    .o(\PWM2/n23 [3]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2610 (
    .a(\PWMB/n24 ),
    .b(\PWMB/n25_neg_lutinv ),
    .c(\PWMB/n26 [19]),
    .d(\PWMB/pnumr [19]),
    .o(_al_u2610_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2611 (
    .a(_al_u2610_o),
    .b(\PWMB/n24 ),
    .c(pnumcntB[19]),
    .d(\PWMB/pnumr [19]),
    .e(pwm_start_stop[27]),
    .o(\PWMB/n31 [19]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2612 (
    .a(\PWMB/n24 ),
    .b(\PWMB/n25_neg_lutinv ),
    .c(\PWMB/n26 [18]),
    .d(\PWMB/pnumr [18]),
    .o(_al_u2612_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2613 (
    .a(_al_u2612_o),
    .b(\PWMB/n24 ),
    .c(pnumcntB[18]),
    .d(\PWMB/pnumr [18]),
    .e(pwm_start_stop[27]),
    .o(\PWMB/n31 [18]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2614 (
    .a(\PWMB/n24 ),
    .b(\PWMB/n25_neg_lutinv ),
    .c(\PWMB/n26 [17]),
    .d(\PWMB/pnumr [17]),
    .o(_al_u2614_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2615 (
    .a(_al_u2614_o),
    .b(\PWMB/n24 ),
    .c(pnumcntB[17]),
    .d(\PWMB/pnumr [17]),
    .e(pwm_start_stop[27]),
    .o(\PWMB/n31 [17]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2616 (
    .a(\PWMB/n24 ),
    .b(\PWMB/n25_neg_lutinv ),
    .c(\PWMB/n26 [16]),
    .d(\PWMB/pnumr [16]),
    .o(_al_u2616_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2617 (
    .a(_al_u2616_o),
    .b(\PWMB/n24 ),
    .c(pnumcntB[16]),
    .d(\PWMB/pnumr [16]),
    .e(pwm_start_stop[27]),
    .o(\PWMB/n31 [16]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2618 (
    .a(\PWMB/n24 ),
    .b(\PWMB/n25_neg_lutinv ),
    .c(\PWMB/n26 [15]),
    .d(\PWMB/pnumr [15]),
    .o(_al_u2618_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2619 (
    .a(_al_u2618_o),
    .b(\PWMB/n24 ),
    .c(pnumcntB[15]),
    .d(\PWMB/pnumr [15]),
    .e(pwm_start_stop[27]),
    .o(\PWMB/n31 [15]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u262 (
    .a(\PWM2/pnumr [29]),
    .b(pnum2[29]),
    .c(pnum2[32]),
    .d(pwm_start_stop[18]),
    .o(\PWM2/n23 [29]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2620 (
    .a(\PWMB/n24 ),
    .b(\PWMB/n25_neg_lutinv ),
    .c(\PWMB/n26 [14]),
    .d(\PWMB/pnumr [14]),
    .o(_al_u2620_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2621 (
    .a(_al_u2620_o),
    .b(\PWMB/n24 ),
    .c(pnumcntB[14]),
    .d(\PWMB/pnumr [14]),
    .e(pwm_start_stop[27]),
    .o(\PWMB/n31 [14]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2622 (
    .a(\PWMB/n24 ),
    .b(\PWMB/n25_neg_lutinv ),
    .c(\PWMB/n26 [13]),
    .d(\PWMB/pnumr [13]),
    .o(_al_u2622_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2623 (
    .a(_al_u2622_o),
    .b(\PWMB/n24 ),
    .c(pnumcntB[13]),
    .d(\PWMB/pnumr [13]),
    .e(pwm_start_stop[27]),
    .o(\PWMB/n31 [13]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2624 (
    .a(\PWMB/n24 ),
    .b(\PWMB/n25_neg_lutinv ),
    .c(\PWMB/n26 [12]),
    .d(\PWMB/pnumr [12]),
    .o(_al_u2624_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2625 (
    .a(_al_u2624_o),
    .b(\PWMB/n24 ),
    .c(pnumcntB[12]),
    .d(\PWMB/pnumr [12]),
    .e(pwm_start_stop[27]),
    .o(\PWMB/n31 [12]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2626 (
    .a(\PWMB/n24 ),
    .b(\PWMB/n25_neg_lutinv ),
    .c(\PWMB/n26 [11]),
    .d(\PWMB/pnumr [11]),
    .o(_al_u2626_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2627 (
    .a(_al_u2626_o),
    .b(\PWMB/n24 ),
    .c(pnumcntB[11]),
    .d(\PWMB/pnumr [11]),
    .e(pwm_start_stop[27]),
    .o(\PWMB/n31 [11]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2628 (
    .a(\PWMB/n24 ),
    .b(\PWMB/n25_neg_lutinv ),
    .c(\PWMB/n26 [10]),
    .d(\PWMB/pnumr [10]),
    .o(_al_u2628_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2629 (
    .a(_al_u2628_o),
    .b(\PWMB/n24 ),
    .c(pnumcntB[10]),
    .d(\PWMB/pnumr [10]),
    .e(pwm_start_stop[27]),
    .o(\PWMB/n31 [10]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u263 (
    .a(\PWM2/pnumr [28]),
    .b(pnum2[28]),
    .c(pnum2[32]),
    .d(pwm_start_stop[18]),
    .o(\PWM2/n23 [28]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2630 (
    .a(\PWMB/n24 ),
    .b(\PWMB/n25_neg_lutinv ),
    .c(\PWMB/n26 [1]),
    .d(\PWMB/pnumr [1]),
    .o(_al_u2630_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2631 (
    .a(_al_u2630_o),
    .b(\PWMB/n24 ),
    .c(pnumcntB[1]),
    .d(\PWMB/pnumr [1]),
    .e(pwm_start_stop[27]),
    .o(\PWMB/n31 [1]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2632 (
    .a(\PWMB/n24 ),
    .b(\PWMB/n25_neg_lutinv ),
    .c(\PWMB/n26 [0]),
    .d(\PWMB/pnumr [0]),
    .o(_al_u2632_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2633 (
    .a(_al_u2632_o),
    .b(\PWMB/n24 ),
    .c(pnumcntB[0]),
    .d(\PWMB/pnumr [0]),
    .e(pwm_start_stop[27]),
    .o(\PWMB/n31 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u2634 (
    .a(\PWMB/FreCnt [19]),
    .b(\PWMB/FreCnt [8]),
    .c(\PWMB/FreCntr [20]),
    .d(\PWMB/FreCntr [9]),
    .o(_al_u2634_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*~C)*~(D*~B))"),
    .INIT(32'h80a088aa))
    _al_u2635 (
    .a(_al_u2634_o),
    .b(\PWMB/FreCnt [17]),
    .c(\PWMB/FreCnt [3]),
    .d(\PWMB/FreCntr [18]),
    .e(\PWMB/FreCntr [4]),
    .o(_al_u2635_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u2636 (
    .a(\PWMB/FreCnt [21]),
    .b(\PWMB/FreCnt [5]),
    .c(\PWMB/FreCntr [22]),
    .d(\PWMB/FreCntr [6]),
    .o(_al_u2636_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(~D*C))"),
    .INIT(16'h8808))
    _al_u2637 (
    .a(_al_u2635_o),
    .b(_al_u2636_o),
    .c(\PWMB/FreCnt [10]),
    .d(\PWMB/FreCntr [11]),
    .o(_al_u2637_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u2638 (
    .a(\PWMB/FreCnt [25]),
    .b(\PWMB/FreCnt [7]),
    .c(\PWMB/FreCntr [26]),
    .d(\PWMB/FreCntr [8]),
    .o(_al_u2638_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*C)*~(D*~B))"),
    .INIT(32'h88aa080a))
    _al_u2639 (
    .a(_al_u2638_o),
    .b(\PWMB/FreCnt [10]),
    .c(\PWMB/FreCnt [3]),
    .d(\PWMB/FreCntr [11]),
    .e(\PWMB/FreCntr [4]),
    .o(_al_u2639_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u264 (
    .a(\PWM2/pnumr [27]),
    .b(pnum2[27]),
    .c(pnum2[32]),
    .d(pwm_start_stop[18]),
    .o(\PWM2/n23 [27]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u2640 (
    .a(\PWMB/FreCnt [1]),
    .b(\PWMB/FreCnt [23]),
    .c(\PWMB/FreCntr [2]),
    .d(\PWMB/FreCntr [24]),
    .o(_al_u2640_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u2641 (
    .a(_al_u2637_o),
    .b(_al_u2639_o),
    .c(_al_u2640_o),
    .d(\PWMB/FreCnt [12]),
    .e(\PWMB/FreCntr [13]),
    .o(_al_u2641_o));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(E@B)*~(~D*A))"),
    .INIT(32'h0c040301))
    _al_u2642 (
    .a(\PWMB/FreCnt [11]),
    .b(\PWMB/FreCnt [2]),
    .c(\PWMB/FreCnt [26]),
    .d(\PWMB/FreCntr [12]),
    .e(\PWMB/FreCntr [3]),
    .o(_al_u2642_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u2643 (
    .a(_al_u2642_o),
    .b(\PWMB/FreCnt [24]),
    .c(\PWMB/FreCnt [4]),
    .d(\PWMB/FreCntr [25]),
    .e(\PWMB/FreCntr [5]),
    .o(_al_u2643_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u2644 (
    .a(\PWMB/FreCnt [20]),
    .b(\PWMB/FreCnt [6]),
    .c(\PWMB/FreCntr [21]),
    .d(\PWMB/FreCntr [7]),
    .o(_al_u2644_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u2645 (
    .a(_al_u2644_o),
    .b(\PWMB/FreCnt [0]),
    .c(\PWMB/FreCntr [1]),
    .o(_al_u2645_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u2646 (
    .a(\PWMB/FreCnt [7]),
    .b(\PWMB/FreCnt [8]),
    .c(\PWMB/FreCntr [8]),
    .d(\PWMB/FreCntr [9]),
    .o(_al_u2646_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*C)*~(~D*B))"),
    .INIT(32'haa220a02))
    _al_u2647 (
    .a(_al_u2646_o),
    .b(\PWMB/FreCnt [17]),
    .c(\PWMB/FreCnt [25]),
    .d(\PWMB/FreCntr [18]),
    .e(\PWMB/FreCntr [26]),
    .o(_al_u2647_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2648 (
    .a(\PWMB/FreCnt [19]),
    .b(\PWMB/FreCntr [20]),
    .o(_al_u2648_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(E@C)*~(D*~B))"),
    .INIT(32'h40500405))
    _al_u2649 (
    .a(_al_u2648_o),
    .b(\PWMB/FreCnt [11]),
    .c(\PWMB/FreCnt [18]),
    .d(\PWMB/FreCntr [12]),
    .e(\PWMB/FreCntr [19]),
    .o(_al_u2649_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u265 (
    .a(\PWM2/pnumr [26]),
    .b(pnum2[26]),
    .c(pnum2[32]),
    .d(pwm_start_stop[18]),
    .o(\PWM2/n23 [26]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u2650 (
    .a(_al_u2643_o),
    .b(_al_u2645_o),
    .c(_al_u2647_o),
    .d(_al_u2649_o),
    .o(_al_u2650_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2651 (
    .a(\PWMB/FreCnt [21]),
    .b(\PWMB/FreCntr [22]),
    .o(_al_u2651_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(~E*C)*~(D@B))"),
    .INIT(32'h44110401))
    _al_u2652 (
    .a(_al_u2651_o),
    .b(\PWMB/FreCnt [13]),
    .c(\PWMB/FreCnt [15]),
    .d(\PWMB/FreCntr [14]),
    .e(\PWMB/FreCntr [16]),
    .o(_al_u2652_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u2653 (
    .a(_al_u2652_o),
    .b(\PWMB/FreCnt [14]),
    .c(\PWMB/FreCnt [22]),
    .d(\PWMB/FreCntr [15]),
    .e(\PWMB/FreCntr [23]),
    .o(_al_u2653_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(~D*A))"),
    .INIT(16'hcf45))
    _al_u2654 (
    .a(\PWMB/FreCnt [23]),
    .b(\PWMB/FreCnt [9]),
    .c(\PWMB/FreCntr [10]),
    .d(\PWMB/FreCntr [24]),
    .o(_al_u2654_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*C)*~(D*~B))"),
    .INIT(32'h88aa080a))
    _al_u2655 (
    .a(_al_u2654_o),
    .b(\PWMB/FreCnt [1]),
    .c(\PWMB/FreCnt [5]),
    .d(\PWMB/FreCntr [2]),
    .e(\PWMB/FreCntr [6]),
    .o(_al_u2655_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2656 (
    .a(\PWMB/FreCnt [15]),
    .b(\PWMB/FreCntr [16]),
    .o(_al_u2656_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(~D*C)*~(E@B))"),
    .INIT(32'h44041101))
    _al_u2657 (
    .a(_al_u2656_o),
    .b(\PWMB/FreCnt [16]),
    .c(\PWMB/FreCnt [9]),
    .d(\PWMB/FreCntr [10]),
    .e(\PWMB/FreCntr [17]),
    .o(_al_u2657_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    _al_u2658 (
    .a(_al_u2641_o),
    .b(_al_u2650_o),
    .c(_al_u2653_o),
    .d(_al_u2655_o),
    .e(_al_u2657_o),
    .o(_al_u2658_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2659 (
    .a(_al_u2658_o),
    .b(pwm_state_read[11]),
    .o(\PWMB/u14_sel_is_1_o ));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u266 (
    .a(\PWM2/pnumr [25]),
    .b(pnum2[25]),
    .c(pnum2[32]),
    .d(pwm_start_stop[18]),
    .o(\PWM2/n23 [25]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2660 (
    .a(\PWMC/n0_lutinv ),
    .b(pwm_state_read[12]),
    .o(\PWMC/n24 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u2661 (
    .a(pnumcntC[18]),
    .b(pnumcntC[19]),
    .c(pnumcntC[1]),
    .d(pnumcntC[20]),
    .o(_al_u2661_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u2662 (
    .a(_al_u2661_o),
    .b(pnumcntC[21]),
    .c(pnumcntC[22]),
    .d(pnumcntC[23]),
    .e(pnumcntC[2]),
    .o(_al_u2662_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u2663 (
    .a(_al_u2662_o),
    .b(pnumcntC[6]),
    .c(pnumcntC[7]),
    .d(pnumcntC[8]),
    .e(pnumcntC[9]),
    .o(_al_u2663_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u2664 (
    .a(pnumcntC[10]),
    .b(pnumcntC[11]),
    .c(pnumcntC[12]),
    .d(pnumcntC[13]),
    .o(_al_u2664_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u2665 (
    .a(_al_u2664_o),
    .b(pnumcntC[14]),
    .c(pnumcntC[15]),
    .d(pnumcntC[16]),
    .e(pnumcntC[17]),
    .o(_al_u2665_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u2666 (
    .a(pnumcntC[3]),
    .b(pnumcntC[4]),
    .c(pnumcntC[5]),
    .o(_al_u2666_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u2667 (
    .a(_al_u2663_o),
    .b(_al_u2665_o),
    .c(_al_u2666_o),
    .d(pnumcntC[0]),
    .o(\PWMC/n25_neg_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2668 (
    .a(\PWMC/n24 ),
    .b(\PWMC/n25_neg_lutinv ),
    .c(\PWMC/n26 [9]),
    .d(\PWMC/pnumr [9]),
    .o(_al_u2668_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2669 (
    .a(_al_u2668_o),
    .b(\PWMC/n24 ),
    .c(pnumcntC[9]),
    .d(\PWMC/pnumr [9]),
    .e(pwm_start_stop[28]),
    .o(\PWMC/n31 [9]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u267 (
    .a(\PWM2/pnumr [24]),
    .b(pnum2[24]),
    .c(pnum2[32]),
    .d(pwm_start_stop[18]),
    .o(\PWM2/n23 [24]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2670 (
    .a(\PWMC/n24 ),
    .b(\PWMC/n25_neg_lutinv ),
    .c(\PWMC/n26 [8]),
    .d(\PWMC/pnumr [8]),
    .o(_al_u2670_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2671 (
    .a(_al_u2670_o),
    .b(\PWMC/n24 ),
    .c(pnumcntC[8]),
    .d(\PWMC/pnumr [8]),
    .e(pwm_start_stop[28]),
    .o(\PWMC/n31 [8]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2672 (
    .a(\PWMC/n24 ),
    .b(\PWMC/n25_neg_lutinv ),
    .c(\PWMC/n26 [7]),
    .d(\PWMC/pnumr [7]),
    .o(_al_u2672_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2673 (
    .a(_al_u2672_o),
    .b(\PWMC/n24 ),
    .c(pnumcntC[7]),
    .d(\PWMC/pnumr [7]),
    .e(pwm_start_stop[28]),
    .o(\PWMC/n31 [7]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2674 (
    .a(\PWMC/n24 ),
    .b(\PWMC/n25_neg_lutinv ),
    .c(\PWMC/n26 [6]),
    .d(\PWMC/pnumr [6]),
    .o(_al_u2674_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2675 (
    .a(_al_u2674_o),
    .b(\PWMC/n24 ),
    .c(pnumcntC[6]),
    .d(\PWMC/pnumr [6]),
    .e(pwm_start_stop[28]),
    .o(\PWMC/n31 [6]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2676 (
    .a(\PWMC/n24 ),
    .b(\PWMC/n25_neg_lutinv ),
    .c(\PWMC/n26 [5]),
    .d(\PWMC/pnumr [5]),
    .o(_al_u2676_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2677 (
    .a(_al_u2676_o),
    .b(\PWMC/n24 ),
    .c(pnumcntC[5]),
    .d(\PWMC/pnumr [5]),
    .e(pwm_start_stop[28]),
    .o(\PWMC/n31 [5]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2678 (
    .a(\PWMC/n24 ),
    .b(\PWMC/n25_neg_lutinv ),
    .c(\PWMC/n26 [4]),
    .d(\PWMC/pnumr [4]),
    .o(_al_u2678_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2679 (
    .a(_al_u2678_o),
    .b(\PWMC/n24 ),
    .c(pnumcntC[4]),
    .d(\PWMC/pnumr [4]),
    .e(pwm_start_stop[28]),
    .o(\PWMC/n31 [4]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u268 (
    .a(\PWM2/pnumr [23]),
    .b(pnum2[23]),
    .c(pnum2[32]),
    .d(pwm_start_stop[18]),
    .o(\PWM2/n23 [23]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2680 (
    .a(\PWMC/n24 ),
    .b(\PWMC/n25_neg_lutinv ),
    .c(\PWMC/n26 [3]),
    .d(\PWMC/pnumr [3]),
    .o(_al_u2680_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2681 (
    .a(_al_u2680_o),
    .b(\PWMC/n24 ),
    .c(pnumcntC[3]),
    .d(\PWMC/pnumr [3]),
    .e(pwm_start_stop[28]),
    .o(\PWMC/n31 [3]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2682 (
    .a(\PWMC/n24 ),
    .b(\PWMC/n25_neg_lutinv ),
    .c(\PWMC/n26 [23]),
    .d(\PWMC/pnumr [23]),
    .o(_al_u2682_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2683 (
    .a(_al_u2682_o),
    .b(\PWMC/n24 ),
    .c(pnumcntC[23]),
    .d(\PWMC/pnumr [23]),
    .e(pwm_start_stop[28]),
    .o(\PWMC/n31 [23]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2684 (
    .a(\PWMC/n24 ),
    .b(\PWMC/n25_neg_lutinv ),
    .c(\PWMC/n26 [22]),
    .d(\PWMC/pnumr [22]),
    .o(_al_u2684_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2685 (
    .a(_al_u2684_o),
    .b(\PWMC/n24 ),
    .c(pnumcntC[22]),
    .d(\PWMC/pnumr [22]),
    .e(pwm_start_stop[28]),
    .o(\PWMC/n31 [22]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2686 (
    .a(\PWMC/n24 ),
    .b(\PWMC/n25_neg_lutinv ),
    .c(\PWMC/n26 [21]),
    .d(\PWMC/pnumr [21]),
    .o(_al_u2686_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2687 (
    .a(_al_u2686_o),
    .b(\PWMC/n24 ),
    .c(pnumcntC[21]),
    .d(\PWMC/pnumr [21]),
    .e(pwm_start_stop[28]),
    .o(\PWMC/n31 [21]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2688 (
    .a(\PWMC/n24 ),
    .b(\PWMC/n25_neg_lutinv ),
    .c(\PWMC/n26 [20]),
    .d(\PWMC/pnumr [20]),
    .o(_al_u2688_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2689 (
    .a(_al_u2688_o),
    .b(\PWMC/n24 ),
    .c(pnumcntC[20]),
    .d(\PWMC/pnumr [20]),
    .e(pwm_start_stop[28]),
    .o(\PWMC/n31 [20]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u269 (
    .a(\PWM2/pnumr [22]),
    .b(pnum2[22]),
    .c(pnum2[32]),
    .d(pwm_start_stop[18]),
    .o(\PWM2/n23 [22]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2690 (
    .a(\PWMC/n24 ),
    .b(\PWMC/n25_neg_lutinv ),
    .c(\PWMC/n26 [2]),
    .d(\PWMC/pnumr [2]),
    .o(_al_u2690_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2691 (
    .a(_al_u2690_o),
    .b(\PWMC/n24 ),
    .c(pnumcntC[2]),
    .d(\PWMC/pnumr [2]),
    .e(pwm_start_stop[28]),
    .o(\PWMC/n31 [2]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2692 (
    .a(\PWMC/n24 ),
    .b(\PWMC/n25_neg_lutinv ),
    .c(\PWMC/n26 [19]),
    .d(\PWMC/pnumr [19]),
    .o(_al_u2692_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2693 (
    .a(_al_u2692_o),
    .b(\PWMC/n24 ),
    .c(pnumcntC[19]),
    .d(\PWMC/pnumr [19]),
    .e(pwm_start_stop[28]),
    .o(\PWMC/n31 [19]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2694 (
    .a(\PWMC/n24 ),
    .b(\PWMC/n25_neg_lutinv ),
    .c(\PWMC/n26 [18]),
    .d(\PWMC/pnumr [18]),
    .o(_al_u2694_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2695 (
    .a(_al_u2694_o),
    .b(\PWMC/n24 ),
    .c(pnumcntC[18]),
    .d(\PWMC/pnumr [18]),
    .e(pwm_start_stop[28]),
    .o(\PWMC/n31 [18]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2696 (
    .a(\PWMC/n24 ),
    .b(\PWMC/n25_neg_lutinv ),
    .c(\PWMC/n26 [17]),
    .d(\PWMC/pnumr [17]),
    .o(_al_u2696_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2697 (
    .a(_al_u2696_o),
    .b(\PWMC/n24 ),
    .c(pnumcntC[17]),
    .d(\PWMC/pnumr [17]),
    .e(pwm_start_stop[28]),
    .o(\PWMC/n31 [17]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2698 (
    .a(\PWMC/n24 ),
    .b(\PWMC/n25_neg_lutinv ),
    .c(\PWMC/n26 [16]),
    .d(\PWMC/pnumr [16]),
    .o(_al_u2698_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2699 (
    .a(_al_u2698_o),
    .b(\PWMC/n24 ),
    .c(pnumcntC[16]),
    .d(\PWMC/pnumr [16]),
    .e(pwm_start_stop[28]),
    .o(\PWMC/n31 [16]));
  EF2_PHY_PAD #(
    //.LOCATION("P43"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u27 (
    .do({open_n846,open_n847,open_n848,dir_pad[11]}),
    .opad(dir[11]));  // CPLD_SOC_AHB_TOP.v(7)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u270 (
    .a(\PWM2/pnumr [21]),
    .b(pnum2[21]),
    .c(pnum2[32]),
    .d(pwm_start_stop[18]),
    .o(\PWM2/n23 [21]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2700 (
    .a(\PWMC/n24 ),
    .b(\PWMC/n25_neg_lutinv ),
    .c(\PWMC/n26 [15]),
    .d(\PWMC/pnumr [15]),
    .o(_al_u2700_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2701 (
    .a(_al_u2700_o),
    .b(\PWMC/n24 ),
    .c(pnumcntC[15]),
    .d(\PWMC/pnumr [15]),
    .e(pwm_start_stop[28]),
    .o(\PWMC/n31 [15]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2702 (
    .a(\PWMC/n24 ),
    .b(\PWMC/n25_neg_lutinv ),
    .c(\PWMC/n26 [14]),
    .d(\PWMC/pnumr [14]),
    .o(_al_u2702_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2703 (
    .a(_al_u2702_o),
    .b(\PWMC/n24 ),
    .c(pnumcntC[14]),
    .d(\PWMC/pnumr [14]),
    .e(pwm_start_stop[28]),
    .o(\PWMC/n31 [14]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2704 (
    .a(\PWMC/n24 ),
    .b(\PWMC/n25_neg_lutinv ),
    .c(\PWMC/n26 [13]),
    .d(\PWMC/pnumr [13]),
    .o(_al_u2704_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2705 (
    .a(_al_u2704_o),
    .b(\PWMC/n24 ),
    .c(pnumcntC[13]),
    .d(\PWMC/pnumr [13]),
    .e(pwm_start_stop[28]),
    .o(\PWMC/n31 [13]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2706 (
    .a(\PWMC/n24 ),
    .b(\PWMC/n25_neg_lutinv ),
    .c(\PWMC/n26 [12]),
    .d(\PWMC/pnumr [12]),
    .o(_al_u2706_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2707 (
    .a(_al_u2706_o),
    .b(\PWMC/n24 ),
    .c(pnumcntC[12]),
    .d(\PWMC/pnumr [12]),
    .e(pwm_start_stop[28]),
    .o(\PWMC/n31 [12]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2708 (
    .a(\PWMC/n24 ),
    .b(\PWMC/n25_neg_lutinv ),
    .c(\PWMC/n26 [11]),
    .d(\PWMC/pnumr [11]),
    .o(_al_u2708_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2709 (
    .a(_al_u2708_o),
    .b(\PWMC/n24 ),
    .c(pnumcntC[11]),
    .d(\PWMC/pnumr [11]),
    .e(pwm_start_stop[28]),
    .o(\PWMC/n31 [11]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u271 (
    .a(\PWM2/pnumr [20]),
    .b(pnum2[20]),
    .c(pnum2[32]),
    .d(pwm_start_stop[18]),
    .o(\PWM2/n23 [20]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2710 (
    .a(\PWMC/n24 ),
    .b(\PWMC/n25_neg_lutinv ),
    .c(\PWMC/n26 [10]),
    .d(\PWMC/pnumr [10]),
    .o(_al_u2710_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2711 (
    .a(_al_u2710_o),
    .b(\PWMC/n24 ),
    .c(pnumcntC[10]),
    .d(\PWMC/pnumr [10]),
    .e(pwm_start_stop[28]),
    .o(\PWMC/n31 [10]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2712 (
    .a(\PWMC/n24 ),
    .b(\PWMC/n25_neg_lutinv ),
    .c(\PWMC/n26 [1]),
    .d(\PWMC/pnumr [1]),
    .o(_al_u2712_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2713 (
    .a(_al_u2712_o),
    .b(\PWMC/n24 ),
    .c(pnumcntC[1]),
    .d(\PWMC/pnumr [1]),
    .e(pwm_start_stop[28]),
    .o(\PWMC/n31 [1]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2714 (
    .a(\PWMC/n24 ),
    .b(\PWMC/n25_neg_lutinv ),
    .c(\PWMC/n26 [0]),
    .d(\PWMC/pnumr [0]),
    .o(_al_u2714_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2715 (
    .a(_al_u2714_o),
    .b(\PWMC/n24 ),
    .c(pnumcntC[0]),
    .d(\PWMC/pnumr [0]),
    .e(pwm_start_stop[28]),
    .o(\PWMC/n31 [0]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2716 (
    .a(\PWMC/FreCnt [25]),
    .b(\PWMC/FreCntr [26]),
    .o(_al_u2716_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(~E*C)*~(D@B))"),
    .INIT(32'h44110401))
    _al_u2717 (
    .a(_al_u2716_o),
    .b(\PWMC/FreCnt [1]),
    .c(\PWMC/FreCnt [21]),
    .d(\PWMC/FreCntr [2]),
    .e(\PWMC/FreCntr [22]),
    .o(_al_u2717_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u2718 (
    .a(\PWMC/FreCnt [10]),
    .b(\PWMC/FreCnt [5]),
    .c(\PWMC/FreCntr [11]),
    .d(\PWMC/FreCntr [6]),
    .o(_al_u2718_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*~C))"),
    .INIT(16'h8088))
    _al_u2719 (
    .a(_al_u2717_o),
    .b(_al_u2718_o),
    .c(\PWMC/FreCnt [23]),
    .d(\PWMC/FreCntr [24]),
    .o(_al_u2719_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u272 (
    .a(\PWM2/pnumr [2]),
    .b(pnum2[2]),
    .c(pnum2[32]),
    .d(pwm_start_stop[18]),
    .o(\PWM2/n23 [2]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u2720 (
    .a(\PWMC/FreCnt [17]),
    .b(\PWMC/FreCnt [21]),
    .c(\PWMC/FreCntr [18]),
    .d(\PWMC/FreCntr [22]),
    .o(_al_u2720_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*C)*~(D*~B))"),
    .INIT(32'h88aa080a))
    _al_u2721 (
    .a(_al_u2720_o),
    .b(\PWMC/FreCnt [15]),
    .c(\PWMC/FreCnt [19]),
    .d(\PWMC/FreCntr [16]),
    .e(\PWMC/FreCntr [20]),
    .o(_al_u2721_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u2722 (
    .a(\PWMC/FreCnt [15]),
    .b(\PWMC/FreCnt [17]),
    .c(\PWMC/FreCntr [16]),
    .d(\PWMC/FreCntr [18]),
    .o(_al_u2722_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u2723 (
    .a(_al_u2719_o),
    .b(_al_u2721_o),
    .c(_al_u2722_o),
    .d(\PWMC/FreCnt [24]),
    .e(\PWMC/FreCntr [25]),
    .o(_al_u2723_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u2724 (
    .a(\PWMC/FreCnt [14]),
    .b(\PWMC/FreCnt [4]),
    .c(\PWMC/FreCntr [15]),
    .d(\PWMC/FreCntr [5]),
    .o(_al_u2724_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u2725 (
    .a(_al_u2724_o),
    .b(\PWMC/FreCnt [13]),
    .c(\PWMC/FreCntr [14]),
    .o(_al_u2725_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u2726 (
    .a(\PWMC/FreCnt [18]),
    .b(\PWMC/FreCnt [2]),
    .c(\PWMC/FreCntr [19]),
    .d(\PWMC/FreCntr [3]),
    .o(_al_u2726_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u2727 (
    .a(_al_u2726_o),
    .b(\PWMC/FreCnt [20]),
    .c(\PWMC/FreCnt [22]),
    .d(\PWMC/FreCntr [21]),
    .e(\PWMC/FreCntr [23]),
    .o(_al_u2727_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u2728 (
    .a(\PWMC/FreCnt [10]),
    .b(\PWMC/FreCnt [3]),
    .c(\PWMC/FreCntr [11]),
    .d(\PWMC/FreCntr [4]),
    .o(_al_u2728_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*C)*~(D*~B))"),
    .INIT(32'h88aa080a))
    _al_u2729 (
    .a(_al_u2728_o),
    .b(\PWMC/FreCnt [16]),
    .c(\PWMC/FreCnt [7]),
    .d(\PWMC/FreCntr [17]),
    .e(\PWMC/FreCntr [8]),
    .o(_al_u2729_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u273 (
    .a(\PWM2/pnumr [19]),
    .b(pnum2[19]),
    .c(pnum2[32]),
    .d(pwm_start_stop[18]),
    .o(\PWM2/n23 [19]));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(~E*B)*~(D@A))"),
    .INIT(32'h0a050201))
    _al_u2730 (
    .a(\PWMC/FreCnt [11]),
    .b(\PWMC/FreCnt [16]),
    .c(\PWMC/FreCnt [26]),
    .d(\PWMC/FreCntr [12]),
    .e(\PWMC/FreCntr [17]),
    .o(_al_u2730_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u2731 (
    .a(_al_u2725_o),
    .b(_al_u2727_o),
    .c(_al_u2729_o),
    .d(_al_u2730_o),
    .o(_al_u2731_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u2732 (
    .a(\PWMC/FreCnt [19]),
    .b(\PWMC/FreCnt [7]),
    .c(\PWMC/FreCntr [20]),
    .d(\PWMC/FreCntr [8]),
    .o(_al_u2732_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*~C)*~(~D*B))"),
    .INIT(32'ha020aa22))
    _al_u2733 (
    .a(_al_u2732_o),
    .b(\PWMC/FreCnt [23]),
    .c(\PWMC/FreCnt [5]),
    .d(\PWMC/FreCntr [24]),
    .e(\PWMC/FreCntr [6]),
    .o(_al_u2733_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u2734 (
    .a(\PWMC/FreCnt [0]),
    .b(\PWMC/FreCnt [8]),
    .c(\PWMC/FreCntr [1]),
    .d(\PWMC/FreCntr [9]),
    .o(_al_u2734_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D@C)*~(E@B))"),
    .INIT(32'h80082002))
    _al_u2735 (
    .a(_al_u2734_o),
    .b(\PWMC/FreCnt [6]),
    .c(\PWMC/FreCnt [9]),
    .d(\PWMC/FreCntr [10]),
    .e(\PWMC/FreCntr [7]),
    .o(_al_u2735_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u2736 (
    .a(\PWMC/FreCnt [25]),
    .b(\PWMC/FreCnt [3]),
    .c(\PWMC/FreCntr [26]),
    .d(\PWMC/FreCntr [4]),
    .o(_al_u2736_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u2737 (
    .a(_al_u2733_o),
    .b(_al_u2735_o),
    .c(_al_u2736_o),
    .d(\PWMC/FreCnt [12]),
    .e(\PWMC/FreCntr [13]),
    .o(_al_u2737_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*A))"),
    .INIT(16'h7f00))
    _al_u2738 (
    .a(_al_u2723_o),
    .b(_al_u2731_o),
    .c(_al_u2737_o),
    .d(pwm_state_read[12]),
    .o(\PWMC/u14_sel_is_1_o ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2739 (
    .a(\PWMD/n0_lutinv ),
    .b(pwm_state_read[13]),
    .o(\PWMD/n24 ));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u274 (
    .a(\PWM2/pnumr [18]),
    .b(pnum2[18]),
    .c(pnum2[32]),
    .d(pwm_start_stop[18]),
    .o(\PWM2/n23 [18]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u2740 (
    .a(pnumcntD[18]),
    .b(pnumcntD[19]),
    .c(pnumcntD[1]),
    .d(pnumcntD[20]),
    .o(_al_u2740_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u2741 (
    .a(_al_u2740_o),
    .b(pnumcntD[21]),
    .c(pnumcntD[22]),
    .d(pnumcntD[23]),
    .e(pnumcntD[2]),
    .o(_al_u2741_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u2742 (
    .a(_al_u2741_o),
    .b(pnumcntD[6]),
    .c(pnumcntD[7]),
    .d(pnumcntD[8]),
    .e(pnumcntD[9]),
    .o(_al_u2742_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u2743 (
    .a(pnumcntD[10]),
    .b(pnumcntD[11]),
    .c(pnumcntD[12]),
    .d(pnumcntD[13]),
    .o(_al_u2743_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u2744 (
    .a(_al_u2743_o),
    .b(pnumcntD[14]),
    .c(pnumcntD[15]),
    .d(pnumcntD[16]),
    .e(pnumcntD[17]),
    .o(_al_u2744_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u2745 (
    .a(pnumcntD[3]),
    .b(pnumcntD[4]),
    .c(pnumcntD[5]),
    .o(_al_u2745_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u2746 (
    .a(_al_u2742_o),
    .b(_al_u2744_o),
    .c(_al_u2745_o),
    .d(pnumcntD[0]),
    .o(\PWMD/n25_neg_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2747 (
    .a(\PWMD/n24 ),
    .b(\PWMD/n25_neg_lutinv ),
    .c(\PWMD/n26 [9]),
    .d(\PWMD/pnumr [9]),
    .o(_al_u2747_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2748 (
    .a(_al_u2747_o),
    .b(\PWMD/n24 ),
    .c(pnumcntD[9]),
    .d(\PWMD/pnumr [9]),
    .e(pwm_start_stop[29]),
    .o(\PWMD/n31 [9]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2749 (
    .a(\PWMD/n24 ),
    .b(\PWMD/n25_neg_lutinv ),
    .c(\PWMD/n26 [8]),
    .d(\PWMD/pnumr [8]),
    .o(_al_u2749_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u275 (
    .a(\PWM2/pnumr [17]),
    .b(pnum2[17]),
    .c(pnum2[32]),
    .d(pwm_start_stop[18]),
    .o(\PWM2/n23 [17]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2750 (
    .a(_al_u2749_o),
    .b(\PWMD/n24 ),
    .c(pnumcntD[8]),
    .d(\PWMD/pnumr [8]),
    .e(pwm_start_stop[29]),
    .o(\PWMD/n31 [8]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2751 (
    .a(\PWMD/n24 ),
    .b(\PWMD/n25_neg_lutinv ),
    .c(\PWMD/n26 [7]),
    .d(\PWMD/pnumr [7]),
    .o(_al_u2751_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2752 (
    .a(_al_u2751_o),
    .b(\PWMD/n24 ),
    .c(pnumcntD[7]),
    .d(\PWMD/pnumr [7]),
    .e(pwm_start_stop[29]),
    .o(\PWMD/n31 [7]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2753 (
    .a(\PWMD/n24 ),
    .b(\PWMD/n25_neg_lutinv ),
    .c(\PWMD/n26 [6]),
    .d(\PWMD/pnumr [6]),
    .o(_al_u2753_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2754 (
    .a(_al_u2753_o),
    .b(\PWMD/n24 ),
    .c(pnumcntD[6]),
    .d(\PWMD/pnumr [6]),
    .e(pwm_start_stop[29]),
    .o(\PWMD/n31 [6]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2755 (
    .a(\PWMD/n24 ),
    .b(\PWMD/n25_neg_lutinv ),
    .c(\PWMD/n26 [5]),
    .d(\PWMD/pnumr [5]),
    .o(_al_u2755_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2756 (
    .a(_al_u2755_o),
    .b(\PWMD/n24 ),
    .c(pnumcntD[5]),
    .d(\PWMD/pnumr [5]),
    .e(pwm_start_stop[29]),
    .o(\PWMD/n31 [5]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2757 (
    .a(\PWMD/n24 ),
    .b(\PWMD/n25_neg_lutinv ),
    .c(\PWMD/n26 [4]),
    .d(\PWMD/pnumr [4]),
    .o(_al_u2757_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2758 (
    .a(_al_u2757_o),
    .b(\PWMD/n24 ),
    .c(pnumcntD[4]),
    .d(\PWMD/pnumr [4]),
    .e(pwm_start_stop[29]),
    .o(\PWMD/n31 [4]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2759 (
    .a(\PWMD/n24 ),
    .b(\PWMD/n25_neg_lutinv ),
    .c(\PWMD/n26 [3]),
    .d(\PWMD/pnumr [3]),
    .o(_al_u2759_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u276 (
    .a(\PWM2/pnumr [16]),
    .b(pnum2[16]),
    .c(pnum2[32]),
    .d(pwm_start_stop[18]),
    .o(\PWM2/n23 [16]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2760 (
    .a(_al_u2759_o),
    .b(\PWMD/n24 ),
    .c(pnumcntD[3]),
    .d(\PWMD/pnumr [3]),
    .e(pwm_start_stop[29]),
    .o(\PWMD/n31 [3]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2761 (
    .a(\PWMD/n24 ),
    .b(\PWMD/n25_neg_lutinv ),
    .c(\PWMD/n26 [23]),
    .d(\PWMD/pnumr [23]),
    .o(_al_u2761_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2762 (
    .a(_al_u2761_o),
    .b(\PWMD/n24 ),
    .c(pnumcntD[23]),
    .d(\PWMD/pnumr [23]),
    .e(pwm_start_stop[29]),
    .o(\PWMD/n31 [23]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2763 (
    .a(\PWMD/n24 ),
    .b(\PWMD/n25_neg_lutinv ),
    .c(\PWMD/n26 [22]),
    .d(\PWMD/pnumr [22]),
    .o(_al_u2763_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2764 (
    .a(_al_u2763_o),
    .b(\PWMD/n24 ),
    .c(pnumcntD[22]),
    .d(\PWMD/pnumr [22]),
    .e(pwm_start_stop[29]),
    .o(\PWMD/n31 [22]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2765 (
    .a(\PWMD/n24 ),
    .b(\PWMD/n25_neg_lutinv ),
    .c(\PWMD/n26 [21]),
    .d(\PWMD/pnumr [21]),
    .o(_al_u2765_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2766 (
    .a(_al_u2765_o),
    .b(\PWMD/n24 ),
    .c(pnumcntD[21]),
    .d(\PWMD/pnumr [21]),
    .e(pwm_start_stop[29]),
    .o(\PWMD/n31 [21]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2767 (
    .a(\PWMD/n24 ),
    .b(\PWMD/n25_neg_lutinv ),
    .c(\PWMD/n26 [20]),
    .d(\PWMD/pnumr [20]),
    .o(_al_u2767_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2768 (
    .a(_al_u2767_o),
    .b(\PWMD/n24 ),
    .c(pnumcntD[20]),
    .d(\PWMD/pnumr [20]),
    .e(pwm_start_stop[29]),
    .o(\PWMD/n31 [20]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2769 (
    .a(\PWMD/n24 ),
    .b(\PWMD/n25_neg_lutinv ),
    .c(\PWMD/n26 [2]),
    .d(\PWMD/pnumr [2]),
    .o(_al_u2769_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u277 (
    .a(\PWM2/pnumr [15]),
    .b(pnum2[15]),
    .c(pnum2[32]),
    .d(pwm_start_stop[18]),
    .o(\PWM2/n23 [15]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2770 (
    .a(_al_u2769_o),
    .b(\PWMD/n24 ),
    .c(pnumcntD[2]),
    .d(\PWMD/pnumr [2]),
    .e(pwm_start_stop[29]),
    .o(\PWMD/n31 [2]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2771 (
    .a(\PWMD/n24 ),
    .b(\PWMD/n25_neg_lutinv ),
    .c(\PWMD/n26 [19]),
    .d(\PWMD/pnumr [19]),
    .o(_al_u2771_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2772 (
    .a(_al_u2771_o),
    .b(\PWMD/n24 ),
    .c(pnumcntD[19]),
    .d(\PWMD/pnumr [19]),
    .e(pwm_start_stop[29]),
    .o(\PWMD/n31 [19]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2773 (
    .a(\PWMD/n24 ),
    .b(\PWMD/n25_neg_lutinv ),
    .c(\PWMD/n26 [18]),
    .d(\PWMD/pnumr [18]),
    .o(_al_u2773_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2774 (
    .a(_al_u2773_o),
    .b(\PWMD/n24 ),
    .c(pnumcntD[18]),
    .d(\PWMD/pnumr [18]),
    .e(pwm_start_stop[29]),
    .o(\PWMD/n31 [18]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2775 (
    .a(\PWMD/n24 ),
    .b(\PWMD/n25_neg_lutinv ),
    .c(\PWMD/n26 [17]),
    .d(\PWMD/pnumr [17]),
    .o(_al_u2775_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2776 (
    .a(_al_u2775_o),
    .b(\PWMD/n24 ),
    .c(pnumcntD[17]),
    .d(\PWMD/pnumr [17]),
    .e(pwm_start_stop[29]),
    .o(\PWMD/n31 [17]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2777 (
    .a(\PWMD/n24 ),
    .b(\PWMD/n25_neg_lutinv ),
    .c(\PWMD/n26 [16]),
    .d(\PWMD/pnumr [16]),
    .o(_al_u2777_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2778 (
    .a(_al_u2777_o),
    .b(\PWMD/n24 ),
    .c(pnumcntD[16]),
    .d(\PWMD/pnumr [16]),
    .e(pwm_start_stop[29]),
    .o(\PWMD/n31 [16]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2779 (
    .a(\PWMD/n24 ),
    .b(\PWMD/n25_neg_lutinv ),
    .c(\PWMD/n26 [15]),
    .d(\PWMD/pnumr [15]),
    .o(_al_u2779_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u278 (
    .a(\PWM2/pnumr [14]),
    .b(pnum2[14]),
    .c(pnum2[32]),
    .d(pwm_start_stop[18]),
    .o(\PWM2/n23 [14]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2780 (
    .a(_al_u2779_o),
    .b(\PWMD/n24 ),
    .c(pnumcntD[15]),
    .d(\PWMD/pnumr [15]),
    .e(pwm_start_stop[29]),
    .o(\PWMD/n31 [15]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2781 (
    .a(\PWMD/n24 ),
    .b(\PWMD/n25_neg_lutinv ),
    .c(\PWMD/n26 [14]),
    .d(\PWMD/pnumr [14]),
    .o(_al_u2781_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2782 (
    .a(_al_u2781_o),
    .b(\PWMD/n24 ),
    .c(pnumcntD[14]),
    .d(\PWMD/pnumr [14]),
    .e(pwm_start_stop[29]),
    .o(\PWMD/n31 [14]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2783 (
    .a(\PWMD/n24 ),
    .b(\PWMD/n25_neg_lutinv ),
    .c(\PWMD/n26 [13]),
    .d(\PWMD/pnumr [13]),
    .o(_al_u2783_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2784 (
    .a(_al_u2783_o),
    .b(\PWMD/n24 ),
    .c(pnumcntD[13]),
    .d(\PWMD/pnumr [13]),
    .e(pwm_start_stop[29]),
    .o(\PWMD/n31 [13]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2785 (
    .a(\PWMD/n24 ),
    .b(\PWMD/n25_neg_lutinv ),
    .c(\PWMD/n26 [12]),
    .d(\PWMD/pnumr [12]),
    .o(_al_u2785_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2786 (
    .a(_al_u2785_o),
    .b(\PWMD/n24 ),
    .c(pnumcntD[12]),
    .d(\PWMD/pnumr [12]),
    .e(pwm_start_stop[29]),
    .o(\PWMD/n31 [12]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2787 (
    .a(\PWMD/n24 ),
    .b(\PWMD/n25_neg_lutinv ),
    .c(\PWMD/n26 [11]),
    .d(\PWMD/pnumr [11]),
    .o(_al_u2787_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2788 (
    .a(_al_u2787_o),
    .b(\PWMD/n24 ),
    .c(pnumcntD[11]),
    .d(\PWMD/pnumr [11]),
    .e(pwm_start_stop[29]),
    .o(\PWMD/n31 [11]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2789 (
    .a(\PWMD/n24 ),
    .b(\PWMD/n25_neg_lutinv ),
    .c(\PWMD/n26 [10]),
    .d(\PWMD/pnumr [10]),
    .o(_al_u2789_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u279 (
    .a(\PWM2/pnumr [13]),
    .b(pnum2[13]),
    .c(pnum2[32]),
    .d(pwm_start_stop[18]),
    .o(\PWM2/n23 [13]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2790 (
    .a(_al_u2789_o),
    .b(\PWMD/n24 ),
    .c(pnumcntD[10]),
    .d(\PWMD/pnumr [10]),
    .e(pwm_start_stop[29]),
    .o(\PWMD/n31 [10]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2791 (
    .a(\PWMD/n24 ),
    .b(\PWMD/n25_neg_lutinv ),
    .c(\PWMD/n26 [1]),
    .d(\PWMD/pnumr [1]),
    .o(_al_u2791_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2792 (
    .a(_al_u2791_o),
    .b(\PWMD/n24 ),
    .c(pnumcntD[1]),
    .d(\PWMD/pnumr [1]),
    .e(pwm_start_stop[29]),
    .o(\PWMD/n31 [1]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2793 (
    .a(\PWMD/n24 ),
    .b(\PWMD/n25_neg_lutinv ),
    .c(\PWMD/n26 [0]),
    .d(\PWMD/pnumr [0]),
    .o(_al_u2793_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2794 (
    .a(_al_u2793_o),
    .b(\PWMD/n24 ),
    .c(pnumcntD[0]),
    .d(\PWMD/pnumr [0]),
    .e(pwm_start_stop[29]),
    .o(\PWMD/n31 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u2795 (
    .a(\PWMD/FreCnt [12]),
    .b(\PWMD/FreCnt [8]),
    .c(\PWMD/FreCntr [13]),
    .d(\PWMD/FreCntr [9]),
    .o(_al_u2795_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*~C)*~(D*~B))"),
    .INIT(32'h80a088aa))
    _al_u2796 (
    .a(_al_u2795_o),
    .b(\PWMD/FreCnt [1]),
    .c(\PWMD/FreCnt [7]),
    .d(\PWMD/FreCntr [2]),
    .e(\PWMD/FreCntr [8]),
    .o(_al_u2796_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*C)*~(D@B))"),
    .INIT(32'h88220802))
    _al_u2797 (
    .a(_al_u2796_o),
    .b(\PWMD/FreCnt [18]),
    .c(\PWMD/FreCnt [7]),
    .d(\PWMD/FreCntr [19]),
    .e(\PWMD/FreCntr [8]),
    .o(_al_u2797_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C@B)*~(D@A))"),
    .INIT(16'h8241))
    _al_u2798 (
    .a(\PWMD/FreCnt [22]),
    .b(\PWMD/FreCnt [9]),
    .c(\PWMD/FreCntr [10]),
    .d(\PWMD/FreCntr [23]),
    .o(_al_u2798_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u2799 (
    .a(\PWMD/FreCnt [15]),
    .b(\PWMD/FreCnt [19]),
    .c(\PWMD/FreCntr [16]),
    .d(\PWMD/FreCntr [20]),
    .o(_al_u2799_o));
  EF2_PHY_SPAD #(
    //.LOCATION("P106"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("16"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u28 (
    .do({open_n870,dir_pad[10]}),
    .ts(1'b1),
    .opad(dir[10]));  // CPLD_SOC_AHB_TOP.v(7)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u280 (
    .a(\PWM2/pnumr [12]),
    .b(pnum2[12]),
    .c(pnum2[32]),
    .d(pwm_start_stop[18]),
    .o(\PWM2/n23 [12]));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u2800 (
    .a(_al_u2797_o),
    .b(_al_u2798_o),
    .c(_al_u2799_o),
    .d(\PWMD/FreCnt [11]),
    .e(\PWMD/FreCntr [12]),
    .o(_al_u2800_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u2801 (
    .a(\PWMD/FreCnt [4]),
    .b(\PWMD/FreCnt [6]),
    .c(\PWMD/FreCntr [5]),
    .d(\PWMD/FreCntr [7]),
    .o(_al_u2801_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u2802 (
    .a(_al_u2801_o),
    .b(\PWMD/FreCnt [24]),
    .c(\PWMD/FreCntr [25]),
    .o(_al_u2802_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u2803 (
    .a(\PWMD/FreCnt [16]),
    .b(\PWMD/FreCnt [2]),
    .c(\PWMD/FreCntr [17]),
    .d(\PWMD/FreCntr [3]),
    .o(_al_u2803_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u2804 (
    .a(_al_u2803_o),
    .b(\PWMD/FreCnt [25]),
    .c(\PWMD/FreCnt [5]),
    .d(\PWMD/FreCntr [26]),
    .e(\PWMD/FreCntr [6]),
    .o(_al_u2804_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u2805 (
    .a(\PWMD/FreCnt [17]),
    .b(\PWMD/FreCnt [23]),
    .c(\PWMD/FreCntr [18]),
    .d(\PWMD/FreCntr [24]),
    .o(_al_u2805_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~D*C)*~(~E*B))"),
    .INIT(32'haa0a2202))
    _al_u2806 (
    .a(_al_u2805_o),
    .b(\PWMD/FreCnt [1]),
    .c(\PWMD/FreCnt [13]),
    .d(\PWMD/FreCntr [14]),
    .e(\PWMD/FreCntr [2]),
    .o(_al_u2806_o));
  AL_MAP_LUT5 #(
    .EQN("(~B*~(E@C)*~(D*~A))"),
    .INIT(32'h20300203))
    _al_u2807 (
    .a(\PWMD/FreCnt [13]),
    .b(\PWMD/FreCnt [26]),
    .c(\PWMD/FreCnt [3]),
    .d(\PWMD/FreCntr [14]),
    .e(\PWMD/FreCntr [4]),
    .o(_al_u2807_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u2808 (
    .a(_al_u2802_o),
    .b(_al_u2804_o),
    .c(_al_u2806_o),
    .d(_al_u2807_o),
    .o(_al_u2808_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2809 (
    .a(\PWMD/FreCnt [17]),
    .b(\PWMD/FreCntr [18]),
    .o(_al_u2809_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u281 (
    .a(\PWM2/pnumr [11]),
    .b(pnum2[11]),
    .c(pnum2[32]),
    .d(pwm_start_stop[18]),
    .o(\PWM2/n23 [11]));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(~E*C)*~(D@B))"),
    .INIT(32'h44110401))
    _al_u2810 (
    .a(_al_u2809_o),
    .b(\PWMD/FreCnt [10]),
    .c(\PWMD/FreCnt [12]),
    .d(\PWMD/FreCntr [11]),
    .e(\PWMD/FreCntr [13]),
    .o(_al_u2810_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u2811 (
    .a(\PWMD/FreCnt [15]),
    .b(\PWMD/FreCnt [19]),
    .c(\PWMD/FreCntr [16]),
    .d(\PWMD/FreCntr [20]),
    .o(_al_u2811_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D@C))"),
    .INIT(16'h8008))
    _al_u2812 (
    .a(_al_u2810_o),
    .b(_al_u2811_o),
    .c(\PWMD/FreCnt [20]),
    .d(\PWMD/FreCntr [21]),
    .o(_al_u2812_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2813 (
    .a(\PWMD/FreCnt [8]),
    .b(\PWMD/FreCntr [9]),
    .o(_al_u2813_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(E@C)*~(D*~B))"),
    .INIT(32'h40500405))
    _al_u2814 (
    .a(_al_u2813_o),
    .b(\PWMD/FreCnt [0]),
    .c(\PWMD/FreCnt [21]),
    .d(\PWMD/FreCntr [1]),
    .e(\PWMD/FreCntr [22]),
    .o(_al_u2814_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2815 (
    .a(\PWMD/FreCnt [0]),
    .b(\PWMD/FreCntr [1]),
    .o(_al_u2815_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(~E*C)*~(D@B))"),
    .INIT(32'h44110401))
    _al_u2816 (
    .a(_al_u2815_o),
    .b(\PWMD/FreCnt [14]),
    .c(\PWMD/FreCnt [23]),
    .d(\PWMD/FreCntr [15]),
    .e(\PWMD/FreCntr [24]),
    .o(_al_u2816_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    _al_u2817 (
    .a(_al_u2800_o),
    .b(_al_u2808_o),
    .c(_al_u2812_o),
    .d(_al_u2814_o),
    .e(_al_u2816_o),
    .o(_al_u2817_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2818 (
    .a(_al_u2817_o),
    .b(pwm_state_read[13]),
    .o(\PWMD/u14_sel_is_1_o ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2819 (
    .a(\PWME/n0_lutinv ),
    .b(pwm_state_read[14]),
    .o(\PWME/n24 ));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u282 (
    .a(\PWM2/pnumr [10]),
    .b(pnum2[10]),
    .c(pnum2[32]),
    .d(pwm_start_stop[18]),
    .o(\PWM2/n23 [10]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u2820 (
    .a(pnumcntE[18]),
    .b(pnumcntE[19]),
    .c(pnumcntE[1]),
    .d(pnumcntE[20]),
    .o(_al_u2820_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u2821 (
    .a(_al_u2820_o),
    .b(pnumcntE[21]),
    .c(pnumcntE[22]),
    .d(pnumcntE[23]),
    .e(pnumcntE[2]),
    .o(_al_u2821_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u2822 (
    .a(_al_u2821_o),
    .b(pnumcntE[6]),
    .c(pnumcntE[7]),
    .d(pnumcntE[8]),
    .e(pnumcntE[9]),
    .o(_al_u2822_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u2823 (
    .a(pnumcntE[10]),
    .b(pnumcntE[11]),
    .c(pnumcntE[12]),
    .d(pnumcntE[13]),
    .o(_al_u2823_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u2824 (
    .a(_al_u2823_o),
    .b(pnumcntE[14]),
    .c(pnumcntE[15]),
    .d(pnumcntE[16]),
    .e(pnumcntE[17]),
    .o(_al_u2824_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u2825 (
    .a(pnumcntE[3]),
    .b(pnumcntE[4]),
    .c(pnumcntE[5]),
    .o(_al_u2825_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u2826 (
    .a(_al_u2822_o),
    .b(_al_u2824_o),
    .c(_al_u2825_o),
    .d(pnumcntE[0]),
    .o(\PWME/n25_neg_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2827 (
    .a(\PWME/n24 ),
    .b(\PWME/n25_neg_lutinv ),
    .c(\PWME/n26 [9]),
    .d(\PWME/pnumr [9]),
    .o(_al_u2827_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2828 (
    .a(_al_u2827_o),
    .b(\PWME/n24 ),
    .c(pnumcntE[9]),
    .d(\PWME/pnumr [9]),
    .e(pwm_start_stop[30]),
    .o(\PWME/n31 [9]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2829 (
    .a(\PWME/n24 ),
    .b(\PWME/n25_neg_lutinv ),
    .c(\PWME/n26 [8]),
    .d(\PWME/pnumr [8]),
    .o(_al_u2829_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u283 (
    .a(\PWM2/pnumr [1]),
    .b(pnum2[1]),
    .c(pnum2[32]),
    .d(pwm_start_stop[18]),
    .o(\PWM2/n23 [1]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2830 (
    .a(_al_u2829_o),
    .b(\PWME/n24 ),
    .c(pnumcntE[8]),
    .d(\PWME/pnumr [8]),
    .e(pwm_start_stop[30]),
    .o(\PWME/n31 [8]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2831 (
    .a(\PWME/n24 ),
    .b(\PWME/n25_neg_lutinv ),
    .c(\PWME/n26 [7]),
    .d(\PWME/pnumr [7]),
    .o(_al_u2831_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2832 (
    .a(_al_u2831_o),
    .b(\PWME/n24 ),
    .c(pnumcntE[7]),
    .d(\PWME/pnumr [7]),
    .e(pwm_start_stop[30]),
    .o(\PWME/n31 [7]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2833 (
    .a(\PWME/n24 ),
    .b(\PWME/n25_neg_lutinv ),
    .c(\PWME/n26 [6]),
    .d(\PWME/pnumr [6]),
    .o(_al_u2833_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2834 (
    .a(_al_u2833_o),
    .b(\PWME/n24 ),
    .c(pnumcntE[6]),
    .d(\PWME/pnumr [6]),
    .e(pwm_start_stop[30]),
    .o(\PWME/n31 [6]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2835 (
    .a(\PWME/n24 ),
    .b(\PWME/n25_neg_lutinv ),
    .c(\PWME/n26 [5]),
    .d(\PWME/pnumr [5]),
    .o(_al_u2835_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2836 (
    .a(_al_u2835_o),
    .b(\PWME/n24 ),
    .c(pnumcntE[5]),
    .d(\PWME/pnumr [5]),
    .e(pwm_start_stop[30]),
    .o(\PWME/n31 [5]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2837 (
    .a(\PWME/n24 ),
    .b(\PWME/n25_neg_lutinv ),
    .c(\PWME/n26 [4]),
    .d(\PWME/pnumr [4]),
    .o(_al_u2837_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2838 (
    .a(_al_u2837_o),
    .b(\PWME/n24 ),
    .c(pnumcntE[4]),
    .d(\PWME/pnumr [4]),
    .e(pwm_start_stop[30]),
    .o(\PWME/n31 [4]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2839 (
    .a(\PWME/n24 ),
    .b(\PWME/n25_neg_lutinv ),
    .c(\PWME/n26 [3]),
    .d(\PWME/pnumr [3]),
    .o(_al_u2839_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u284 (
    .a(\PWM2/pnumr [0]),
    .b(pnum2[0]),
    .c(pnum2[32]),
    .d(pwm_start_stop[18]),
    .o(\PWM2/n23 [0]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2840 (
    .a(_al_u2839_o),
    .b(\PWME/n24 ),
    .c(pnumcntE[3]),
    .d(\PWME/pnumr [3]),
    .e(pwm_start_stop[30]),
    .o(\PWME/n31 [3]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2841 (
    .a(\PWME/n24 ),
    .b(\PWME/n25_neg_lutinv ),
    .c(\PWME/n26 [23]),
    .d(\PWME/pnumr [23]),
    .o(_al_u2841_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2842 (
    .a(_al_u2841_o),
    .b(\PWME/n24 ),
    .c(pnumcntE[23]),
    .d(\PWME/pnumr [23]),
    .e(pwm_start_stop[30]),
    .o(\PWME/n31 [23]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2843 (
    .a(\PWME/n24 ),
    .b(\PWME/n25_neg_lutinv ),
    .c(\PWME/n26 [22]),
    .d(\PWME/pnumr [22]),
    .o(_al_u2843_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2844 (
    .a(_al_u2843_o),
    .b(\PWME/n24 ),
    .c(pnumcntE[22]),
    .d(\PWME/pnumr [22]),
    .e(pwm_start_stop[30]),
    .o(\PWME/n31 [22]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2845 (
    .a(\PWME/n24 ),
    .b(\PWME/n25_neg_lutinv ),
    .c(\PWME/n26 [21]),
    .d(\PWME/pnumr [21]),
    .o(_al_u2845_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2846 (
    .a(_al_u2845_o),
    .b(\PWME/n24 ),
    .c(pnumcntE[21]),
    .d(\PWME/pnumr [21]),
    .e(pwm_start_stop[30]),
    .o(\PWME/n31 [21]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2847 (
    .a(\PWME/n24 ),
    .b(\PWME/n25_neg_lutinv ),
    .c(\PWME/n26 [20]),
    .d(\PWME/pnumr [20]),
    .o(_al_u2847_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2848 (
    .a(_al_u2847_o),
    .b(\PWME/n24 ),
    .c(pnumcntE[20]),
    .d(\PWME/pnumr [20]),
    .e(pwm_start_stop[30]),
    .o(\PWME/n31 [20]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2849 (
    .a(\PWME/n24 ),
    .b(\PWME/n25_neg_lutinv ),
    .c(\PWME/n26 [2]),
    .d(\PWME/pnumr [2]),
    .o(_al_u2849_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u285 (
    .a(\PWM3/pnumr [9]),
    .b(pnum3[32]),
    .c(pnum3[9]),
    .d(pwm_start_stop[19]),
    .o(\PWM3/n23 [9]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2850 (
    .a(_al_u2849_o),
    .b(\PWME/n24 ),
    .c(pnumcntE[2]),
    .d(\PWME/pnumr [2]),
    .e(pwm_start_stop[30]),
    .o(\PWME/n31 [2]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2851 (
    .a(\PWME/n24 ),
    .b(\PWME/n25_neg_lutinv ),
    .c(\PWME/n26 [19]),
    .d(\PWME/pnumr [19]),
    .o(_al_u2851_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2852 (
    .a(_al_u2851_o),
    .b(\PWME/n24 ),
    .c(pnumcntE[19]),
    .d(\PWME/pnumr [19]),
    .e(pwm_start_stop[30]),
    .o(\PWME/n31 [19]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2853 (
    .a(\PWME/n24 ),
    .b(\PWME/n25_neg_lutinv ),
    .c(\PWME/n26 [18]),
    .d(\PWME/pnumr [18]),
    .o(_al_u2853_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2854 (
    .a(_al_u2853_o),
    .b(\PWME/n24 ),
    .c(pnumcntE[18]),
    .d(\PWME/pnumr [18]),
    .e(pwm_start_stop[30]),
    .o(\PWME/n31 [18]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2855 (
    .a(\PWME/n24 ),
    .b(\PWME/n25_neg_lutinv ),
    .c(\PWME/n26 [17]),
    .d(\PWME/pnumr [17]),
    .o(_al_u2855_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2856 (
    .a(_al_u2855_o),
    .b(\PWME/n24 ),
    .c(pnumcntE[17]),
    .d(\PWME/pnumr [17]),
    .e(pwm_start_stop[30]),
    .o(\PWME/n31 [17]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2857 (
    .a(\PWME/n24 ),
    .b(\PWME/n25_neg_lutinv ),
    .c(\PWME/n26 [16]),
    .d(\PWME/pnumr [16]),
    .o(_al_u2857_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2858 (
    .a(_al_u2857_o),
    .b(\PWME/n24 ),
    .c(pnumcntE[16]),
    .d(\PWME/pnumr [16]),
    .e(pwm_start_stop[30]),
    .o(\PWME/n31 [16]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2859 (
    .a(\PWME/n24 ),
    .b(\PWME/n25_neg_lutinv ),
    .c(\PWME/n26 [15]),
    .d(\PWME/pnumr [15]),
    .o(_al_u2859_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u286 (
    .a(\PWM3/pnumr [8]),
    .b(pnum3[32]),
    .c(pnum3[8]),
    .d(pwm_start_stop[19]),
    .o(\PWM3/n23 [8]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2860 (
    .a(_al_u2859_o),
    .b(\PWME/n24 ),
    .c(pnumcntE[15]),
    .d(\PWME/pnumr [15]),
    .e(pwm_start_stop[30]),
    .o(\PWME/n31 [15]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2861 (
    .a(\PWME/n24 ),
    .b(\PWME/n25_neg_lutinv ),
    .c(\PWME/n26 [14]),
    .d(\PWME/pnumr [14]),
    .o(_al_u2861_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2862 (
    .a(_al_u2861_o),
    .b(\PWME/n24 ),
    .c(pnumcntE[14]),
    .d(\PWME/pnumr [14]),
    .e(pwm_start_stop[30]),
    .o(\PWME/n31 [14]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2863 (
    .a(\PWME/n24 ),
    .b(\PWME/n25_neg_lutinv ),
    .c(\PWME/n26 [13]),
    .d(\PWME/pnumr [13]),
    .o(_al_u2863_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2864 (
    .a(_al_u2863_o),
    .b(\PWME/n24 ),
    .c(pnumcntE[13]),
    .d(\PWME/pnumr [13]),
    .e(pwm_start_stop[30]),
    .o(\PWME/n31 [13]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2865 (
    .a(\PWME/n24 ),
    .b(\PWME/n25_neg_lutinv ),
    .c(\PWME/n26 [12]),
    .d(\PWME/pnumr [12]),
    .o(_al_u2865_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2866 (
    .a(_al_u2865_o),
    .b(\PWME/n24 ),
    .c(pnumcntE[12]),
    .d(\PWME/pnumr [12]),
    .e(pwm_start_stop[30]),
    .o(\PWME/n31 [12]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2867 (
    .a(\PWME/n24 ),
    .b(\PWME/n25_neg_lutinv ),
    .c(\PWME/n26 [11]),
    .d(\PWME/pnumr [11]),
    .o(_al_u2867_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2868 (
    .a(_al_u2867_o),
    .b(\PWME/n24 ),
    .c(pnumcntE[11]),
    .d(\PWME/pnumr [11]),
    .e(pwm_start_stop[30]),
    .o(\PWME/n31 [11]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2869 (
    .a(\PWME/n24 ),
    .b(\PWME/n25_neg_lutinv ),
    .c(\PWME/n26 [10]),
    .d(\PWME/pnumr [10]),
    .o(_al_u2869_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u287 (
    .a(\PWM3/pnumr [7]),
    .b(pnum3[32]),
    .c(pnum3[7]),
    .d(pwm_start_stop[19]),
    .o(\PWM3/n23 [7]));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2870 (
    .a(_al_u2869_o),
    .b(\PWME/n24 ),
    .c(pnumcntE[10]),
    .d(\PWME/pnumr [10]),
    .e(pwm_start_stop[30]),
    .o(\PWME/n31 [10]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2871 (
    .a(\PWME/n24 ),
    .b(\PWME/n25_neg_lutinv ),
    .c(\PWME/n26 [1]),
    .d(\PWME/pnumr [1]),
    .o(_al_u2871_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2872 (
    .a(_al_u2871_o),
    .b(\PWME/n24 ),
    .c(pnumcntE[1]),
    .d(\PWME/pnumr [1]),
    .e(pwm_start_stop[30]),
    .o(\PWME/n31 [1]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2873 (
    .a(\PWME/n24 ),
    .b(\PWME/n25_neg_lutinv ),
    .c(\PWME/n26 [0]),
    .d(\PWME/pnumr [0]),
    .o(_al_u2873_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2874 (
    .a(_al_u2873_o),
    .b(\PWME/n24 ),
    .c(pnumcntE[0]),
    .d(\PWME/pnumr [0]),
    .e(pwm_start_stop[30]),
    .o(\PWME/n31 [0]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2875 (
    .a(\PWME/FreCnt [5]),
    .b(\PWME/FreCntr [6]),
    .o(_al_u2875_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(~E*C)*~(D@B))"),
    .INIT(32'h44110401))
    _al_u2876 (
    .a(_al_u2875_o),
    .b(\PWME/FreCnt [12]),
    .c(\PWME/FreCnt [23]),
    .d(\PWME/FreCntr [13]),
    .e(\PWME/FreCntr [24]),
    .o(_al_u2876_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(~D*B))"),
    .INIT(32'ha0200a02))
    _al_u2877 (
    .a(_al_u2876_o),
    .b(\PWME/FreCnt [10]),
    .c(\PWME/FreCnt [24]),
    .d(\PWME/FreCntr [11]),
    .e(\PWME/FreCntr [25]),
    .o(_al_u2877_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u2878 (
    .a(\PWME/FreCnt [3]),
    .b(\PWME/FreCnt [5]),
    .c(\PWME/FreCntr [4]),
    .d(\PWME/FreCntr [6]),
    .o(_al_u2878_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u2879 (
    .a(\PWME/FreCnt [0]),
    .b(\PWME/FreCnt [14]),
    .c(\PWME/FreCntr [1]),
    .d(\PWME/FreCntr [15]),
    .o(_al_u2879_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u288 (
    .a(\PWM3/pnumr [6]),
    .b(pnum3[32]),
    .c(pnum3[6]),
    .d(pwm_start_stop[19]),
    .o(\PWM3/n23 [6]));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u2880 (
    .a(_al_u2877_o),
    .b(_al_u2878_o),
    .c(_al_u2879_o),
    .d(\PWME/FreCnt [9]),
    .e(\PWME/FreCntr [10]),
    .o(_al_u2880_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2881 (
    .a(\PWME/FreCnt [17]),
    .b(\PWME/FreCntr [18]),
    .o(_al_u2881_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(E@C)*~(D*~B))"),
    .INIT(32'h40500405))
    _al_u2882 (
    .a(_al_u2881_o),
    .b(\PWME/FreCnt [21]),
    .c(\PWME/FreCnt [8]),
    .d(\PWME/FreCntr [22]),
    .e(\PWME/FreCntr [9]),
    .o(_al_u2882_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u2883 (
    .a(\PWME/FreCnt [15]),
    .b(\PWME/FreCnt [3]),
    .c(\PWME/FreCntr [16]),
    .d(\PWME/FreCntr [4]),
    .o(_al_u2883_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D@C))"),
    .INIT(16'h8008))
    _al_u2884 (
    .a(_al_u2882_o),
    .b(_al_u2883_o),
    .c(\PWME/FreCnt [16]),
    .d(\PWME/FreCntr [17]),
    .o(_al_u2884_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(D*~A))"),
    .INIT(16'h8acf))
    _al_u2885 (
    .a(\PWME/FreCnt [1]),
    .b(\PWME/FreCnt [15]),
    .c(\PWME/FreCntr [16]),
    .d(\PWME/FreCntr [2]),
    .o(_al_u2885_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*C)*~(D*~B))"),
    .INIT(32'h88aa080a))
    _al_u2886 (
    .a(_al_u2885_o),
    .b(\PWME/FreCnt [10]),
    .c(\PWME/FreCnt [19]),
    .d(\PWME/FreCntr [11]),
    .e(\PWME/FreCntr [20]),
    .o(_al_u2886_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u2887 (
    .a(\PWME/FreCnt [13]),
    .b(\PWME/FreCnt [21]),
    .c(\PWME/FreCntr [14]),
    .d(\PWME/FreCntr [22]),
    .o(_al_u2887_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u2888 (
    .a(_al_u2884_o),
    .b(_al_u2886_o),
    .c(_al_u2887_o),
    .d(\PWME/FreCnt [11]),
    .e(\PWME/FreCntr [12]),
    .o(_al_u2888_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u2889 (
    .a(\PWME/FreCnt [22]),
    .b(\PWME/FreCnt [4]),
    .c(\PWME/FreCntr [23]),
    .d(\PWME/FreCntr [5]),
    .o(_al_u2889_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u289 (
    .a(\PWM3/pnumr [5]),
    .b(pnum3[32]),
    .c(pnum3[5]),
    .d(pwm_start_stop[19]),
    .o(\PWM3/n23 [5]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u2890 (
    .a(_al_u2889_o),
    .b(\PWME/FreCnt [6]),
    .c(\PWME/FreCntr [7]),
    .o(_al_u2890_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C@B)*~(D@A))"),
    .INIT(16'h8241))
    _al_u2891 (
    .a(\PWME/FreCnt [2]),
    .b(\PWME/FreCnt [20]),
    .c(\PWME/FreCntr [21]),
    .d(\PWME/FreCntr [3]),
    .o(_al_u2891_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u2892 (
    .a(_al_u2891_o),
    .b(\PWME/FreCnt [18]),
    .c(\PWME/FreCnt [25]),
    .d(\PWME/FreCntr [19]),
    .e(\PWME/FreCntr [26]),
    .o(_al_u2892_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u2893 (
    .a(\PWME/FreCnt [17]),
    .b(\PWME/FreCnt [23]),
    .c(\PWME/FreCntr [18]),
    .d(\PWME/FreCntr [24]),
    .o(_al_u2893_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*~C)*~(~D*B))"),
    .INIT(32'ha020aa22))
    _al_u2894 (
    .a(_al_u2893_o),
    .b(\PWME/FreCnt [1]),
    .c(\PWME/FreCnt [19]),
    .d(\PWME/FreCntr [2]),
    .e(\PWME/FreCntr [20]),
    .o(_al_u2894_o));
  AL_MAP_LUT5 #(
    .EQN("(~B*~(E@C)*~(~D*A))"),
    .INIT(32'h30100301))
    _al_u2895 (
    .a(\PWME/FreCnt [13]),
    .b(\PWME/FreCnt [26]),
    .c(\PWME/FreCnt [7]),
    .d(\PWME/FreCntr [14]),
    .e(\PWME/FreCntr [8]),
    .o(_al_u2895_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u2896 (
    .a(_al_u2890_o),
    .b(_al_u2892_o),
    .c(_al_u2894_o),
    .d(_al_u2895_o),
    .o(_al_u2896_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*A))"),
    .INIT(16'h7f00))
    _al_u2897 (
    .a(_al_u2880_o),
    .b(_al_u2888_o),
    .c(_al_u2896_o),
    .d(pwm_state_read[14]),
    .o(\PWME/u14_sel_is_1_o ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u2898 (
    .a(\PWMF/n0_lutinv ),
    .b(pwm_state_read[15]),
    .o(\PWMF/n24 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u2899 (
    .a(pnumcntF[18]),
    .b(pnumcntF[19]),
    .c(pnumcntF[1]),
    .d(pnumcntF[20]),
    .o(_al_u2899_o));
  EF2_PHY_PAD #(
    //.LOCATION("P42"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u29 (
    .do({open_n878,open_n879,open_n880,dir_pad[9]}),
    .opad(dir[9]));  // CPLD_SOC_AHB_TOP.v(7)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u290 (
    .a(\PWM3/pnumr [4]),
    .b(pnum3[32]),
    .c(pnum3[4]),
    .d(pwm_start_stop[19]),
    .o(\PWM3/n23 [4]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u2900 (
    .a(_al_u2899_o),
    .b(pnumcntF[21]),
    .c(pnumcntF[22]),
    .d(pnumcntF[23]),
    .e(pnumcntF[2]),
    .o(_al_u2900_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u2901 (
    .a(_al_u2900_o),
    .b(pnumcntF[6]),
    .c(pnumcntF[7]),
    .d(pnumcntF[8]),
    .e(pnumcntF[9]),
    .o(_al_u2901_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u2902 (
    .a(pnumcntF[10]),
    .b(pnumcntF[11]),
    .c(pnumcntF[12]),
    .d(pnumcntF[13]),
    .o(_al_u2902_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u2903 (
    .a(_al_u2902_o),
    .b(pnumcntF[14]),
    .c(pnumcntF[15]),
    .d(pnumcntF[16]),
    .e(pnumcntF[17]),
    .o(_al_u2903_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u2904 (
    .a(pnumcntF[3]),
    .b(pnumcntF[4]),
    .c(pnumcntF[5]),
    .o(_al_u2904_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u2905 (
    .a(_al_u2901_o),
    .b(_al_u2903_o),
    .c(_al_u2904_o),
    .d(pnumcntF[0]),
    .o(\PWMF/n25_neg_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2906 (
    .a(\PWMF/n24 ),
    .b(\PWMF/n25_neg_lutinv ),
    .c(\PWMF/n26 [9]),
    .d(\PWMF/pnumr [9]),
    .o(_al_u2906_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2907 (
    .a(_al_u2906_o),
    .b(\PWMF/n24 ),
    .c(pnumcntF[9]),
    .d(\PWMF/pnumr [9]),
    .e(pwm_start_stop[31]),
    .o(\PWMF/n31 [9]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2908 (
    .a(\PWMF/n24 ),
    .b(\PWMF/n25_neg_lutinv ),
    .c(\PWMF/n26 [8]),
    .d(\PWMF/pnumr [8]),
    .o(_al_u2908_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2909 (
    .a(_al_u2908_o),
    .b(\PWMF/n24 ),
    .c(pnumcntF[8]),
    .d(\PWMF/pnumr [8]),
    .e(pwm_start_stop[31]),
    .o(\PWMF/n31 [8]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u291 (
    .a(\PWM3/pnumr [31]),
    .b(pnum3[31]),
    .c(pnum3[32]),
    .d(pwm_start_stop[19]),
    .o(\PWM3/n23 [31]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2910 (
    .a(\PWMF/n24 ),
    .b(\PWMF/n25_neg_lutinv ),
    .c(\PWMF/n26 [7]),
    .d(\PWMF/pnumr [7]),
    .o(_al_u2910_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2911 (
    .a(_al_u2910_o),
    .b(\PWMF/n24 ),
    .c(pnumcntF[7]),
    .d(\PWMF/pnumr [7]),
    .e(pwm_start_stop[31]),
    .o(\PWMF/n31 [7]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2912 (
    .a(\PWMF/n24 ),
    .b(\PWMF/n25_neg_lutinv ),
    .c(\PWMF/n26 [6]),
    .d(\PWMF/pnumr [6]),
    .o(_al_u2912_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2913 (
    .a(_al_u2912_o),
    .b(\PWMF/n24 ),
    .c(pnumcntF[6]),
    .d(\PWMF/pnumr [6]),
    .e(pwm_start_stop[31]),
    .o(\PWMF/n31 [6]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2914 (
    .a(\PWMF/n24 ),
    .b(\PWMF/n25_neg_lutinv ),
    .c(\PWMF/n26 [5]),
    .d(\PWMF/pnumr [5]),
    .o(_al_u2914_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2915 (
    .a(_al_u2914_o),
    .b(\PWMF/n24 ),
    .c(pnumcntF[5]),
    .d(\PWMF/pnumr [5]),
    .e(pwm_start_stop[31]),
    .o(\PWMF/n31 [5]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2916 (
    .a(\PWMF/n24 ),
    .b(\PWMF/n25_neg_lutinv ),
    .c(\PWMF/n26 [4]),
    .d(\PWMF/pnumr [4]),
    .o(_al_u2916_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2917 (
    .a(_al_u2916_o),
    .b(\PWMF/n24 ),
    .c(pnumcntF[4]),
    .d(\PWMF/pnumr [4]),
    .e(pwm_start_stop[31]),
    .o(\PWMF/n31 [4]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2918 (
    .a(\PWMF/n24 ),
    .b(\PWMF/n25_neg_lutinv ),
    .c(\PWMF/n26 [3]),
    .d(\PWMF/pnumr [3]),
    .o(_al_u2918_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2919 (
    .a(_al_u2918_o),
    .b(\PWMF/n24 ),
    .c(pnumcntF[3]),
    .d(\PWMF/pnumr [3]),
    .e(pwm_start_stop[31]),
    .o(\PWMF/n31 [3]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u292 (
    .a(\PWM3/pnumr [30]),
    .b(pnum3[30]),
    .c(pnum3[32]),
    .d(pwm_start_stop[19]),
    .o(\PWM3/n23 [30]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2920 (
    .a(\PWMF/n24 ),
    .b(\PWMF/n25_neg_lutinv ),
    .c(\PWMF/n26 [23]),
    .d(\PWMF/pnumr [23]),
    .o(_al_u2920_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2921 (
    .a(_al_u2920_o),
    .b(\PWMF/n24 ),
    .c(pnumcntF[23]),
    .d(\PWMF/pnumr [23]),
    .e(pwm_start_stop[31]),
    .o(\PWMF/n31 [23]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2922 (
    .a(\PWMF/n24 ),
    .b(\PWMF/n25_neg_lutinv ),
    .c(\PWMF/n26 [22]),
    .d(\PWMF/pnumr [22]),
    .o(_al_u2922_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2923 (
    .a(_al_u2922_o),
    .b(\PWMF/n24 ),
    .c(pnumcntF[22]),
    .d(\PWMF/pnumr [22]),
    .e(pwm_start_stop[31]),
    .o(\PWMF/n31 [22]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2924 (
    .a(\PWMF/n24 ),
    .b(\PWMF/n25_neg_lutinv ),
    .c(\PWMF/n26 [21]),
    .d(\PWMF/pnumr [21]),
    .o(_al_u2924_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2925 (
    .a(_al_u2924_o),
    .b(\PWMF/n24 ),
    .c(pnumcntF[21]),
    .d(\PWMF/pnumr [21]),
    .e(pwm_start_stop[31]),
    .o(\PWMF/n31 [21]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2926 (
    .a(\PWMF/n24 ),
    .b(\PWMF/n25_neg_lutinv ),
    .c(\PWMF/n26 [20]),
    .d(\PWMF/pnumr [20]),
    .o(_al_u2926_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2927 (
    .a(_al_u2926_o),
    .b(\PWMF/n24 ),
    .c(pnumcntF[20]),
    .d(\PWMF/pnumr [20]),
    .e(pwm_start_stop[31]),
    .o(\PWMF/n31 [20]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2928 (
    .a(\PWMF/n24 ),
    .b(\PWMF/n25_neg_lutinv ),
    .c(\PWMF/n26 [2]),
    .d(\PWMF/pnumr [2]),
    .o(_al_u2928_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2929 (
    .a(_al_u2928_o),
    .b(\PWMF/n24 ),
    .c(pnumcntF[2]),
    .d(\PWMF/pnumr [2]),
    .e(pwm_start_stop[31]),
    .o(\PWMF/n31 [2]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u293 (
    .a(\PWM3/pnumr [3]),
    .b(pnum3[3]),
    .c(pnum3[32]),
    .d(pwm_start_stop[19]),
    .o(\PWM3/n23 [3]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2930 (
    .a(\PWMF/n24 ),
    .b(\PWMF/n25_neg_lutinv ),
    .c(\PWMF/n26 [19]),
    .d(\PWMF/pnumr [19]),
    .o(_al_u2930_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2931 (
    .a(_al_u2930_o),
    .b(\PWMF/n24 ),
    .c(pnumcntF[19]),
    .d(\PWMF/pnumr [19]),
    .e(pwm_start_stop[31]),
    .o(\PWMF/n31 [19]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2932 (
    .a(\PWMF/n24 ),
    .b(\PWMF/n25_neg_lutinv ),
    .c(\PWMF/n26 [18]),
    .d(\PWMF/pnumr [18]),
    .o(_al_u2932_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2933 (
    .a(_al_u2932_o),
    .b(\PWMF/n24 ),
    .c(pnumcntF[18]),
    .d(\PWMF/pnumr [18]),
    .e(pwm_start_stop[31]),
    .o(\PWMF/n31 [18]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2934 (
    .a(\PWMF/n24 ),
    .b(\PWMF/n25_neg_lutinv ),
    .c(\PWMF/n26 [17]),
    .d(\PWMF/pnumr [17]),
    .o(_al_u2934_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2935 (
    .a(_al_u2934_o),
    .b(\PWMF/n24 ),
    .c(pnumcntF[17]),
    .d(\PWMF/pnumr [17]),
    .e(pwm_start_stop[31]),
    .o(\PWMF/n31 [17]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2936 (
    .a(\PWMF/n24 ),
    .b(\PWMF/n25_neg_lutinv ),
    .c(\PWMF/n26 [16]),
    .d(\PWMF/pnumr [16]),
    .o(_al_u2936_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2937 (
    .a(_al_u2936_o),
    .b(\PWMF/n24 ),
    .c(pnumcntF[16]),
    .d(\PWMF/pnumr [16]),
    .e(pwm_start_stop[31]),
    .o(\PWMF/n31 [16]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2938 (
    .a(\PWMF/n24 ),
    .b(\PWMF/n25_neg_lutinv ),
    .c(\PWMF/n26 [15]),
    .d(\PWMF/pnumr [15]),
    .o(_al_u2938_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2939 (
    .a(_al_u2938_o),
    .b(\PWMF/n24 ),
    .c(pnumcntF[15]),
    .d(\PWMF/pnumr [15]),
    .e(pwm_start_stop[31]),
    .o(\PWMF/n31 [15]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u294 (
    .a(\PWM3/pnumr [29]),
    .b(pnum3[29]),
    .c(pnum3[32]),
    .d(pwm_start_stop[19]),
    .o(\PWM3/n23 [29]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2940 (
    .a(\PWMF/n24 ),
    .b(\PWMF/n25_neg_lutinv ),
    .c(\PWMF/n26 [14]),
    .d(\PWMF/pnumr [14]),
    .o(_al_u2940_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2941 (
    .a(_al_u2940_o),
    .b(\PWMF/n24 ),
    .c(pnumcntF[14]),
    .d(\PWMF/pnumr [14]),
    .e(pwm_start_stop[31]),
    .o(\PWMF/n31 [14]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2942 (
    .a(\PWMF/n24 ),
    .b(\PWMF/n25_neg_lutinv ),
    .c(\PWMF/n26 [13]),
    .d(\PWMF/pnumr [13]),
    .o(_al_u2942_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2943 (
    .a(_al_u2942_o),
    .b(\PWMF/n24 ),
    .c(pnumcntF[13]),
    .d(\PWMF/pnumr [13]),
    .e(pwm_start_stop[31]),
    .o(\PWMF/n31 [13]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2944 (
    .a(\PWMF/n24 ),
    .b(\PWMF/n25_neg_lutinv ),
    .c(\PWMF/n26 [12]),
    .d(\PWMF/pnumr [12]),
    .o(_al_u2944_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2945 (
    .a(_al_u2944_o),
    .b(\PWMF/n24 ),
    .c(pnumcntF[12]),
    .d(\PWMF/pnumr [12]),
    .e(pwm_start_stop[31]),
    .o(\PWMF/n31 [12]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2946 (
    .a(\PWMF/n24 ),
    .b(\PWMF/n25_neg_lutinv ),
    .c(\PWMF/n26 [11]),
    .d(\PWMF/pnumr [11]),
    .o(_al_u2946_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2947 (
    .a(_al_u2946_o),
    .b(\PWMF/n24 ),
    .c(pnumcntF[11]),
    .d(\PWMF/pnumr [11]),
    .e(pwm_start_stop[31]),
    .o(\PWMF/n31 [11]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2948 (
    .a(\PWMF/n24 ),
    .b(\PWMF/n25_neg_lutinv ),
    .c(\PWMF/n26 [10]),
    .d(\PWMF/pnumr [10]),
    .o(_al_u2948_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2949 (
    .a(_al_u2948_o),
    .b(\PWMF/n24 ),
    .c(pnumcntF[10]),
    .d(\PWMF/pnumr [10]),
    .e(pwm_start_stop[31]),
    .o(\PWMF/n31 [10]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u295 (
    .a(\PWM3/pnumr [28]),
    .b(pnum3[28]),
    .c(pnum3[32]),
    .d(pwm_start_stop[19]),
    .o(\PWM3/n23 [28]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2950 (
    .a(\PWMF/n24 ),
    .b(\PWMF/n25_neg_lutinv ),
    .c(\PWMF/n26 [1]),
    .d(\PWMF/pnumr [1]),
    .o(_al_u2950_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2951 (
    .a(_al_u2950_o),
    .b(\PWMF/n24 ),
    .c(pnumcntF[1]),
    .d(\PWMF/pnumr [1]),
    .e(pwm_start_stop[31]),
    .o(\PWMF/n31 [1]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u2952 (
    .a(\PWMF/n24 ),
    .b(\PWMF/n25_neg_lutinv ),
    .c(\PWMF/n26 [0]),
    .d(\PWMF/pnumr [0]),
    .o(_al_u2952_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~A*~(C*~B))*~(D)*~(E)+~(~A*~(C*~B))*D*~(E)+~(~(~A*~(C*~B)))*D*E+~(~A*~(C*~B))*D*E)"),
    .INIT(32'hff00baba))
    _al_u2953 (
    .a(_al_u2952_o),
    .b(\PWMF/n24 ),
    .c(pnumcntF[0]),
    .d(\PWMF/pnumr [0]),
    .e(pwm_start_stop[31]),
    .o(\PWMF/n31 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u2954 (
    .a(\PWMF/FreCnt [14]),
    .b(\PWMF/FreCnt [5]),
    .c(\PWMF/FreCntr [15]),
    .d(\PWMF/FreCntr [6]),
    .o(_al_u2954_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C@B)*~(D@A))"),
    .INIT(16'h8241))
    _al_u2955 (
    .a(\PWMF/FreCnt [2]),
    .b(\PWMF/FreCnt [24]),
    .c(\PWMF/FreCntr [25]),
    .d(\PWMF/FreCntr [3]),
    .o(_al_u2955_o));
  AL_MAP_LUT5 #(
    .EQN("(~D*B*A*~(~E*C))"),
    .INIT(32'h00880008))
    _al_u2956 (
    .a(_al_u2954_o),
    .b(_al_u2955_o),
    .c(\PWMF/FreCnt [10]),
    .d(\PWMF/FreCnt [26]),
    .e(\PWMF/FreCntr [11]),
    .o(_al_u2956_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u2957 (
    .a(\PWMF/FreCnt [11]),
    .b(\PWMF/FreCnt [6]),
    .c(\PWMF/FreCntr [12]),
    .d(\PWMF/FreCntr [7]),
    .o(_al_u2957_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u2958 (
    .a(_al_u2957_o),
    .b(\PWMF/FreCnt [4]),
    .c(\PWMF/FreCntr [5]),
    .o(_al_u2958_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u2959 (
    .a(\PWMF/FreCnt [15]),
    .b(\PWMF/FreCnt [7]),
    .c(\PWMF/FreCntr [16]),
    .d(\PWMF/FreCntr [8]),
    .o(_al_u2959_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u296 (
    .a(\PWM3/pnumr [27]),
    .b(pnum3[27]),
    .c(pnum3[32]),
    .d(pwm_start_stop[19]),
    .o(\PWM3/n23 [27]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*~C)*~(~E*B))"),
    .INIT(32'ha0aa2022))
    _al_u2960 (
    .a(_al_u2959_o),
    .b(\PWMF/FreCnt [1]),
    .c(\PWMF/FreCnt [14]),
    .d(\PWMF/FreCntr [15]),
    .e(\PWMF/FreCntr [2]),
    .o(_al_u2960_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u2961 (
    .a(\PWMF/FreCnt [8]),
    .b(\PWMF/FreCntr [9]),
    .o(_al_u2961_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(E@C)*~(~D*B))"),
    .INIT(32'h50100501))
    _al_u2962 (
    .a(_al_u2961_o),
    .b(\PWMF/FreCnt [19]),
    .c(\PWMF/FreCnt [22]),
    .d(\PWMF/FreCntr [20]),
    .e(\PWMF/FreCntr [23]),
    .o(_al_u2962_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u2963 (
    .a(_al_u2956_o),
    .b(_al_u2958_o),
    .c(_al_u2960_o),
    .d(_al_u2962_o),
    .o(_al_u2963_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u2964 (
    .a(\PWMF/FreCnt [18]),
    .b(\PWMF/FreCnt [20]),
    .c(\PWMF/FreCntr [19]),
    .d(\PWMF/FreCntr [21]),
    .o(_al_u2964_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u2965 (
    .a(\PWMF/FreCnt [10]),
    .b(\PWMF/FreCnt [21]),
    .c(\PWMF/FreCntr [11]),
    .d(\PWMF/FreCntr [22]),
    .o(_al_u2965_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D@C))"),
    .INIT(16'h8008))
    _al_u2966 (
    .a(_al_u2964_o),
    .b(_al_u2965_o),
    .c(\PWMF/FreCnt [16]),
    .d(\PWMF/FreCntr [17]),
    .o(_al_u2966_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(~C*A))"),
    .INIT(16'hf531))
    _al_u2967 (
    .a(\PWMF/FreCnt [13]),
    .b(\PWMF/FreCnt [23]),
    .c(\PWMF/FreCntr [14]),
    .d(\PWMF/FreCntr [24]),
    .o(_al_u2967_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*~C)*~(~D*B))"),
    .INIT(32'ha020aa22))
    _al_u2968 (
    .a(_al_u2967_o),
    .b(\PWMF/FreCnt [3]),
    .c(\PWMF/FreCnt [7]),
    .d(\PWMF/FreCntr [4]),
    .e(\PWMF/FreCntr [8]),
    .o(_al_u2968_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(~C*A))"),
    .INIT(16'hc4f5))
    _al_u2969 (
    .a(\PWMF/FreCnt [15]),
    .b(\PWMF/FreCnt [25]),
    .c(\PWMF/FreCntr [16]),
    .d(\PWMF/FreCntr [26]),
    .o(_al_u2969_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u297 (
    .a(\PWM3/pnumr [26]),
    .b(pnum3[26]),
    .c(pnum3[32]),
    .d(pwm_start_stop[19]),
    .o(\PWM3/n23 [26]));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u2970 (
    .a(_al_u2966_o),
    .b(_al_u2968_o),
    .c(_al_u2969_o),
    .d(\PWMF/FreCnt [12]),
    .e(\PWMF/FreCntr [13]),
    .o(_al_u2970_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*~A))"),
    .INIT(16'h8caf))
    _al_u2971 (
    .a(\PWMF/FreCnt [23]),
    .b(\PWMF/FreCnt [3]),
    .c(\PWMF/FreCntr [24]),
    .d(\PWMF/FreCntr [4]),
    .o(_al_u2971_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*~C)*~(~E*B))"),
    .INIT(32'ha0aa2022))
    _al_u2972 (
    .a(_al_u2971_o),
    .b(\PWMF/FreCnt [25]),
    .c(\PWMF/FreCnt [9]),
    .d(\PWMF/FreCntr [10]),
    .e(\PWMF/FreCntr [26]),
    .o(_al_u2972_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*C)*~(D@B))"),
    .INIT(32'h88220802))
    _al_u2973 (
    .a(_al_u2972_o),
    .b(\PWMF/FreCnt [0]),
    .c(\PWMF/FreCnt [5]),
    .d(\PWMF/FreCntr [1]),
    .e(\PWMF/FreCntr [6]),
    .o(_al_u2973_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(D*~A))"),
    .INIT(16'ha2f3))
    _al_u2974 (
    .a(\PWMF/FreCnt [8]),
    .b(\PWMF/FreCnt [9]),
    .c(\PWMF/FreCntr [10]),
    .d(\PWMF/FreCntr [9]),
    .o(_al_u2974_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*~C)*~(D*~B))"),
    .INIT(32'h80a088aa))
    _al_u2975 (
    .a(_al_u2974_o),
    .b(\PWMF/FreCnt [13]),
    .c(\PWMF/FreCnt [17]),
    .d(\PWMF/FreCntr [14]),
    .e(\PWMF/FreCntr [18]),
    .o(_al_u2975_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*B)*~(C*~A))"),
    .INIT(16'haf23))
    _al_u2976 (
    .a(\PWMF/FreCnt [1]),
    .b(\PWMF/FreCnt [21]),
    .c(\PWMF/FreCntr [2]),
    .d(\PWMF/FreCntr [22]),
    .o(_al_u2976_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*~C)*~(~D*B))"),
    .INIT(32'ha020aa22))
    _al_u2977 (
    .a(_al_u2976_o),
    .b(\PWMF/FreCnt [17]),
    .c(\PWMF/FreCnt [19]),
    .d(\PWMF/FreCntr [18]),
    .e(\PWMF/FreCntr [20]),
    .o(_al_u2977_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    _al_u2978 (
    .a(_al_u2963_o),
    .b(_al_u2970_o),
    .c(_al_u2973_o),
    .d(_al_u2975_o),
    .e(_al_u2977_o),
    .o(_al_u2978_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2979 (
    .a(_al_u2978_o),
    .b(pwm_state_read[15]),
    .o(\PWMF/u14_sel_is_1_o ));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u298 (
    .a(\PWM3/pnumr [25]),
    .b(pnum3[25]),
    .c(pnum3[32]),
    .d(pwm_start_stop[19]),
    .o(\PWM3/n23 [25]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*~A)"),
    .INIT(16'h4000))
    _al_u2980 (
    .a(timer[12]),
    .b(timer[13]),
    .c(timer[14]),
    .d(timer[15]),
    .o(_al_u2980_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*D*~C*B*A)"),
    .INIT(32'h00000800))
    _al_u2981 (
    .a(_al_u2980_o),
    .b(timer[16]),
    .c(timer[17]),
    .d(timer[18]),
    .e(timer[19]),
    .o(_al_u2981_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*D*~C*B*A)"),
    .INIT(32'h00000800))
    _al_u2982 (
    .a(_al_u2981_o),
    .b(timer[24]),
    .c(timer[25]),
    .d(timer[26]),
    .e(timer[27]),
    .o(_al_u2982_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u2983 (
    .a(_al_u2982_o),
    .b(_al_u1640_o),
    .c(_al_u1648_o),
    .o(_al_u2983_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u2984 (
    .a(_al_u2983_o),
    .b(n4_neg),
    .o(_al_u2984_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u2985 (
    .a(timer[14]),
    .b(timer[15]),
    .c(timer[26]),
    .d(timer[27]),
    .o(_al_u2985_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*B*A)"),
    .INIT(32'h00000008))
    _al_u2986 (
    .a(_al_u2985_o),
    .b(timer[12]),
    .c(timer[13]),
    .d(timer[16]),
    .e(timer[17]),
    .o(_al_u2986_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u2987 (
    .a(_al_u1639_o),
    .b(timer[18]),
    .c(timer[19]),
    .d(timer[24]),
    .e(timer[25]),
    .o(_al_u2987_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u2988 (
    .a(_al_u1647_o),
    .b(_al_u1642_o),
    .c(_al_u2986_o),
    .d(_al_u2987_o),
    .o(_al_u2988_o));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(~C*~(~D*~B)))"),
    .INIT(16'h5f5d))
    _al_u2989 (
    .a(_al_u2984_o),
    .b(_al_u1652_o),
    .c(_al_u2988_o),
    .d(ledout_pad[2]),
    .o(n10[2]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u299 (
    .a(\PWM3/pnumr [24]),
    .b(pnum3[24]),
    .c(pnum3[32]),
    .d(pwm_start_stop[19]),
    .o(\PWM3/n23 [24]));
  AL_MAP_LUT5 #(
    .EQN("(D*~(C)*~((~E*~(B*A)))+D*C*~((~E*~(B*A)))+~(D)*C*(~E*~(B*A))+D*C*(~E*~(B*A)))"),
    .INIT(32'hff00f870))
    _al_u2990 (
    .a(\PWM0/n24 ),
    .b(\PWM0/n25_neg_lutinv ),
    .c(dir_pad[0]),
    .d(\PWM0/pnumr [31]),
    .e(pwm_start_stop[16]),
    .o(\PWM0/n32 ));
  AL_MAP_LUT5 #(
    .EQN("(D*~(C)*~((~E*~(B*A)))+D*C*~((~E*~(B*A)))+~(D)*C*(~E*~(B*A))+D*C*(~E*~(B*A)))"),
    .INIT(32'hff00f870))
    _al_u2991 (
    .a(\PWM1/n24 ),
    .b(\PWM1/n25_neg_lutinv ),
    .c(dir_pad[1]),
    .d(\PWM1/pnumr [31]),
    .e(pwm_start_stop[17]),
    .o(\PWM1/n32 ));
  AL_MAP_LUT5 #(
    .EQN("(D*~(C)*~((~E*~(B*A)))+D*C*~((~E*~(B*A)))+~(D)*C*(~E*~(B*A))+D*C*(~E*~(B*A)))"),
    .INIT(32'hff00f870))
    _al_u2992 (
    .a(\PWM2/n24 ),
    .b(\PWM2/n25_neg_lutinv ),
    .c(dir_pad[2]),
    .d(\PWM2/pnumr [31]),
    .e(pwm_start_stop[18]),
    .o(\PWM2/n32 ));
  AL_MAP_LUT5 #(
    .EQN("(D*~(C)*~((~E*~(B*A)))+D*C*~((~E*~(B*A)))+~(D)*C*(~E*~(B*A))+D*C*(~E*~(B*A)))"),
    .INIT(32'hff00f870))
    _al_u2993 (
    .a(\PWM3/n24 ),
    .b(\PWM3/n25_neg_lutinv ),
    .c(dir_pad[3]),
    .d(\PWM3/pnumr [31]),
    .e(pwm_start_stop[19]),
    .o(\PWM3/n32 ));
  AL_MAP_LUT5 #(
    .EQN("(D*~(C)*~((~E*~(B*A)))+D*C*~((~E*~(B*A)))+~(D)*C*(~E*~(B*A))+D*C*(~E*~(B*A)))"),
    .INIT(32'hff00f870))
    _al_u2994 (
    .a(\PWM4/n24 ),
    .b(\PWM4/n25_neg_lutinv ),
    .c(dir_pad[4]),
    .d(\PWM4/pnumr [31]),
    .e(pwm_start_stop[20]),
    .o(\PWM4/n32 ));
  AL_MAP_LUT5 #(
    .EQN("(D*~(C)*~((~E*~(B*A)))+D*C*~((~E*~(B*A)))+~(D)*C*(~E*~(B*A))+D*C*(~E*~(B*A)))"),
    .INIT(32'hff00f870))
    _al_u2995 (
    .a(\PWM5/n24 ),
    .b(\PWM5/n25_neg_lutinv ),
    .c(dir_pad[5]),
    .d(\PWM5/pnumr [31]),
    .e(pwm_start_stop[21]),
    .o(\PWM5/n32 ));
  AL_MAP_LUT5 #(
    .EQN("(D*~(C)*~((~E*~(B*A)))+D*C*~((~E*~(B*A)))+~(D)*C*(~E*~(B*A))+D*C*(~E*~(B*A)))"),
    .INIT(32'hff00f870))
    _al_u2996 (
    .a(\PWM6/n24 ),
    .b(\PWM6/n25_neg_lutinv ),
    .c(dir_pad[6]),
    .d(\PWM6/pnumr [31]),
    .e(pwm_start_stop[22]),
    .o(\PWM6/n32 ));
  AL_MAP_LUT5 #(
    .EQN("(D*~(C)*~((~E*~(B*A)))+D*C*~((~E*~(B*A)))+~(D)*C*(~E*~(B*A))+D*C*(~E*~(B*A)))"),
    .INIT(32'hff00f870))
    _al_u2997 (
    .a(\PWM7/n24 ),
    .b(\PWM7/n25_neg_lutinv ),
    .c(dir_pad[7]),
    .d(\PWM7/pnumr [31]),
    .e(pwm_start_stop[23]),
    .o(\PWM7/n32 ));
  AL_MAP_LUT5 #(
    .EQN("(D*~(C)*~((~E*~(B*A)))+D*C*~((~E*~(B*A)))+~(D)*C*(~E*~(B*A))+D*C*(~E*~(B*A)))"),
    .INIT(32'hff00f870))
    _al_u2998 (
    .a(\PWM8/n24 ),
    .b(\PWM8/n25_neg_lutinv ),
    .c(dir_pad[8]),
    .d(\PWM8/pnumr [31]),
    .e(pwm_start_stop[24]),
    .o(\PWM8/n32 ));
  AL_MAP_LUT5 #(
    .EQN("(D*~(C)*~((~E*~(B*A)))+D*C*~((~E*~(B*A)))+~(D)*C*(~E*~(B*A))+D*C*(~E*~(B*A)))"),
    .INIT(32'hff00f870))
    _al_u2999 (
    .a(\PWM9/n24 ),
    .b(\PWM9/n25_neg_lutinv ),
    .c(dir_pad[9]),
    .d(\PWM9/pnumr [31]),
    .e(pwm_start_stop[25]),
    .o(\PWM9/n32 ));
  EF2_PHY_PAD #(
    //.LOCATION("P114"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u30 (
    .do({open_n901,open_n902,open_n903,dir_pad[8]}),
    .opad(dir[8]));  // CPLD_SOC_AHB_TOP.v(7)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u300 (
    .a(\PWM3/pnumr [23]),
    .b(pnum3[23]),
    .c(pnum3[32]),
    .d(pwm_start_stop[19]),
    .o(\PWM3/n23 [23]));
  AL_MAP_LUT5 #(
    .EQN("(D*~(C)*~((~E*~(B*A)))+D*C*~((~E*~(B*A)))+~(D)*C*(~E*~(B*A))+D*C*(~E*~(B*A)))"),
    .INIT(32'hff00f870))
    _al_u3000 (
    .a(\PWMA/n24 ),
    .b(\PWMA/n25_neg_lutinv ),
    .c(dir_pad[10]),
    .d(\PWMA/pnumr [31]),
    .e(pwm_start_stop[26]),
    .o(\PWMA/n32 ));
  AL_MAP_LUT5 #(
    .EQN("(D*~(C)*~((~E*~(B*A)))+D*C*~((~E*~(B*A)))+~(D)*C*(~E*~(B*A))+D*C*(~E*~(B*A)))"),
    .INIT(32'hff00f870))
    _al_u3001 (
    .a(\PWMB/n24 ),
    .b(\PWMB/n25_neg_lutinv ),
    .c(dir_pad[11]),
    .d(\PWMB/pnumr [31]),
    .e(pwm_start_stop[27]),
    .o(\PWMB/n32 ));
  AL_MAP_LUT5 #(
    .EQN("(D*~(C)*~((~E*~(B*A)))+D*C*~((~E*~(B*A)))+~(D)*C*(~E*~(B*A))+D*C*(~E*~(B*A)))"),
    .INIT(32'hff00f870))
    _al_u3002 (
    .a(\PWMC/n24 ),
    .b(\PWMC/n25_neg_lutinv ),
    .c(dir_pad[12]),
    .d(\PWMC/pnumr [31]),
    .e(pwm_start_stop[28]),
    .o(\PWMC/n32 ));
  AL_MAP_LUT5 #(
    .EQN("(D*~(C)*~((~E*~(B*A)))+D*C*~((~E*~(B*A)))+~(D)*C*(~E*~(B*A))+D*C*(~E*~(B*A)))"),
    .INIT(32'hff00f870))
    _al_u3003 (
    .a(\PWMD/n24 ),
    .b(\PWMD/n25_neg_lutinv ),
    .c(dir_pad[13]),
    .d(\PWMD/pnumr [31]),
    .e(pwm_start_stop[29]),
    .o(\PWMD/n32 ));
  AL_MAP_LUT5 #(
    .EQN("(D*~(C)*~((~E*~(B*A)))+D*C*~((~E*~(B*A)))+~(D)*C*(~E*~(B*A))+D*C*(~E*~(B*A)))"),
    .INIT(32'hff00f870))
    _al_u3004 (
    .a(\PWME/n24 ),
    .b(\PWME/n25_neg_lutinv ),
    .c(dir_pad[14]),
    .d(\PWME/pnumr [31]),
    .e(pwm_start_stop[30]),
    .o(\PWME/n32 ));
  AL_MAP_LUT5 #(
    .EQN("(D*~(C)*~((~E*~(B*A)))+D*C*~((~E*~(B*A)))+~(D)*C*(~E*~(B*A))+D*C*(~E*~(B*A)))"),
    .INIT(32'hff00f870))
    _al_u3005 (
    .a(\PWMF/n24 ),
    .b(\PWMF/n25_neg_lutinv ),
    .c(dir_pad[15]),
    .d(\PWMF/pnumr [31]),
    .e(pwm_start_stop[31]),
    .o(\PWMF/n32 ));
  AL_MAP_LUT4 #(
    .EQN("~(~C*A*~(D*~B))"),
    .INIT(16'hf7f5))
    _al_u3006 (
    .a(_al_u2984_o),
    .b(_al_u1652_o),
    .c(_al_u2988_o),
    .d(ledout_pad[3]),
    .o(n10[3]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(D*C*B*A))"),
    .INIT(32'h00007fff))
    _al_u3007 (
    .a(_al_u1688_o),
    .b(_al_u1690_o),
    .c(_al_u1691_o),
    .d(pnumcnt0[0]),
    .e(\PWM0/stopreq ),
    .o(_al_u3007_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3008 (
    .a(\PWM0/n11 ),
    .b(limit_r_pad[0]),
    .c(limit_l_pad[0]),
    .o(_al_u3008_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*B*~A))"),
    .INIT(16'hf0b0))
    _al_u3009 (
    .a(_al_u3007_o),
    .b(\PWM0/n0_lutinv ),
    .c(_al_u3008_o),
    .d(pwm_start_stop[16]),
    .o(\PWM0/n10 ));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u301 (
    .a(\PWM3/pnumr [22]),
    .b(pnum3[22]),
    .c(pnum3[32]),
    .d(pwm_start_stop[19]),
    .o(\PWM3/n23 [22]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(D*C*B*A))"),
    .INIT(32'h00007fff))
    _al_u3010 (
    .a(_al_u1770_o),
    .b(_al_u1772_o),
    .c(_al_u1773_o),
    .d(pnumcnt1[0]),
    .e(\PWM1/stopreq ),
    .o(_al_u3010_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3011 (
    .a(\PWM1/n11 ),
    .b(limit_r_pad[1]),
    .c(limit_l_pad[1]),
    .o(_al_u3011_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*B*~A))"),
    .INIT(16'hf0b0))
    _al_u3012 (
    .a(_al_u3010_o),
    .b(\PWM1/n0_lutinv ),
    .c(_al_u3011_o),
    .d(pwm_start_stop[17]),
    .o(\PWM1/n10 ));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(D*C*B*A))"),
    .INIT(32'h00007fff))
    _al_u3013 (
    .a(_al_u1852_o),
    .b(_al_u1854_o),
    .c(_al_u1855_o),
    .d(pnumcnt2[0]),
    .e(\PWM2/stopreq ),
    .o(_al_u3013_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3014 (
    .a(\PWM2/n11 ),
    .b(limit_r_pad[2]),
    .c(limit_l_pad[2]),
    .o(_al_u3014_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*B*~A))"),
    .INIT(16'hf0b0))
    _al_u3015 (
    .a(_al_u3013_o),
    .b(\PWM2/n0_lutinv ),
    .c(_al_u3014_o),
    .d(pwm_start_stop[18]),
    .o(\PWM2/n10 ));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(D*C*B*A))"),
    .INIT(32'h00007fff))
    _al_u3016 (
    .a(_al_u1932_o),
    .b(_al_u1934_o),
    .c(_al_u1935_o),
    .d(pnumcnt3[0]),
    .e(\PWM3/stopreq ),
    .o(_al_u3016_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3017 (
    .a(\PWM3/n11 ),
    .b(limit_r_pad[3]),
    .c(limit_l_pad[3]),
    .o(_al_u3017_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*B*~A))"),
    .INIT(16'hf0b0))
    _al_u3018 (
    .a(_al_u3016_o),
    .b(\PWM3/n0_lutinv ),
    .c(_al_u3017_o),
    .d(pwm_start_stop[19]),
    .o(\PWM3/n10 ));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(D*C*B*A))"),
    .INIT(32'h00007fff))
    _al_u3019 (
    .a(_al_u2014_o),
    .b(_al_u2016_o),
    .c(_al_u2017_o),
    .d(pnumcnt4[0]),
    .e(\PWM4/stopreq ),
    .o(_al_u3019_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u302 (
    .a(\PWM3/pnumr [21]),
    .b(pnum3[21]),
    .c(pnum3[32]),
    .d(pwm_start_stop[19]),
    .o(\PWM3/n23 [21]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3020 (
    .a(\PWM4/n11 ),
    .b(limit_r_pad[4]),
    .c(limit_l_pad[4]),
    .o(_al_u3020_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*B*~A))"),
    .INIT(16'hf0b0))
    _al_u3021 (
    .a(_al_u3019_o),
    .b(\PWM4/n0_lutinv ),
    .c(_al_u3020_o),
    .d(pwm_start_stop[20]),
    .o(\PWM4/n10 ));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(D*C*B*A))"),
    .INIT(32'h00007fff))
    _al_u3022 (
    .a(_al_u2096_o),
    .b(_al_u2098_o),
    .c(_al_u2099_o),
    .d(pnumcnt5[0]),
    .e(\PWM5/stopreq ),
    .o(_al_u3022_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3023 (
    .a(\PWM5/n11 ),
    .b(limit_r_pad[5]),
    .c(limit_l_pad[5]),
    .o(_al_u3023_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*B*~A))"),
    .INIT(16'hf0b0))
    _al_u3024 (
    .a(_al_u3022_o),
    .b(\PWM5/n0_lutinv ),
    .c(_al_u3023_o),
    .d(pwm_start_stop[21]),
    .o(\PWM5/n10 ));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(D*C*B*A))"),
    .INIT(32'h00007fff))
    _al_u3025 (
    .a(_al_u2178_o),
    .b(_al_u2180_o),
    .c(_al_u2181_o),
    .d(pnumcnt6[0]),
    .e(\PWM6/stopreq ),
    .o(_al_u3025_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3026 (
    .a(\PWM6/n11 ),
    .b(limit_l_pad[6]),
    .c(limit_r_pad[6]),
    .o(_al_u3026_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*B*~A))"),
    .INIT(16'hf0b0))
    _al_u3027 (
    .a(_al_u3025_o),
    .b(\PWM6/n0_lutinv ),
    .c(_al_u3026_o),
    .d(pwm_start_stop[22]),
    .o(\PWM6/n10 ));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(D*C*B*A))"),
    .INIT(32'h00007fff))
    _al_u3028 (
    .a(_al_u2258_o),
    .b(_al_u2260_o),
    .c(_al_u2261_o),
    .d(pnumcnt7[0]),
    .e(\PWM7/stopreq ),
    .o(_al_u3028_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3029 (
    .a(\PWM7/n11 ),
    .b(limit_l_pad[7]),
    .c(limit_r_pad[7]),
    .o(_al_u3029_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u303 (
    .a(\PWM3/pnumr [20]),
    .b(pnum3[20]),
    .c(pnum3[32]),
    .d(pwm_start_stop[19]),
    .o(\PWM3/n23 [20]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*B*~A))"),
    .INIT(16'hf0b0))
    _al_u3030 (
    .a(_al_u3028_o),
    .b(\PWM7/n0_lutinv ),
    .c(_al_u3029_o),
    .d(pwm_start_stop[23]),
    .o(\PWM7/n10 ));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(D*C*B*A))"),
    .INIT(32'h00007fff))
    _al_u3031 (
    .a(_al_u2340_o),
    .b(_al_u2342_o),
    .c(_al_u2343_o),
    .d(pnumcnt8[0]),
    .e(\PWM8/stopreq ),
    .o(_al_u3031_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3032 (
    .a(\PWM8/n11 ),
    .b(limit_l_pad[8]),
    .c(limit_r_pad[8]),
    .o(_al_u3032_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*B*~A))"),
    .INIT(16'hf0b0))
    _al_u3033 (
    .a(_al_u3031_o),
    .b(\PWM8/n0_lutinv ),
    .c(_al_u3032_o),
    .d(pwm_start_stop[24]),
    .o(\PWM8/n10 ));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(D*C*B*A))"),
    .INIT(32'h00007fff))
    _al_u3034 (
    .a(_al_u2420_o),
    .b(_al_u2422_o),
    .c(_al_u2423_o),
    .d(pnumcnt9[0]),
    .e(\PWM9/stopreq ),
    .o(_al_u3034_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3035 (
    .a(\PWM9/n11 ),
    .b(limit_l_pad[9]),
    .c(limit_r_pad[9]),
    .o(_al_u3035_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*B*~A))"),
    .INIT(16'hf0b0))
    _al_u3036 (
    .a(_al_u3034_o),
    .b(\PWM9/n0_lutinv ),
    .c(_al_u3035_o),
    .d(pwm_start_stop[25]),
    .o(\PWM9/n10 ));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(D*C*B*A))"),
    .INIT(32'h00007fff))
    _al_u3037 (
    .a(_al_u2502_o),
    .b(_al_u2504_o),
    .c(_al_u2505_o),
    .d(pnumcntA[0]),
    .e(\PWMA/stopreq ),
    .o(_al_u3037_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3038 (
    .a(\PWMA/n11 ),
    .b(limit_l_pad[10]),
    .c(limit_r_pad[10]),
    .o(_al_u3038_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*B*~A))"),
    .INIT(16'hf0b0))
    _al_u3039 (
    .a(_al_u3037_o),
    .b(\PWMA/n0_lutinv ),
    .c(_al_u3038_o),
    .d(pwm_start_stop[26]),
    .o(\PWMA/n10 ));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u304 (
    .a(\PWM3/pnumr [2]),
    .b(pnum3[2]),
    .c(pnum3[32]),
    .d(pwm_start_stop[19]),
    .o(\PWM3/n23 [2]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(D*C*B*A))"),
    .INIT(32'h00007fff))
    _al_u3040 (
    .a(_al_u2581_o),
    .b(_al_u2583_o),
    .c(_al_u2584_o),
    .d(pnumcntB[0]),
    .e(\PWMB/stopreq ),
    .o(_al_u3040_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3041 (
    .a(\PWMB/n11 ),
    .b(limit_l_pad[11]),
    .c(limit_r_pad[11]),
    .o(_al_u3041_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*B*~A))"),
    .INIT(16'hf0b0))
    _al_u3042 (
    .a(_al_u3040_o),
    .b(\PWMB/n0_lutinv ),
    .c(_al_u3041_o),
    .d(pwm_start_stop[27]),
    .o(\PWMB/n10 ));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(D*C*B*A))"),
    .INIT(32'h00007fff))
    _al_u3043 (
    .a(_al_u2663_o),
    .b(_al_u2665_o),
    .c(_al_u2666_o),
    .d(pnumcntC[0]),
    .e(\PWMC/stopreq ),
    .o(_al_u3043_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3044 (
    .a(\PWMC/n11 ),
    .b(limit_l_pad[12]),
    .c(limit_r_pad[12]),
    .o(_al_u3044_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*B*~A))"),
    .INIT(16'hf0b0))
    _al_u3045 (
    .a(_al_u3043_o),
    .b(\PWMC/n0_lutinv ),
    .c(_al_u3044_o),
    .d(pwm_start_stop[28]),
    .o(\PWMC/n10 ));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(D*C*B*A))"),
    .INIT(32'h00007fff))
    _al_u3046 (
    .a(_al_u2742_o),
    .b(_al_u2744_o),
    .c(_al_u2745_o),
    .d(pnumcntD[0]),
    .e(\PWMD/stopreq ),
    .o(_al_u3046_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3047 (
    .a(\PWMD/n11 ),
    .b(limit_l_pad[13]),
    .c(limit_r_pad[13]),
    .o(_al_u3047_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*B*~A))"),
    .INIT(16'hf0b0))
    _al_u3048 (
    .a(_al_u3046_o),
    .b(\PWMD/n0_lutinv ),
    .c(_al_u3047_o),
    .d(pwm_start_stop[29]),
    .o(\PWMD/n10 ));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(D*C*B*A))"),
    .INIT(32'h00007fff))
    _al_u3049 (
    .a(_al_u2822_o),
    .b(_al_u2824_o),
    .c(_al_u2825_o),
    .d(pnumcntE[0]),
    .e(\PWME/stopreq ),
    .o(_al_u3049_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u305 (
    .a(\PWM3/pnumr [19]),
    .b(pnum3[19]),
    .c(pnum3[32]),
    .d(pwm_start_stop[19]),
    .o(\PWM3/n23 [19]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3050 (
    .a(\PWME/n11 ),
    .b(limit_l_pad[14]),
    .c(limit_r_pad[14]),
    .o(_al_u3050_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*B*~A))"),
    .INIT(16'hf0b0))
    _al_u3051 (
    .a(_al_u3049_o),
    .b(\PWME/n0_lutinv ),
    .c(_al_u3050_o),
    .d(pwm_start_stop[30]),
    .o(\PWME/n10 ));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(D*C*B*A))"),
    .INIT(32'h00007fff))
    _al_u3052 (
    .a(_al_u2901_o),
    .b(_al_u2903_o),
    .c(_al_u2904_o),
    .d(pnumcntF[0]),
    .e(\PWMF/stopreq ),
    .o(_al_u3052_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u3053 (
    .a(\PWMF/n11 ),
    .b(limit_l_pad[15]),
    .c(limit_r_pad[15]),
    .o(_al_u3053_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*B*~A))"),
    .INIT(16'hf0b0))
    _al_u3054 (
    .a(_al_u3052_o),
    .b(\PWMF/n0_lutinv ),
    .c(_al_u3053_o),
    .d(pwm_start_stop[31]),
    .o(\PWMF/n10 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3055 (
    .a(_al_u1652_o),
    .b(_al_u2988_o),
    .o(_al_u3055_o));
  AL_MAP_LUT2 #(
    .EQN("~(B*A)"),
    .INIT(4'h7))
    _al_u3056 (
    .a(_al_u2984_o),
    .b(_al_u3055_o),
    .o(_al_n1_en));
  AL_MAP_LUT4 #(
    .EQN("~(C*~(~B*~(~D*A)))"),
    .INIT(16'h3f1f))
    _al_u3057 (
    .a(_al_u3055_o),
    .b(_al_u2983_o),
    .c(n4_neg),
    .d(ledout_pad[1]),
    .o(n10[1]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*~A)"),
    .INIT(32'h00000001))
    _al_u3058 (
    .a(\U_AHB/h2h_haddr [2]),
    .b(\U_AHB/h2h_haddr [3]),
    .c(\U_AHB/h2h_haddr [4]),
    .d(\U_AHB/h2h_haddr [5]),
    .e(\U_AHB/h2h_haddr [6]),
    .o(\U_AHB/n95_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3059 (
    .a(\U_AHB/n95_lutinv ),
    .b(\U_AHB/h2h_haddr [7]),
    .o(\U_AHB/n96 ));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u306 (
    .a(\PWM3/pnumr [18]),
    .b(pnum3[18]),
    .c(pnum3[32]),
    .d(pwm_start_stop[19]),
    .o(\PWM3/n23 [18]));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    _al_u3060 (
    .a(\U_AHB/n95_lutinv ),
    .b(\U_AHB/h2h_haddr [7]),
    .c(\U_AHB/h2h_haddr [8]),
    .d(\U_AHB/h2h_haddr [9]),
    .o(\U_AHB/n102 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u3061 (
    .a(\U_AHB/h2h_hwrite ),
    .b(\U_AHB/h2h_haddr [14]),
    .o(_al_u3061_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~(E*B)*~(D*A)))"),
    .INIT(32'he0c0a000))
    _al_u3062 (
    .a(\U_AHB/n96 ),
    .b(\U_AHB/n102 ),
    .c(_al_u3061_o),
    .d(pwm_state_read[15]),
    .e(limit_l_pad[15]),
    .o(_al_u3062_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u3063 (
    .a(\U_AHB/n95_lutinv ),
    .b(\U_AHB/h2h_haddr [7]),
    .c(\U_AHB/h2h_haddr [8]),
    .d(\U_AHB/h2h_haddr [9]),
    .o(\U_AHB/n104_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u3064 (
    .a(\U_AHB/n104_lutinv ),
    .b(\U_AHB/h2h_haddr [12]),
    .c(\U_AHB/h2h_haddr [10]),
    .d(\U_AHB/h2h_haddr [11]),
    .o(\U_AHB/n113_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u3065 (
    .a(\U_AHB/n104_lutinv ),
    .b(_al_u3061_o),
    .o(_al_u3065_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u3066 (
    .a(\U_AHB/h2h_hwrite ),
    .b(\U_AHB/h2h_haddr [13]),
    .c(\U_AHB/h2h_haddr [14]),
    .o(\U_AHB/n82 ));
  AL_MAP_LUT5 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8caf00aa))
    _al_u3067 (
    .a(_al_u3062_o),
    .b(\U_AHB/n113_lutinv ),
    .c(_al_u3065_o),
    .d(\U_AHB/n82 ),
    .e(\U_AHB/h2h_hrdata [31]),
    .o(\U_AHB/n118 [31]));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~(E*B)*~(D*A)))"),
    .INIT(32'he0c0a000))
    _al_u3068 (
    .a(\U_AHB/n96 ),
    .b(\U_AHB/n102 ),
    .c(_al_u3061_o),
    .d(pwm_state_read[14]),
    .e(limit_l_pad[14]),
    .o(_al_u3068_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8caf00aa))
    _al_u3069 (
    .a(_al_u3068_o),
    .b(\U_AHB/n113_lutinv ),
    .c(_al_u3065_o),
    .d(\U_AHB/n82 ),
    .e(\U_AHB/h2h_hrdata [30]),
    .o(\U_AHB/n118 [30]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u307 (
    .a(\PWM3/pnumr [17]),
    .b(pnum3[17]),
    .c(pnum3[32]),
    .d(pwm_start_stop[19]),
    .o(\PWM3/n23 [17]));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~(E*B)*~(D*A)))"),
    .INIT(32'he0c0a000))
    _al_u3070 (
    .a(\U_AHB/n96 ),
    .b(\U_AHB/n102 ),
    .c(_al_u3061_o),
    .d(pwm_state_read[13]),
    .e(limit_l_pad[13]),
    .o(_al_u3070_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8caf00aa))
    _al_u3071 (
    .a(_al_u3070_o),
    .b(\U_AHB/n113_lutinv ),
    .c(_al_u3065_o),
    .d(\U_AHB/n82 ),
    .e(\U_AHB/h2h_hrdata [29]),
    .o(\U_AHB/n118 [29]));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~(E*B)*~(D*A)))"),
    .INIT(32'he0c0a000))
    _al_u3072 (
    .a(\U_AHB/n96 ),
    .b(\U_AHB/n102 ),
    .c(_al_u3061_o),
    .d(pwm_state_read[12]),
    .e(limit_l_pad[12]),
    .o(_al_u3072_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8caf00aa))
    _al_u3073 (
    .a(_al_u3072_o),
    .b(\U_AHB/n113_lutinv ),
    .c(_al_u3065_o),
    .d(\U_AHB/n82 ),
    .e(\U_AHB/h2h_hrdata [28]),
    .o(\U_AHB/n118 [28]));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~(E*B)*~(D*A)))"),
    .INIT(32'he0c0a000))
    _al_u3074 (
    .a(\U_AHB/n96 ),
    .b(\U_AHB/n102 ),
    .c(_al_u3061_o),
    .d(pwm_state_read[11]),
    .e(limit_l_pad[11]),
    .o(_al_u3074_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8caf00aa))
    _al_u3075 (
    .a(_al_u3074_o),
    .b(\U_AHB/n113_lutinv ),
    .c(_al_u3065_o),
    .d(\U_AHB/n82 ),
    .e(\U_AHB/h2h_hrdata [27]),
    .o(\U_AHB/n118 [27]));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~(E*B)*~(D*A)))"),
    .INIT(32'he0c0a000))
    _al_u3076 (
    .a(\U_AHB/n96 ),
    .b(\U_AHB/n102 ),
    .c(_al_u3061_o),
    .d(pwm_state_read[10]),
    .e(limit_l_pad[10]),
    .o(_al_u3076_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8caf00aa))
    _al_u3077 (
    .a(_al_u3076_o),
    .b(\U_AHB/n113_lutinv ),
    .c(_al_u3065_o),
    .d(\U_AHB/n82 ),
    .e(\U_AHB/h2h_hrdata [26]),
    .o(\U_AHB/n118 [26]));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~(E*B)*~(D*A)))"),
    .INIT(32'he0c0a000))
    _al_u3078 (
    .a(\U_AHB/n96 ),
    .b(\U_AHB/n102 ),
    .c(_al_u3061_o),
    .d(pwm_state_read[9]),
    .e(limit_l_pad[9]),
    .o(_al_u3078_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8caf00aa))
    _al_u3079 (
    .a(_al_u3078_o),
    .b(\U_AHB/n113_lutinv ),
    .c(_al_u3065_o),
    .d(\U_AHB/n82 ),
    .e(\U_AHB/h2h_hrdata [25]),
    .o(\U_AHB/n118 [25]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u308 (
    .a(\PWM3/pnumr [16]),
    .b(pnum3[16]),
    .c(pnum3[32]),
    .d(pwm_start_stop[19]),
    .o(\PWM3/n23 [16]));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~(E*B)*~(D*A)))"),
    .INIT(32'he0c0a000))
    _al_u3080 (
    .a(\U_AHB/n96 ),
    .b(\U_AHB/n102 ),
    .c(_al_u3061_o),
    .d(pwm_state_read[8]),
    .e(limit_l_pad[8]),
    .o(_al_u3080_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8caf00aa))
    _al_u3081 (
    .a(_al_u3080_o),
    .b(\U_AHB/n113_lutinv ),
    .c(_al_u3065_o),
    .d(\U_AHB/n82 ),
    .e(\U_AHB/h2h_hrdata [24]),
    .o(\U_AHB/n118 [24]));
  AL_MAP_LUT4 #(
    .EQN("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    .INIT(16'h535f))
    _al_u3082 (
    .a(pnumcnt0[9]),
    .b(pnumcnt1[9]),
    .c(\U_AHB/h2h_haddr [2]),
    .d(\U_AHB/h2h_haddr [3]),
    .o(_al_u3082_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    _al_u3083 (
    .a(\U_AHB/h2h_haddr [2]),
    .b(\U_AHB/h2h_haddr [3]),
    .c(\U_AHB/h2h_haddr [4]),
    .d(\U_AHB/h2h_haddr [5]),
    .o(\U_AHB/n90 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u3084 (
    .a(\U_AHB/h2h_haddr [2]),
    .b(\U_AHB/h2h_haddr [3]),
    .c(\U_AHB/h2h_haddr [4]),
    .o(\U_AHB/n87 ));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3085 (
    .a(_al_u3082_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcnt2[9]),
    .e(pnumcnt3[9]),
    .o(_al_u3085_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*~B*~A)"),
    .INIT(32'h00010000))
    _al_u3086 (
    .a(\U_AHB/h2h_haddr [2]),
    .b(\U_AHB/h2h_haddr [3]),
    .c(\U_AHB/h2h_haddr [4]),
    .d(\U_AHB/h2h_haddr [5]),
    .e(\U_AHB/h2h_haddr [6]),
    .o(\U_AHB/n93 ));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3087 (
    .a(_al_u3085_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcnt4[9]),
    .e(pnumcnt5[9]),
    .o(_al_u3087_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u3088 (
    .a(\U_AHB/n95_lutinv ),
    .b(\U_AHB/h2h_haddr [7]),
    .c(\U_AHB/h2h_haddr [8]),
    .o(\U_AHB/n99 ));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3089 (
    .a(_al_u3087_o),
    .b(\U_AHB/n102 ),
    .c(\U_AHB/n99 ),
    .d(pnumcnt6[9]),
    .e(pnumcnt7[9]),
    .o(_al_u3089_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u309 (
    .a(\PWM3/pnumr [15]),
    .b(pnum3[15]),
    .c(pnum3[32]),
    .d(pwm_start_stop[19]),
    .o(\PWM3/n23 [15]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u3090 (
    .a(\U_AHB/n104_lutinv ),
    .b(\U_AHB/h2h_haddr [10]),
    .c(\U_AHB/h2h_haddr [11]),
    .o(\U_AHB/n108 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u3091 (
    .a(\U_AHB/n104_lutinv ),
    .b(\U_AHB/h2h_haddr [10]),
    .o(\U_AHB/n105 ));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3092 (
    .a(_al_u3089_o),
    .b(\U_AHB/n108 ),
    .c(\U_AHB/n105 ),
    .d(pnumcnt8[9]),
    .e(pnumcnt9[9]),
    .o(_al_u3092_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u3093 (
    .a(\U_AHB/n104_lutinv ),
    .b(\U_AHB/h2h_haddr [12]),
    .c(\U_AHB/h2h_haddr [10]),
    .d(\U_AHB/h2h_haddr [11]),
    .o(\U_AHB/n111 ));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3094 (
    .a(_al_u3092_o),
    .b(\U_AHB/n113_lutinv ),
    .c(\U_AHB/n111 ),
    .d(pnumcntA[9]),
    .e(\U_AHB/h2h_hrdata [9]),
    .o(_al_u3094_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((E*C)*~(B)*~(D)+(E*C)*B*~(D)+~((E*C))*B*D+(E*C)*B*D))"),
    .INIT(32'h220a22aa))
    _al_u3095 (
    .a(_al_u3061_o),
    .b(pnumcntB[9]),
    .c(pnumcntC[9]),
    .d(\U_AHB/h2h_haddr [2]),
    .e(\U_AHB/h2h_haddr [3]),
    .o(_al_u3095_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3096 (
    .a(_al_u3095_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcntD[9]),
    .e(pnumcntE[9]),
    .o(_al_u3096_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3097 (
    .a(_al_u3096_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcntF[9]),
    .e(pwm_state_read[9]),
    .o(_al_u3097_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*C)*~(D*B))"),
    .INIT(32'h020a22aa))
    _al_u3098 (
    .a(_al_u3097_o),
    .b(\U_AHB/n104_lutinv ),
    .c(\U_AHB/n102 ),
    .d(\U_AHB/h2h_hrdata [9]),
    .e(limit_r_pad[9]),
    .o(_al_u3098_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h33533050))
    _al_u3099 (
    .a(_al_u3094_o),
    .b(_al_u3098_o),
    .c(_al_u3061_o),
    .d(\U_AHB/h2h_haddr [13]),
    .e(\U_AHB/h2h_hrdata [9]),
    .o(\U_AHB/n118 [9]));
  EF2_PHY_PAD #(
    //.LOCATION("P122"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u31 (
    .do({open_n924,open_n925,open_n926,dir_pad[7]}),
    .opad(dir[7]));  // CPLD_SOC_AHB_TOP.v(7)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u310 (
    .a(\PWM3/pnumr [14]),
    .b(pnum3[14]),
    .c(pnum3[32]),
    .d(pwm_start_stop[19]),
    .o(\PWM3/n23 [14]));
  AL_MAP_LUT4 #(
    .EQN("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    .INIT(16'h535f))
    _al_u3100 (
    .a(pnumcnt0[8]),
    .b(pnumcnt1[8]),
    .c(\U_AHB/h2h_haddr [2]),
    .d(\U_AHB/h2h_haddr [3]),
    .o(_al_u3100_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3101 (
    .a(_al_u3100_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcnt2[8]),
    .e(pnumcnt3[8]),
    .o(_al_u3101_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3102 (
    .a(_al_u3101_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcnt4[8]),
    .e(pnumcnt5[8]),
    .o(_al_u3102_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3103 (
    .a(_al_u3102_o),
    .b(\U_AHB/n102 ),
    .c(\U_AHB/n99 ),
    .d(pnumcnt6[8]),
    .e(pnumcnt7[8]),
    .o(_al_u3103_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3104 (
    .a(_al_u3103_o),
    .b(\U_AHB/n108 ),
    .c(\U_AHB/n105 ),
    .d(pnumcnt8[8]),
    .e(pnumcnt9[8]),
    .o(_al_u3104_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3105 (
    .a(_al_u3104_o),
    .b(\U_AHB/n113_lutinv ),
    .c(\U_AHB/n111 ),
    .d(pnumcntA[8]),
    .e(\U_AHB/h2h_hrdata [8]),
    .o(_al_u3105_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((E*C)*~(B)*~(D)+(E*C)*B*~(D)+~((E*C))*B*D+(E*C)*B*D))"),
    .INIT(32'h220a22aa))
    _al_u3106 (
    .a(_al_u3061_o),
    .b(pnumcntB[8]),
    .c(pnumcntC[8]),
    .d(\U_AHB/h2h_haddr [2]),
    .e(\U_AHB/h2h_haddr [3]),
    .o(_al_u3106_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3107 (
    .a(_al_u3106_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcntD[8]),
    .e(pnumcntE[8]),
    .o(_al_u3107_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3108 (
    .a(_al_u3107_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcntF[8]),
    .e(pwm_state_read[8]),
    .o(_al_u3108_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*C)*~(D*B))"),
    .INIT(32'h020a22aa))
    _al_u3109 (
    .a(_al_u3108_o),
    .b(\U_AHB/n104_lutinv ),
    .c(\U_AHB/n102 ),
    .d(\U_AHB/h2h_hrdata [8]),
    .e(limit_r_pad[8]),
    .o(_al_u3109_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u311 (
    .a(\PWM3/pnumr [13]),
    .b(pnum3[13]),
    .c(pnum3[32]),
    .d(pwm_start_stop[19]),
    .o(\PWM3/n23 [13]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h33533050))
    _al_u3110 (
    .a(_al_u3105_o),
    .b(_al_u3109_o),
    .c(_al_u3061_o),
    .d(\U_AHB/h2h_haddr [13]),
    .e(\U_AHB/h2h_hrdata [8]),
    .o(\U_AHB/n118 [8]));
  AL_MAP_LUT4 #(
    .EQN("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    .INIT(16'h535f))
    _al_u3111 (
    .a(pnumcnt0[7]),
    .b(pnumcnt1[7]),
    .c(\U_AHB/h2h_haddr [2]),
    .d(\U_AHB/h2h_haddr [3]),
    .o(_al_u3111_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3112 (
    .a(_al_u3111_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcnt2[7]),
    .e(pnumcnt3[7]),
    .o(_al_u3112_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3113 (
    .a(_al_u3112_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcnt4[7]),
    .e(pnumcnt5[7]),
    .o(_al_u3113_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3114 (
    .a(_al_u3113_o),
    .b(\U_AHB/n102 ),
    .c(\U_AHB/n99 ),
    .d(pnumcnt6[7]),
    .e(pnumcnt7[7]),
    .o(_al_u3114_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3115 (
    .a(_al_u3114_o),
    .b(\U_AHB/n108 ),
    .c(\U_AHB/n105 ),
    .d(pnumcnt8[7]),
    .e(pnumcnt9[7]),
    .o(_al_u3115_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3116 (
    .a(_al_u3115_o),
    .b(\U_AHB/n113_lutinv ),
    .c(\U_AHB/n111 ),
    .d(pnumcntA[7]),
    .e(\U_AHB/h2h_hrdata [7]),
    .o(_al_u3116_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((E*C)*~(B)*~(D)+(E*C)*B*~(D)+~((E*C))*B*D+(E*C)*B*D))"),
    .INIT(32'h220a22aa))
    _al_u3117 (
    .a(_al_u3061_o),
    .b(pnumcntB[7]),
    .c(pnumcntC[7]),
    .d(\U_AHB/h2h_haddr [2]),
    .e(\U_AHB/h2h_haddr [3]),
    .o(_al_u3117_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3118 (
    .a(_al_u3117_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcntD[7]),
    .e(pnumcntE[7]),
    .o(_al_u3118_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3119 (
    .a(_al_u3118_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcntF[7]),
    .e(pwm_state_read[7]),
    .o(_al_u3119_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u312 (
    .a(\PWM3/pnumr [12]),
    .b(pnum3[12]),
    .c(pnum3[32]),
    .d(pwm_start_stop[19]),
    .o(\PWM3/n23 [12]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*C)*~(D*B))"),
    .INIT(32'h020a22aa))
    _al_u3120 (
    .a(_al_u3119_o),
    .b(\U_AHB/n104_lutinv ),
    .c(\U_AHB/n102 ),
    .d(\U_AHB/h2h_hrdata [7]),
    .e(limit_r_pad[7]),
    .o(_al_u3120_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h33533050))
    _al_u3121 (
    .a(_al_u3116_o),
    .b(_al_u3120_o),
    .c(_al_u3061_o),
    .d(\U_AHB/h2h_haddr [13]),
    .e(\U_AHB/h2h_hrdata [7]),
    .o(\U_AHB/n118 [7]));
  AL_MAP_LUT4 #(
    .EQN("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    .INIT(16'h535f))
    _al_u3122 (
    .a(pnumcnt0[6]),
    .b(pnumcnt1[6]),
    .c(\U_AHB/h2h_haddr [2]),
    .d(\U_AHB/h2h_haddr [3]),
    .o(_al_u3122_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3123 (
    .a(_al_u3122_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcnt2[6]),
    .e(pnumcnt3[6]),
    .o(_al_u3123_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3124 (
    .a(_al_u3123_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcnt4[6]),
    .e(pnumcnt5[6]),
    .o(_al_u3124_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3125 (
    .a(_al_u3124_o),
    .b(\U_AHB/n102 ),
    .c(\U_AHB/n99 ),
    .d(pnumcnt6[6]),
    .e(pnumcnt7[6]),
    .o(_al_u3125_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3126 (
    .a(_al_u3125_o),
    .b(\U_AHB/n108 ),
    .c(\U_AHB/n105 ),
    .d(pnumcnt8[6]),
    .e(pnumcnt9[6]),
    .o(_al_u3126_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3127 (
    .a(_al_u3126_o),
    .b(\U_AHB/n113_lutinv ),
    .c(\U_AHB/n111 ),
    .d(pnumcntA[6]),
    .e(\U_AHB/h2h_hrdata [6]),
    .o(_al_u3127_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((E*C)*~(B)*~(D)+(E*C)*B*~(D)+~((E*C))*B*D+(E*C)*B*D))"),
    .INIT(32'h220a22aa))
    _al_u3128 (
    .a(_al_u3061_o),
    .b(pnumcntB[6]),
    .c(pnumcntC[6]),
    .d(\U_AHB/h2h_haddr [2]),
    .e(\U_AHB/h2h_haddr [3]),
    .o(_al_u3128_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3129 (
    .a(_al_u3128_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcntD[6]),
    .e(pnumcntE[6]),
    .o(_al_u3129_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u313 (
    .a(\PWM3/pnumr [11]),
    .b(pnum3[11]),
    .c(pnum3[32]),
    .d(pwm_start_stop[19]),
    .o(\PWM3/n23 [11]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3130 (
    .a(_al_u3129_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcntF[6]),
    .e(pwm_state_read[6]),
    .o(_al_u3130_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*C)*~(D*B))"),
    .INIT(32'h020a22aa))
    _al_u3131 (
    .a(_al_u3130_o),
    .b(\U_AHB/n104_lutinv ),
    .c(\U_AHB/n102 ),
    .d(\U_AHB/h2h_hrdata [6]),
    .e(limit_r_pad[6]),
    .o(_al_u3131_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h33533050))
    _al_u3132 (
    .a(_al_u3127_o),
    .b(_al_u3131_o),
    .c(_al_u3061_o),
    .d(\U_AHB/h2h_haddr [13]),
    .e(\U_AHB/h2h_hrdata [6]),
    .o(\U_AHB/n118 [6]));
  AL_MAP_LUT4 #(
    .EQN("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    .INIT(16'h535f))
    _al_u3133 (
    .a(pnumcnt0[5]),
    .b(pnumcnt1[5]),
    .c(\U_AHB/h2h_haddr [2]),
    .d(\U_AHB/h2h_haddr [3]),
    .o(_al_u3133_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3134 (
    .a(_al_u3133_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcnt2[5]),
    .e(pnumcnt3[5]),
    .o(_al_u3134_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3135 (
    .a(_al_u3134_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcnt4[5]),
    .e(pnumcnt5[5]),
    .o(_al_u3135_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3136 (
    .a(_al_u3135_o),
    .b(\U_AHB/n102 ),
    .c(\U_AHB/n99 ),
    .d(pnumcnt6[5]),
    .e(pnumcnt7[5]),
    .o(_al_u3136_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3137 (
    .a(_al_u3136_o),
    .b(\U_AHB/n108 ),
    .c(\U_AHB/n105 ),
    .d(pnumcnt8[5]),
    .e(pnumcnt9[5]),
    .o(_al_u3137_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3138 (
    .a(_al_u3137_o),
    .b(\U_AHB/n113_lutinv ),
    .c(\U_AHB/n111 ),
    .d(pnumcntA[5]),
    .e(\U_AHB/h2h_hrdata [5]),
    .o(_al_u3138_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u3139 (
    .a(\U_AHB/n96 ),
    .b(_al_u3061_o),
    .c(pwm_state_read[5]),
    .o(_al_u3139_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u314 (
    .a(\PWM3/pnumr [10]),
    .b(pnum3[10]),
    .c(pnum3[32]),
    .d(pwm_start_stop[19]),
    .o(\PWM3/n23 [10]));
  AL_MAP_LUT4 #(
    .EQN("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    .INIT(16'h535f))
    _al_u3140 (
    .a(pnumcntB[5]),
    .b(pnumcntC[5]),
    .c(\U_AHB/h2h_haddr [2]),
    .d(\U_AHB/h2h_haddr [3]),
    .o(_al_u3140_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3141 (
    .a(_al_u3140_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcntD[5]),
    .e(pnumcntE[5]),
    .o(_al_u3141_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u3142 (
    .a(_al_u3139_o),
    .b(_al_u3141_o),
    .c(\U_AHB/n93 ),
    .d(pnumcntF[5]),
    .o(_al_u3142_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*C)*~(D*B))"),
    .INIT(32'h020a22aa))
    _al_u3143 (
    .a(_al_u3142_o),
    .b(\U_AHB/n104_lutinv ),
    .c(\U_AHB/n102 ),
    .d(\U_AHB/h2h_hrdata [5]),
    .e(limit_r_pad[5]),
    .o(_al_u3143_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h33533050))
    _al_u3144 (
    .a(_al_u3138_o),
    .b(_al_u3143_o),
    .c(_al_u3061_o),
    .d(\U_AHB/h2h_haddr [13]),
    .e(\U_AHB/h2h_hrdata [5]),
    .o(\U_AHB/n118 [5]));
  AL_MAP_LUT4 #(
    .EQN("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    .INIT(16'h535f))
    _al_u3145 (
    .a(pnumcnt0[4]),
    .b(pnumcnt1[4]),
    .c(\U_AHB/h2h_haddr [2]),
    .d(\U_AHB/h2h_haddr [3]),
    .o(_al_u3145_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3146 (
    .a(_al_u3145_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcnt2[4]),
    .e(pnumcnt3[4]),
    .o(_al_u3146_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3147 (
    .a(_al_u3146_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcnt4[4]),
    .e(pnumcnt5[4]),
    .o(_al_u3147_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3148 (
    .a(_al_u3147_o),
    .b(\U_AHB/n102 ),
    .c(\U_AHB/n99 ),
    .d(pnumcnt6[4]),
    .e(pnumcnt7[4]),
    .o(_al_u3148_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3149 (
    .a(_al_u3148_o),
    .b(\U_AHB/n108 ),
    .c(\U_AHB/n105 ),
    .d(pnumcnt8[4]),
    .e(pnumcnt9[4]),
    .o(_al_u3149_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u315 (
    .a(\PWM3/pnumr [1]),
    .b(pnum3[1]),
    .c(pnum3[32]),
    .d(pwm_start_stop[19]),
    .o(\PWM3/n23 [1]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3150 (
    .a(_al_u3149_o),
    .b(\U_AHB/n113_lutinv ),
    .c(\U_AHB/n111 ),
    .d(pnumcntA[4]),
    .e(\U_AHB/h2h_hrdata [4]),
    .o(_al_u3150_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((E*C)*~(B)*~(D)+(E*C)*B*~(D)+~((E*C))*B*D+(E*C)*B*D))"),
    .INIT(32'h220a22aa))
    _al_u3151 (
    .a(_al_u3061_o),
    .b(pnumcntB[4]),
    .c(pnumcntC[4]),
    .d(\U_AHB/h2h_haddr [2]),
    .e(\U_AHB/h2h_haddr [3]),
    .o(_al_u3151_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3152 (
    .a(_al_u3151_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcntD[4]),
    .e(pnumcntE[4]),
    .o(_al_u3152_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3153 (
    .a(_al_u3152_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcntF[4]),
    .e(pwm_state_read[4]),
    .o(_al_u3153_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*C)*~(D*B))"),
    .INIT(32'h020a22aa))
    _al_u3154 (
    .a(_al_u3153_o),
    .b(\U_AHB/n104_lutinv ),
    .c(\U_AHB/n102 ),
    .d(\U_AHB/h2h_hrdata [4]),
    .e(limit_r_pad[4]),
    .o(_al_u3154_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h33533050))
    _al_u3155 (
    .a(_al_u3150_o),
    .b(_al_u3154_o),
    .c(_al_u3061_o),
    .d(\U_AHB/h2h_haddr [13]),
    .e(\U_AHB/h2h_hrdata [4]),
    .o(\U_AHB/n118 [4]));
  AL_MAP_LUT4 #(
    .EQN("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    .INIT(16'h535f))
    _al_u3156 (
    .a(pnumcnt0[3]),
    .b(pnumcnt1[3]),
    .c(\U_AHB/h2h_haddr [2]),
    .d(\U_AHB/h2h_haddr [3]),
    .o(_al_u3156_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3157 (
    .a(_al_u3156_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcnt2[3]),
    .e(pnumcnt3[3]),
    .o(_al_u3157_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3158 (
    .a(_al_u3157_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcnt4[3]),
    .e(pnumcnt5[3]),
    .o(_al_u3158_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3159 (
    .a(_al_u3158_o),
    .b(\U_AHB/n102 ),
    .c(\U_AHB/n99 ),
    .d(pnumcnt6[3]),
    .e(pnumcnt7[3]),
    .o(_al_u3159_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u316 (
    .a(\PWM3/pnumr [0]),
    .b(pnum3[0]),
    .c(pnum3[32]),
    .d(pwm_start_stop[19]),
    .o(\PWM3/n23 [0]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3160 (
    .a(_al_u3159_o),
    .b(\U_AHB/n108 ),
    .c(\U_AHB/n105 ),
    .d(pnumcnt8[3]),
    .e(pnumcnt9[3]),
    .o(_al_u3160_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3161 (
    .a(_al_u3160_o),
    .b(\U_AHB/n113_lutinv ),
    .c(\U_AHB/n111 ),
    .d(pnumcntA[3]),
    .e(\U_AHB/h2h_hrdata [3]),
    .o(_al_u3161_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((E*C)*~(B)*~(D)+(E*C)*B*~(D)+~((E*C))*B*D+(E*C)*B*D))"),
    .INIT(32'h220a22aa))
    _al_u3162 (
    .a(_al_u3061_o),
    .b(pnumcntB[3]),
    .c(pnumcntC[3]),
    .d(\U_AHB/h2h_haddr [2]),
    .e(\U_AHB/h2h_haddr [3]),
    .o(_al_u3162_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3163 (
    .a(_al_u3162_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcntD[3]),
    .e(pnumcntE[3]),
    .o(_al_u3163_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3164 (
    .a(_al_u3163_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcntF[3]),
    .e(pwm_state_read[3]),
    .o(_al_u3164_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*C)*~(D*B))"),
    .INIT(32'h020a22aa))
    _al_u3165 (
    .a(_al_u3164_o),
    .b(\U_AHB/n104_lutinv ),
    .c(\U_AHB/n102 ),
    .d(\U_AHB/h2h_hrdata [3]),
    .e(limit_r_pad[3]),
    .o(_al_u3165_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h33533050))
    _al_u3166 (
    .a(_al_u3161_o),
    .b(_al_u3165_o),
    .c(_al_u3061_o),
    .d(\U_AHB/h2h_haddr [13]),
    .e(\U_AHB/h2h_hrdata [3]),
    .o(\U_AHB/n118 [3]));
  AL_MAP_LUT4 #(
    .EQN("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    .INIT(16'h535f))
    _al_u3167 (
    .a(pnumcnt0[23]),
    .b(pnumcnt1[23]),
    .c(\U_AHB/h2h_haddr [2]),
    .d(\U_AHB/h2h_haddr [3]),
    .o(_al_u3167_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3168 (
    .a(_al_u3167_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcnt2[23]),
    .e(pnumcnt3[23]),
    .o(_al_u3168_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3169 (
    .a(_al_u3168_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcnt4[23]),
    .e(pnumcnt5[23]),
    .o(_al_u3169_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u317 (
    .a(\PWM4/pnumr [9]),
    .b(pnum4[32]),
    .c(pnum4[9]),
    .d(pwm_start_stop[20]),
    .o(\PWM4/n23 [9]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3170 (
    .a(_al_u3169_o),
    .b(\U_AHB/n102 ),
    .c(\U_AHB/n99 ),
    .d(pnumcnt6[23]),
    .e(pnumcnt7[23]),
    .o(_al_u3170_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3171 (
    .a(_al_u3170_o),
    .b(\U_AHB/n108 ),
    .c(\U_AHB/n105 ),
    .d(pnumcnt8[23]),
    .e(pnumcnt9[23]),
    .o(_al_u3171_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3172 (
    .a(_al_u3171_o),
    .b(\U_AHB/n113_lutinv ),
    .c(\U_AHB/n111 ),
    .d(pnumcntA[23]),
    .e(\U_AHB/h2h_hrdata [23]),
    .o(_al_u3172_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((E*C)*~(B)*~(D)+(E*C)*B*~(D)+~((E*C))*B*D+(E*C)*B*D))"),
    .INIT(32'h220a22aa))
    _al_u3173 (
    .a(_al_u3061_o),
    .b(pnumcntB[23]),
    .c(pnumcntC[23]),
    .d(\U_AHB/h2h_haddr [2]),
    .e(\U_AHB/h2h_haddr [3]),
    .o(_al_u3173_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3174 (
    .a(_al_u3173_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcntD[23]),
    .e(pnumcntE[23]),
    .o(_al_u3174_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3175 (
    .a(_al_u3174_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcntF[23]),
    .e(pwm_state_read[7]),
    .o(_al_u3175_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*C)*~(D*B))"),
    .INIT(32'h020a22aa))
    _al_u3176 (
    .a(_al_u3175_o),
    .b(\U_AHB/n104_lutinv ),
    .c(\U_AHB/n102 ),
    .d(\U_AHB/h2h_hrdata [23]),
    .e(limit_l_pad[7]),
    .o(_al_u3176_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h33533050))
    _al_u3177 (
    .a(_al_u3172_o),
    .b(_al_u3176_o),
    .c(_al_u3061_o),
    .d(\U_AHB/h2h_haddr [13]),
    .e(\U_AHB/h2h_hrdata [23]),
    .o(\U_AHB/n118 [23]));
  AL_MAP_LUT4 #(
    .EQN("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    .INIT(16'h535f))
    _al_u3178 (
    .a(pnumcnt0[22]),
    .b(pnumcnt1[22]),
    .c(\U_AHB/h2h_haddr [2]),
    .d(\U_AHB/h2h_haddr [3]),
    .o(_al_u3178_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3179 (
    .a(_al_u3178_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcnt2[22]),
    .e(pnumcnt3[22]),
    .o(_al_u3179_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u318 (
    .a(\PWM4/pnumr [8]),
    .b(pnum4[32]),
    .c(pnum4[8]),
    .d(pwm_start_stop[20]),
    .o(\PWM4/n23 [8]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3180 (
    .a(_al_u3179_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcnt4[22]),
    .e(pnumcnt5[22]),
    .o(_al_u3180_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3181 (
    .a(_al_u3180_o),
    .b(\U_AHB/n102 ),
    .c(\U_AHB/n99 ),
    .d(pnumcnt6[22]),
    .e(pnumcnt7[22]),
    .o(_al_u3181_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3182 (
    .a(_al_u3181_o),
    .b(\U_AHB/n108 ),
    .c(\U_AHB/n105 ),
    .d(pnumcnt8[22]),
    .e(pnumcnt9[22]),
    .o(_al_u3182_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3183 (
    .a(_al_u3182_o),
    .b(\U_AHB/n113_lutinv ),
    .c(\U_AHB/n111 ),
    .d(pnumcntA[22]),
    .e(\U_AHB/h2h_hrdata [22]),
    .o(_al_u3183_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((E*C)*~(B)*~(D)+(E*C)*B*~(D)+~((E*C))*B*D+(E*C)*B*D))"),
    .INIT(32'h220a22aa))
    _al_u3184 (
    .a(_al_u3061_o),
    .b(pnumcntB[22]),
    .c(pnumcntC[22]),
    .d(\U_AHB/h2h_haddr [2]),
    .e(\U_AHB/h2h_haddr [3]),
    .o(_al_u3184_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3185 (
    .a(_al_u3184_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcntD[22]),
    .e(pnumcntE[22]),
    .o(_al_u3185_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3186 (
    .a(_al_u3185_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcntF[22]),
    .e(pwm_state_read[6]),
    .o(_al_u3186_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*C)*~(D*B))"),
    .INIT(32'h020a22aa))
    _al_u3187 (
    .a(_al_u3186_o),
    .b(\U_AHB/n104_lutinv ),
    .c(\U_AHB/n102 ),
    .d(\U_AHB/h2h_hrdata [22]),
    .e(limit_l_pad[6]),
    .o(_al_u3187_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h33533050))
    _al_u3188 (
    .a(_al_u3183_o),
    .b(_al_u3187_o),
    .c(_al_u3061_o),
    .d(\U_AHB/h2h_haddr [13]),
    .e(\U_AHB/h2h_hrdata [22]),
    .o(\U_AHB/n118 [22]));
  AL_MAP_LUT4 #(
    .EQN("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    .INIT(16'h535f))
    _al_u3189 (
    .a(pnumcnt0[21]),
    .b(pnumcnt1[21]),
    .c(\U_AHB/h2h_haddr [2]),
    .d(\U_AHB/h2h_haddr [3]),
    .o(_al_u3189_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u319 (
    .a(\PWM4/pnumr [7]),
    .b(pnum4[32]),
    .c(pnum4[7]),
    .d(pwm_start_stop[20]),
    .o(\PWM4/n23 [7]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3190 (
    .a(_al_u3189_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcnt2[21]),
    .e(pnumcnt3[21]),
    .o(_al_u3190_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3191 (
    .a(_al_u3190_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcnt4[21]),
    .e(pnumcnt5[21]),
    .o(_al_u3191_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3192 (
    .a(_al_u3191_o),
    .b(\U_AHB/n102 ),
    .c(\U_AHB/n99 ),
    .d(pnumcnt6[21]),
    .e(pnumcnt7[21]),
    .o(_al_u3192_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3193 (
    .a(_al_u3192_o),
    .b(\U_AHB/n108 ),
    .c(\U_AHB/n105 ),
    .d(pnumcnt8[21]),
    .e(pnumcnt9[21]),
    .o(_al_u3193_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3194 (
    .a(_al_u3193_o),
    .b(\U_AHB/n113_lutinv ),
    .c(\U_AHB/n111 ),
    .d(pnumcntA[21]),
    .e(\U_AHB/h2h_hrdata [21]),
    .o(_al_u3194_o));
  AL_MAP_LUT4 #(
    .EQN("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    .INIT(16'h535f))
    _al_u3195 (
    .a(pnumcntB[21]),
    .b(pnumcntC[21]),
    .c(\U_AHB/h2h_haddr [2]),
    .d(\U_AHB/h2h_haddr [3]),
    .o(_al_u3195_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3196 (
    .a(_al_u3195_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcntD[21]),
    .e(pnumcntE[21]),
    .o(_al_u3196_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u3197 (
    .a(_al_u3139_o),
    .b(_al_u3196_o),
    .c(\U_AHB/n93 ),
    .d(pnumcntF[21]),
    .o(_al_u3197_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*C)*~(D*B))"),
    .INIT(32'h020a22aa))
    _al_u3198 (
    .a(_al_u3197_o),
    .b(\U_AHB/n104_lutinv ),
    .c(\U_AHB/n102 ),
    .d(\U_AHB/h2h_hrdata [21]),
    .e(limit_l_pad[5]),
    .o(_al_u3198_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h33533050))
    _al_u3199 (
    .a(_al_u3194_o),
    .b(_al_u3198_o),
    .c(_al_u3061_o),
    .d(\U_AHB/h2h_haddr [13]),
    .e(\U_AHB/h2h_hrdata [21]),
    .o(\U_AHB/n118 [21]));
  EF2_PHY_SPAD #(
    //.LOCATION("P24"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("16"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u32 (
    .do({open_n948,dir_pad[6]}),
    .ts(1'b1),
    .opad(dir[6]));  // CPLD_SOC_AHB_TOP.v(7)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u320 (
    .a(\PWM4/pnumr [6]),
    .b(pnum4[32]),
    .c(pnum4[6]),
    .d(pwm_start_stop[20]),
    .o(\PWM4/n23 [6]));
  AL_MAP_LUT4 #(
    .EQN("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    .INIT(16'h535f))
    _al_u3200 (
    .a(pnumcnt0[20]),
    .b(pnumcnt1[20]),
    .c(\U_AHB/h2h_haddr [2]),
    .d(\U_AHB/h2h_haddr [3]),
    .o(_al_u3200_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3201 (
    .a(_al_u3200_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcnt2[20]),
    .e(pnumcnt3[20]),
    .o(_al_u3201_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3202 (
    .a(_al_u3201_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcnt4[20]),
    .e(pnumcnt5[20]),
    .o(_al_u3202_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3203 (
    .a(_al_u3202_o),
    .b(\U_AHB/n102 ),
    .c(\U_AHB/n99 ),
    .d(pnumcnt6[20]),
    .e(pnumcnt7[20]),
    .o(_al_u3203_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3204 (
    .a(_al_u3203_o),
    .b(\U_AHB/n108 ),
    .c(\U_AHB/n105 ),
    .d(pnumcnt8[20]),
    .e(pnumcnt9[20]),
    .o(_al_u3204_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3205 (
    .a(_al_u3204_o),
    .b(\U_AHB/n113_lutinv ),
    .c(\U_AHB/n111 ),
    .d(pnumcntA[20]),
    .e(\U_AHB/h2h_hrdata [20]),
    .o(_al_u3205_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((E*C)*~(B)*~(D)+(E*C)*B*~(D)+~((E*C))*B*D+(E*C)*B*D))"),
    .INIT(32'h220a22aa))
    _al_u3206 (
    .a(_al_u3061_o),
    .b(pnumcntB[20]),
    .c(pnumcntC[20]),
    .d(\U_AHB/h2h_haddr [2]),
    .e(\U_AHB/h2h_haddr [3]),
    .o(_al_u3206_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3207 (
    .a(_al_u3206_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcntD[20]),
    .e(pnumcntE[20]),
    .o(_al_u3207_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3208 (
    .a(_al_u3207_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcntF[20]),
    .e(pwm_state_read[4]),
    .o(_al_u3208_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*C)*~(D*B))"),
    .INIT(32'h020a22aa))
    _al_u3209 (
    .a(_al_u3208_o),
    .b(\U_AHB/n104_lutinv ),
    .c(\U_AHB/n102 ),
    .d(\U_AHB/h2h_hrdata [20]),
    .e(limit_l_pad[4]),
    .o(_al_u3209_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u321 (
    .a(\PWM4/pnumr [5]),
    .b(pnum4[32]),
    .c(pnum4[5]),
    .d(pwm_start_stop[20]),
    .o(\PWM4/n23 [5]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h33533050))
    _al_u3210 (
    .a(_al_u3205_o),
    .b(_al_u3209_o),
    .c(_al_u3061_o),
    .d(\U_AHB/h2h_haddr [13]),
    .e(\U_AHB/h2h_hrdata [20]),
    .o(\U_AHB/n118 [20]));
  AL_MAP_LUT4 #(
    .EQN("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    .INIT(16'h535f))
    _al_u3211 (
    .a(pnumcnt0[2]),
    .b(pnumcnt1[2]),
    .c(\U_AHB/h2h_haddr [2]),
    .d(\U_AHB/h2h_haddr [3]),
    .o(_al_u3211_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3212 (
    .a(_al_u3211_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcnt2[2]),
    .e(pnumcnt3[2]),
    .o(_al_u3212_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3213 (
    .a(_al_u3212_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcnt4[2]),
    .e(pnumcnt5[2]),
    .o(_al_u3213_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3214 (
    .a(_al_u3213_o),
    .b(\U_AHB/n102 ),
    .c(\U_AHB/n99 ),
    .d(pnumcnt6[2]),
    .e(pnumcnt7[2]),
    .o(_al_u3214_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3215 (
    .a(_al_u3214_o),
    .b(\U_AHB/n108 ),
    .c(\U_AHB/n105 ),
    .d(pnumcnt8[2]),
    .e(pnumcnt9[2]),
    .o(_al_u3215_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3216 (
    .a(_al_u3215_o),
    .b(\U_AHB/n113_lutinv ),
    .c(\U_AHB/n111 ),
    .d(pnumcntA[2]),
    .e(\U_AHB/h2h_hrdata [2]),
    .o(_al_u3216_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((E*C)*~(B)*~(D)+(E*C)*B*~(D)+~((E*C))*B*D+(E*C)*B*D))"),
    .INIT(32'h220a22aa))
    _al_u3217 (
    .a(_al_u3061_o),
    .b(pnumcntB[2]),
    .c(pnumcntC[2]),
    .d(\U_AHB/h2h_haddr [2]),
    .e(\U_AHB/h2h_haddr [3]),
    .o(_al_u3217_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3218 (
    .a(_al_u3217_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcntD[2]),
    .e(pnumcntE[2]),
    .o(_al_u3218_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3219 (
    .a(_al_u3218_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcntF[2]),
    .e(pwm_state_read[2]),
    .o(_al_u3219_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u322 (
    .a(\PWM4/pnumr [4]),
    .b(pnum4[32]),
    .c(pnum4[4]),
    .d(pwm_start_stop[20]),
    .o(\PWM4/n23 [4]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*C)*~(D*B))"),
    .INIT(32'h020a22aa))
    _al_u3220 (
    .a(_al_u3219_o),
    .b(\U_AHB/n104_lutinv ),
    .c(\U_AHB/n102 ),
    .d(\U_AHB/h2h_hrdata [2]),
    .e(limit_r_pad[2]),
    .o(_al_u3220_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h33533050))
    _al_u3221 (
    .a(_al_u3216_o),
    .b(_al_u3220_o),
    .c(_al_u3061_o),
    .d(\U_AHB/h2h_haddr [13]),
    .e(\U_AHB/h2h_hrdata [2]),
    .o(\U_AHB/n118 [2]));
  AL_MAP_LUT4 #(
    .EQN("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    .INIT(16'h535f))
    _al_u3222 (
    .a(pnumcnt0[19]),
    .b(pnumcnt1[19]),
    .c(\U_AHB/h2h_haddr [2]),
    .d(\U_AHB/h2h_haddr [3]),
    .o(_al_u3222_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3223 (
    .a(_al_u3222_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcnt2[19]),
    .e(pnumcnt3[19]),
    .o(_al_u3223_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3224 (
    .a(_al_u3223_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcnt4[19]),
    .e(pnumcnt5[19]),
    .o(_al_u3224_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3225 (
    .a(_al_u3224_o),
    .b(\U_AHB/n102 ),
    .c(\U_AHB/n99 ),
    .d(pnumcnt6[19]),
    .e(pnumcnt7[19]),
    .o(_al_u3225_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3226 (
    .a(_al_u3225_o),
    .b(\U_AHB/n108 ),
    .c(\U_AHB/n105 ),
    .d(pnumcnt8[19]),
    .e(pnumcnt9[19]),
    .o(_al_u3226_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3227 (
    .a(_al_u3226_o),
    .b(\U_AHB/n113_lutinv ),
    .c(\U_AHB/n111 ),
    .d(pnumcntA[19]),
    .e(\U_AHB/h2h_hrdata [19]),
    .o(_al_u3227_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((E*C)*~(B)*~(D)+(E*C)*B*~(D)+~((E*C))*B*D+(E*C)*B*D))"),
    .INIT(32'h220a22aa))
    _al_u3228 (
    .a(_al_u3061_o),
    .b(pnumcntB[19]),
    .c(pnumcntC[19]),
    .d(\U_AHB/h2h_haddr [2]),
    .e(\U_AHB/h2h_haddr [3]),
    .o(_al_u3228_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3229 (
    .a(_al_u3228_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcntD[19]),
    .e(pnumcntE[19]),
    .o(_al_u3229_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u323 (
    .a(\PWM4/pnumr [31]),
    .b(pnum4[31]),
    .c(pnum4[32]),
    .d(pwm_start_stop[20]),
    .o(\PWM4/n23 [31]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3230 (
    .a(_al_u3229_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcntF[19]),
    .e(pwm_state_read[3]),
    .o(_al_u3230_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*C)*~(D*B))"),
    .INIT(32'h020a22aa))
    _al_u3231 (
    .a(_al_u3230_o),
    .b(\U_AHB/n104_lutinv ),
    .c(\U_AHB/n102 ),
    .d(\U_AHB/h2h_hrdata [19]),
    .e(limit_l_pad[3]),
    .o(_al_u3231_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h33533050))
    _al_u3232 (
    .a(_al_u3227_o),
    .b(_al_u3231_o),
    .c(_al_u3061_o),
    .d(\U_AHB/h2h_haddr [13]),
    .e(\U_AHB/h2h_hrdata [19]),
    .o(\U_AHB/n118 [19]));
  AL_MAP_LUT5 #(
    .EQN("(A*~((E*C)*~(B)*~(D)+(E*C)*B*~(D)+~((E*C))*B*D+(E*C)*B*D))"),
    .INIT(32'h220a22aa))
    _al_u3233 (
    .a(\U_AHB/n82 ),
    .b(pnumcnt0[18]),
    .c(pnumcnt1[18]),
    .d(\U_AHB/h2h_haddr [2]),
    .e(\U_AHB/h2h_haddr [3]),
    .o(_al_u3233_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3234 (
    .a(_al_u3233_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcnt2[18]),
    .e(pnumcnt3[18]),
    .o(_al_u3234_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3235 (
    .a(_al_u3234_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcnt4[18]),
    .e(pnumcnt5[18]),
    .o(_al_u3235_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3236 (
    .a(_al_u3235_o),
    .b(\U_AHB/n102 ),
    .c(\U_AHB/n99 ),
    .d(pnumcnt6[18]),
    .e(pnumcnt7[18]),
    .o(_al_u3236_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3237 (
    .a(_al_u3236_o),
    .b(\U_AHB/n108 ),
    .c(\U_AHB/n105 ),
    .d(pnumcnt8[18]),
    .e(pnumcnt9[18]),
    .o(_al_u3237_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C))"),
    .INIT(32'h535f0000))
    _al_u3238 (
    .a(pnumcntB[18]),
    .b(pnumcntC[18]),
    .c(\U_AHB/h2h_haddr [2]),
    .d(\U_AHB/h2h_haddr [3]),
    .e(\U_AHB/h2h_haddr [13]),
    .o(_al_u3238_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3239 (
    .a(_al_u3238_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcntD[18]),
    .e(pnumcntE[18]),
    .o(_al_u3239_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u324 (
    .a(\PWM4/pnumr [30]),
    .b(pnum4[30]),
    .c(pnum4[32]),
    .d(pwm_start_stop[20]),
    .o(\PWM4/n23 [30]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3240 (
    .a(_al_u3239_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcntF[18]),
    .e(pwm_state_read[2]),
    .o(_al_u3240_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(D*B)))"),
    .INIT(16'hd050))
    _al_u3241 (
    .a(_al_u3240_o),
    .b(\U_AHB/n102 ),
    .c(_al_u3061_o),
    .d(limit_l_pad[2]),
    .o(_al_u3241_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u3242 (
    .a(\U_AHB/n113_lutinv ),
    .b(\U_AHB/n111 ),
    .c(pnumcntA[18]),
    .d(\U_AHB/h2h_hrdata [18]),
    .o(_al_u3242_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~(E*~D)*~B)*~(C*A))"),
    .INIT(32'h4c5f4c4c))
    _al_u3243 (
    .a(_al_u3237_o),
    .b(_al_u3241_o),
    .c(_al_u3242_o),
    .d(_al_u3065_o),
    .e(\U_AHB/h2h_hrdata [18]),
    .o(\U_AHB/n118 [18]));
  AL_MAP_LUT4 #(
    .EQN("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    .INIT(16'h535f))
    _al_u3244 (
    .a(pnumcnt0[17]),
    .b(pnumcnt1[17]),
    .c(\U_AHB/h2h_haddr [2]),
    .d(\U_AHB/h2h_haddr [3]),
    .o(_al_u3244_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3245 (
    .a(_al_u3244_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcnt2[17]),
    .e(pnumcnt3[17]),
    .o(_al_u3245_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3246 (
    .a(_al_u3245_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcnt4[17]),
    .e(pnumcnt5[17]),
    .o(_al_u3246_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3247 (
    .a(_al_u3246_o),
    .b(\U_AHB/n102 ),
    .c(\U_AHB/n99 ),
    .d(pnumcnt6[17]),
    .e(pnumcnt7[17]),
    .o(_al_u3247_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3248 (
    .a(_al_u3247_o),
    .b(\U_AHB/n108 ),
    .c(\U_AHB/n105 ),
    .d(pnumcnt8[17]),
    .e(pnumcnt9[17]),
    .o(_al_u3248_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3249 (
    .a(_al_u3248_o),
    .b(\U_AHB/n113_lutinv ),
    .c(\U_AHB/n111 ),
    .d(pnumcntA[17]),
    .e(\U_AHB/h2h_hrdata [17]),
    .o(_al_u3249_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u325 (
    .a(\PWM4/pnumr [3]),
    .b(pnum4[3]),
    .c(pnum4[32]),
    .d(pwm_start_stop[20]),
    .o(\PWM4/n23 [3]));
  AL_MAP_LUT5 #(
    .EQN("(A*~((E*C)*~(B)*~(D)+(E*C)*B*~(D)+~((E*C))*B*D+(E*C)*B*D))"),
    .INIT(32'h220a22aa))
    _al_u3250 (
    .a(_al_u3061_o),
    .b(pnumcntB[17]),
    .c(pnumcntC[17]),
    .d(\U_AHB/h2h_haddr [2]),
    .e(\U_AHB/h2h_haddr [3]),
    .o(_al_u3250_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3251 (
    .a(_al_u3250_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcntD[17]),
    .e(pnumcntE[17]),
    .o(_al_u3251_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3252 (
    .a(_al_u3251_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcntF[17]),
    .e(pwm_state_read[1]),
    .o(_al_u3252_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*C)*~(D*B))"),
    .INIT(32'h020a22aa))
    _al_u3253 (
    .a(_al_u3252_o),
    .b(\U_AHB/n104_lutinv ),
    .c(\U_AHB/n102 ),
    .d(\U_AHB/h2h_hrdata [17]),
    .e(limit_l_pad[1]),
    .o(_al_u3253_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h33533050))
    _al_u3254 (
    .a(_al_u3249_o),
    .b(_al_u3253_o),
    .c(_al_u3061_o),
    .d(\U_AHB/h2h_haddr [13]),
    .e(\U_AHB/h2h_hrdata [17]),
    .o(\U_AHB/n118 [17]));
  AL_MAP_LUT4 #(
    .EQN("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    .INIT(16'h535f))
    _al_u3255 (
    .a(pnumcnt0[16]),
    .b(pnumcnt1[16]),
    .c(\U_AHB/h2h_haddr [2]),
    .d(\U_AHB/h2h_haddr [3]),
    .o(_al_u3255_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3256 (
    .a(_al_u3255_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcnt2[16]),
    .e(pnumcnt3[16]),
    .o(_al_u3256_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3257 (
    .a(_al_u3256_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcnt4[16]),
    .e(pnumcnt5[16]),
    .o(_al_u3257_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3258 (
    .a(_al_u3257_o),
    .b(\U_AHB/n102 ),
    .c(\U_AHB/n99 ),
    .d(pnumcnt6[16]),
    .e(pnumcnt7[16]),
    .o(_al_u3258_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3259 (
    .a(_al_u3258_o),
    .b(\U_AHB/n108 ),
    .c(\U_AHB/n105 ),
    .d(pnumcnt8[16]),
    .e(pnumcnt9[16]),
    .o(_al_u3259_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u326 (
    .a(\PWM4/pnumr [29]),
    .b(pnum4[29]),
    .c(pnum4[32]),
    .d(pwm_start_stop[20]),
    .o(\PWM4/n23 [29]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3260 (
    .a(_al_u3259_o),
    .b(\U_AHB/n113_lutinv ),
    .c(\U_AHB/n111 ),
    .d(pnumcntA[16]),
    .e(\U_AHB/h2h_hrdata [16]),
    .o(_al_u3260_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((E*C)*~(B)*~(D)+(E*C)*B*~(D)+~((E*C))*B*D+(E*C)*B*D))"),
    .INIT(32'h220a22aa))
    _al_u3261 (
    .a(_al_u3061_o),
    .b(pnumcntB[16]),
    .c(pnumcntC[16]),
    .d(\U_AHB/h2h_haddr [2]),
    .e(\U_AHB/h2h_haddr [3]),
    .o(_al_u3261_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3262 (
    .a(_al_u3261_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcntD[16]),
    .e(pnumcntE[16]),
    .o(_al_u3262_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3263 (
    .a(_al_u3262_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcntF[16]),
    .e(pwm_state_read[0]),
    .o(_al_u3263_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*C)*~(D*B))"),
    .INIT(32'h020a22aa))
    _al_u3264 (
    .a(_al_u3263_o),
    .b(\U_AHB/n104_lutinv ),
    .c(\U_AHB/n102 ),
    .d(\U_AHB/h2h_hrdata [16]),
    .e(limit_l_pad[0]),
    .o(_al_u3264_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h33533050))
    _al_u3265 (
    .a(_al_u3260_o),
    .b(_al_u3264_o),
    .c(_al_u3061_o),
    .d(\U_AHB/h2h_haddr [13]),
    .e(\U_AHB/h2h_hrdata [16]),
    .o(\U_AHB/n118 [16]));
  AL_MAP_LUT4 #(
    .EQN("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    .INIT(16'h535f))
    _al_u3266 (
    .a(pnumcnt0[15]),
    .b(pnumcnt1[15]),
    .c(\U_AHB/h2h_haddr [2]),
    .d(\U_AHB/h2h_haddr [3]),
    .o(_al_u3266_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3267 (
    .a(_al_u3266_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcnt2[15]),
    .e(pnumcnt3[15]),
    .o(_al_u3267_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3268 (
    .a(_al_u3267_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcnt4[15]),
    .e(pnumcnt5[15]),
    .o(_al_u3268_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3269 (
    .a(_al_u3268_o),
    .b(\U_AHB/n102 ),
    .c(\U_AHB/n99 ),
    .d(pnumcnt6[15]),
    .e(pnumcnt7[15]),
    .o(_al_u3269_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u327 (
    .a(\PWM4/pnumr [28]),
    .b(pnum4[28]),
    .c(pnum4[32]),
    .d(pwm_start_stop[20]),
    .o(\PWM4/n23 [28]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3270 (
    .a(_al_u3269_o),
    .b(\U_AHB/n108 ),
    .c(\U_AHB/n105 ),
    .d(pnumcnt8[15]),
    .e(pnumcnt9[15]),
    .o(_al_u3270_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3271 (
    .a(_al_u3270_o),
    .b(\U_AHB/n113_lutinv ),
    .c(\U_AHB/n111 ),
    .d(pnumcntA[15]),
    .e(\U_AHB/h2h_hrdata [15]),
    .o(_al_u3271_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((E*C)*~(B)*~(D)+(E*C)*B*~(D)+~((E*C))*B*D+(E*C)*B*D))"),
    .INIT(32'h220a22aa))
    _al_u3272 (
    .a(_al_u3061_o),
    .b(pnumcntB[15]),
    .c(pnumcntC[15]),
    .d(\U_AHB/h2h_haddr [2]),
    .e(\U_AHB/h2h_haddr [3]),
    .o(_al_u3272_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3273 (
    .a(_al_u3272_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcntD[15]),
    .e(pnumcntE[15]),
    .o(_al_u3273_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3274 (
    .a(_al_u3273_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcntF[15]),
    .e(pwm_state_read[15]),
    .o(_al_u3274_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*C)*~(D*B))"),
    .INIT(32'h020a22aa))
    _al_u3275 (
    .a(_al_u3274_o),
    .b(\U_AHB/n104_lutinv ),
    .c(\U_AHB/n102 ),
    .d(\U_AHB/h2h_hrdata [15]),
    .e(limit_r_pad[15]),
    .o(_al_u3275_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h33533050))
    _al_u3276 (
    .a(_al_u3271_o),
    .b(_al_u3275_o),
    .c(_al_u3061_o),
    .d(\U_AHB/h2h_haddr [13]),
    .e(\U_AHB/h2h_hrdata [15]),
    .o(\U_AHB/n118 [15]));
  AL_MAP_LUT4 #(
    .EQN("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    .INIT(16'h535f))
    _al_u3277 (
    .a(pnumcnt0[14]),
    .b(pnumcnt1[14]),
    .c(\U_AHB/h2h_haddr [2]),
    .d(\U_AHB/h2h_haddr [3]),
    .o(_al_u3277_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3278 (
    .a(_al_u3277_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcnt2[14]),
    .e(pnumcnt3[14]),
    .o(_al_u3278_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3279 (
    .a(_al_u3278_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcnt4[14]),
    .e(pnumcnt5[14]),
    .o(_al_u3279_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u328 (
    .a(\PWM4/pnumr [27]),
    .b(pnum4[27]),
    .c(pnum4[32]),
    .d(pwm_start_stop[20]),
    .o(\PWM4/n23 [27]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3280 (
    .a(_al_u3279_o),
    .b(\U_AHB/n102 ),
    .c(\U_AHB/n99 ),
    .d(pnumcnt6[14]),
    .e(pnumcnt7[14]),
    .o(_al_u3280_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3281 (
    .a(_al_u3280_o),
    .b(\U_AHB/n108 ),
    .c(\U_AHB/n105 ),
    .d(pnumcnt8[14]),
    .e(pnumcnt9[14]),
    .o(_al_u3281_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3282 (
    .a(_al_u3281_o),
    .b(\U_AHB/n113_lutinv ),
    .c(\U_AHB/n111 ),
    .d(pnumcntA[14]),
    .e(\U_AHB/h2h_hrdata [14]),
    .o(_al_u3282_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((E*C)*~(B)*~(D)+(E*C)*B*~(D)+~((E*C))*B*D+(E*C)*B*D))"),
    .INIT(32'h220a22aa))
    _al_u3283 (
    .a(_al_u3061_o),
    .b(pnumcntB[14]),
    .c(pnumcntC[14]),
    .d(\U_AHB/h2h_haddr [2]),
    .e(\U_AHB/h2h_haddr [3]),
    .o(_al_u3283_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3284 (
    .a(_al_u3283_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcntD[14]),
    .e(pnumcntE[14]),
    .o(_al_u3284_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3285 (
    .a(_al_u3284_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcntF[14]),
    .e(pwm_state_read[14]),
    .o(_al_u3285_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*C)*~(D*B))"),
    .INIT(32'h020a22aa))
    _al_u3286 (
    .a(_al_u3285_o),
    .b(\U_AHB/n104_lutinv ),
    .c(\U_AHB/n102 ),
    .d(\U_AHB/h2h_hrdata [14]),
    .e(limit_r_pad[14]),
    .o(_al_u3286_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h33533050))
    _al_u3287 (
    .a(_al_u3282_o),
    .b(_al_u3286_o),
    .c(_al_u3061_o),
    .d(\U_AHB/h2h_haddr [13]),
    .e(\U_AHB/h2h_hrdata [14]),
    .o(\U_AHB/n118 [14]));
  AL_MAP_LUT4 #(
    .EQN("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    .INIT(16'h535f))
    _al_u3288 (
    .a(pnumcnt0[13]),
    .b(pnumcnt1[13]),
    .c(\U_AHB/h2h_haddr [2]),
    .d(\U_AHB/h2h_haddr [3]),
    .o(_al_u3288_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3289 (
    .a(_al_u3288_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcnt2[13]),
    .e(pnumcnt3[13]),
    .o(_al_u3289_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u329 (
    .a(\PWM4/pnumr [26]),
    .b(pnum4[26]),
    .c(pnum4[32]),
    .d(pwm_start_stop[20]),
    .o(\PWM4/n23 [26]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3290 (
    .a(_al_u3289_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcnt4[13]),
    .e(pnumcnt5[13]),
    .o(_al_u3290_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3291 (
    .a(_al_u3290_o),
    .b(\U_AHB/n102 ),
    .c(\U_AHB/n99 ),
    .d(pnumcnt6[13]),
    .e(pnumcnt7[13]),
    .o(_al_u3291_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3292 (
    .a(_al_u3291_o),
    .b(\U_AHB/n108 ),
    .c(\U_AHB/n105 ),
    .d(pnumcnt8[13]),
    .e(pnumcnt9[13]),
    .o(_al_u3292_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3293 (
    .a(_al_u3292_o),
    .b(\U_AHB/n113_lutinv ),
    .c(\U_AHB/n111 ),
    .d(pnumcntA[13]),
    .e(\U_AHB/h2h_hrdata [13]),
    .o(_al_u3293_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((E*C)*~(B)*~(D)+(E*C)*B*~(D)+~((E*C))*B*D+(E*C)*B*D))"),
    .INIT(32'h220a22aa))
    _al_u3294 (
    .a(_al_u3061_o),
    .b(pnumcntB[13]),
    .c(pnumcntC[13]),
    .d(\U_AHB/h2h_haddr [2]),
    .e(\U_AHB/h2h_haddr [3]),
    .o(_al_u3294_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3295 (
    .a(_al_u3294_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcntD[13]),
    .e(pnumcntE[13]),
    .o(_al_u3295_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3296 (
    .a(_al_u3295_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcntF[13]),
    .e(pwm_state_read[13]),
    .o(_al_u3296_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*C)*~(D*B))"),
    .INIT(32'h020a22aa))
    _al_u3297 (
    .a(_al_u3296_o),
    .b(\U_AHB/n104_lutinv ),
    .c(\U_AHB/n102 ),
    .d(\U_AHB/h2h_hrdata [13]),
    .e(limit_r_pad[13]),
    .o(_al_u3297_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h33533050))
    _al_u3298 (
    .a(_al_u3293_o),
    .b(_al_u3297_o),
    .c(_al_u3061_o),
    .d(\U_AHB/h2h_haddr [13]),
    .e(\U_AHB/h2h_hrdata [13]),
    .o(\U_AHB/n118 [13]));
  AL_MAP_LUT4 #(
    .EQN("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    .INIT(16'h535f))
    _al_u3299 (
    .a(pnumcnt0[12]),
    .b(pnumcnt1[12]),
    .c(\U_AHB/h2h_haddr [2]),
    .d(\U_AHB/h2h_haddr [3]),
    .o(_al_u3299_o));
  EF2_PHY_SPAD #(
    //.LOCATION("P23"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("16"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u33 (
    .do({open_n957,dir_pad[5]}),
    .ts(1'b1),
    .opad(dir[5]));  // CPLD_SOC_AHB_TOP.v(7)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u330 (
    .a(\PWM4/pnumr [25]),
    .b(pnum4[25]),
    .c(pnum4[32]),
    .d(pwm_start_stop[20]),
    .o(\PWM4/n23 [25]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3300 (
    .a(_al_u3299_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcnt2[12]),
    .e(pnumcnt3[12]),
    .o(_al_u3300_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3301 (
    .a(_al_u3300_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcnt4[12]),
    .e(pnumcnt5[12]),
    .o(_al_u3301_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3302 (
    .a(_al_u3301_o),
    .b(\U_AHB/n102 ),
    .c(\U_AHB/n99 ),
    .d(pnumcnt6[12]),
    .e(pnumcnt7[12]),
    .o(_al_u3302_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3303 (
    .a(_al_u3302_o),
    .b(\U_AHB/n108 ),
    .c(\U_AHB/n105 ),
    .d(pnumcnt8[12]),
    .e(pnumcnt9[12]),
    .o(_al_u3303_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3304 (
    .a(_al_u3303_o),
    .b(\U_AHB/n113_lutinv ),
    .c(\U_AHB/n111 ),
    .d(pnumcntA[12]),
    .e(\U_AHB/h2h_hrdata [12]),
    .o(_al_u3304_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((E*C)*~(B)*~(D)+(E*C)*B*~(D)+~((E*C))*B*D+(E*C)*B*D))"),
    .INIT(32'h220a22aa))
    _al_u3305 (
    .a(_al_u3061_o),
    .b(pnumcntB[12]),
    .c(pnumcntC[12]),
    .d(\U_AHB/h2h_haddr [2]),
    .e(\U_AHB/h2h_haddr [3]),
    .o(_al_u3305_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3306 (
    .a(_al_u3305_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcntD[12]),
    .e(pnumcntE[12]),
    .o(_al_u3306_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3307 (
    .a(_al_u3306_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcntF[12]),
    .e(pwm_state_read[12]),
    .o(_al_u3307_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*C)*~(D*B))"),
    .INIT(32'h020a22aa))
    _al_u3308 (
    .a(_al_u3307_o),
    .b(\U_AHB/n104_lutinv ),
    .c(\U_AHB/n102 ),
    .d(\U_AHB/h2h_hrdata [12]),
    .e(limit_r_pad[12]),
    .o(_al_u3308_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h33533050))
    _al_u3309 (
    .a(_al_u3304_o),
    .b(_al_u3308_o),
    .c(_al_u3061_o),
    .d(\U_AHB/h2h_haddr [13]),
    .e(\U_AHB/h2h_hrdata [12]),
    .o(\U_AHB/n118 [12]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u331 (
    .a(\PWM4/pnumr [24]),
    .b(pnum4[24]),
    .c(pnum4[32]),
    .d(pwm_start_stop[20]),
    .o(\PWM4/n23 [24]));
  AL_MAP_LUT4 #(
    .EQN("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    .INIT(16'h535f))
    _al_u3310 (
    .a(pnumcnt0[11]),
    .b(pnumcnt1[11]),
    .c(\U_AHB/h2h_haddr [2]),
    .d(\U_AHB/h2h_haddr [3]),
    .o(_al_u3310_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3311 (
    .a(_al_u3310_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcnt2[11]),
    .e(pnumcnt3[11]),
    .o(_al_u3311_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3312 (
    .a(_al_u3311_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcnt4[11]),
    .e(pnumcnt5[11]),
    .o(_al_u3312_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3313 (
    .a(_al_u3312_o),
    .b(\U_AHB/n102 ),
    .c(\U_AHB/n99 ),
    .d(pnumcnt6[11]),
    .e(pnumcnt7[11]),
    .o(_al_u3313_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3314 (
    .a(_al_u3313_o),
    .b(\U_AHB/n108 ),
    .c(\U_AHB/n105 ),
    .d(pnumcnt8[11]),
    .e(pnumcnt9[11]),
    .o(_al_u3314_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3315 (
    .a(_al_u3314_o),
    .b(\U_AHB/n113_lutinv ),
    .c(\U_AHB/n111 ),
    .d(pnumcntA[11]),
    .e(\U_AHB/h2h_hrdata [11]),
    .o(_al_u3315_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((E*C)*~(B)*~(D)+(E*C)*B*~(D)+~((E*C))*B*D+(E*C)*B*D))"),
    .INIT(32'h220a22aa))
    _al_u3316 (
    .a(_al_u3061_o),
    .b(pnumcntB[11]),
    .c(pnumcntC[11]),
    .d(\U_AHB/h2h_haddr [2]),
    .e(\U_AHB/h2h_haddr [3]),
    .o(_al_u3316_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3317 (
    .a(_al_u3316_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcntD[11]),
    .e(pnumcntE[11]),
    .o(_al_u3317_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3318 (
    .a(_al_u3317_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcntF[11]),
    .e(pwm_state_read[11]),
    .o(_al_u3318_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*C)*~(D*B))"),
    .INIT(32'h020a22aa))
    _al_u3319 (
    .a(_al_u3318_o),
    .b(\U_AHB/n104_lutinv ),
    .c(\U_AHB/n102 ),
    .d(\U_AHB/h2h_hrdata [11]),
    .e(limit_r_pad[11]),
    .o(_al_u3319_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u332 (
    .a(\PWM4/pnumr [23]),
    .b(pnum4[23]),
    .c(pnum4[32]),
    .d(pwm_start_stop[20]),
    .o(\PWM4/n23 [23]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h33533050))
    _al_u3320 (
    .a(_al_u3315_o),
    .b(_al_u3319_o),
    .c(_al_u3061_o),
    .d(\U_AHB/h2h_haddr [13]),
    .e(\U_AHB/h2h_hrdata [11]),
    .o(\U_AHB/n118 [11]));
  AL_MAP_LUT4 #(
    .EQN("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    .INIT(16'h535f))
    _al_u3321 (
    .a(pnumcnt0[10]),
    .b(pnumcnt1[10]),
    .c(\U_AHB/h2h_haddr [2]),
    .d(\U_AHB/h2h_haddr [3]),
    .o(_al_u3321_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3322 (
    .a(_al_u3321_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcnt2[10]),
    .e(pnumcnt3[10]),
    .o(_al_u3322_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3323 (
    .a(_al_u3322_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcnt4[10]),
    .e(pnumcnt5[10]),
    .o(_al_u3323_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3324 (
    .a(_al_u3323_o),
    .b(\U_AHB/n102 ),
    .c(\U_AHB/n99 ),
    .d(pnumcnt6[10]),
    .e(pnumcnt7[10]),
    .o(_al_u3324_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3325 (
    .a(_al_u3324_o),
    .b(\U_AHB/n108 ),
    .c(\U_AHB/n105 ),
    .d(pnumcnt8[10]),
    .e(pnumcnt9[10]),
    .o(_al_u3325_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3326 (
    .a(_al_u3325_o),
    .b(\U_AHB/n113_lutinv ),
    .c(\U_AHB/n111 ),
    .d(pnumcntA[10]),
    .e(\U_AHB/h2h_hrdata [10]),
    .o(_al_u3326_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((E*C)*~(B)*~(D)+(E*C)*B*~(D)+~((E*C))*B*D+(E*C)*B*D))"),
    .INIT(32'h220a22aa))
    _al_u3327 (
    .a(_al_u3061_o),
    .b(pnumcntB[10]),
    .c(pnumcntC[10]),
    .d(\U_AHB/h2h_haddr [2]),
    .e(\U_AHB/h2h_haddr [3]),
    .o(_al_u3327_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3328 (
    .a(_al_u3327_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcntD[10]),
    .e(pnumcntE[10]),
    .o(_al_u3328_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3329 (
    .a(_al_u3328_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcntF[10]),
    .e(pwm_state_read[10]),
    .o(_al_u3329_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u333 (
    .a(\PWM4/pnumr [22]),
    .b(pnum4[22]),
    .c(pnum4[32]),
    .d(pwm_start_stop[20]),
    .o(\PWM4/n23 [22]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*C)*~(D*B))"),
    .INIT(32'h020a22aa))
    _al_u3330 (
    .a(_al_u3329_o),
    .b(\U_AHB/n104_lutinv ),
    .c(\U_AHB/n102 ),
    .d(\U_AHB/h2h_hrdata [10]),
    .e(limit_r_pad[10]),
    .o(_al_u3330_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h33533050))
    _al_u3331 (
    .a(_al_u3326_o),
    .b(_al_u3330_o),
    .c(_al_u3061_o),
    .d(\U_AHB/h2h_haddr [13]),
    .e(\U_AHB/h2h_hrdata [10]),
    .o(\U_AHB/n118 [10]));
  AL_MAP_LUT4 #(
    .EQN("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    .INIT(16'h535f))
    _al_u3332 (
    .a(pnumcnt0[1]),
    .b(pnumcnt1[1]),
    .c(\U_AHB/h2h_haddr [2]),
    .d(\U_AHB/h2h_haddr [3]),
    .o(_al_u3332_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3333 (
    .a(_al_u3332_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcnt2[1]),
    .e(pnumcnt3[1]),
    .o(_al_u3333_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3334 (
    .a(_al_u3333_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcnt4[1]),
    .e(pnumcnt5[1]),
    .o(_al_u3334_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3335 (
    .a(_al_u3334_o),
    .b(\U_AHB/n102 ),
    .c(\U_AHB/n99 ),
    .d(pnumcnt6[1]),
    .e(pnumcnt7[1]),
    .o(_al_u3335_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3336 (
    .a(_al_u3335_o),
    .b(\U_AHB/n108 ),
    .c(\U_AHB/n105 ),
    .d(pnumcnt8[1]),
    .e(pnumcnt9[1]),
    .o(_al_u3336_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3337 (
    .a(_al_u3336_o),
    .b(\U_AHB/n113_lutinv ),
    .c(\U_AHB/n111 ),
    .d(pnumcntA[1]),
    .e(\U_AHB/h2h_hrdata [1]),
    .o(_al_u3337_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((E*C)*~(B)*~(D)+(E*C)*B*~(D)+~((E*C))*B*D+(E*C)*B*D))"),
    .INIT(32'h220a22aa))
    _al_u3338 (
    .a(_al_u3061_o),
    .b(pnumcntB[1]),
    .c(pnumcntC[1]),
    .d(\U_AHB/h2h_haddr [2]),
    .e(\U_AHB/h2h_haddr [3]),
    .o(_al_u3338_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3339 (
    .a(_al_u3338_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcntD[1]),
    .e(pnumcntE[1]),
    .o(_al_u3339_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u334 (
    .a(\PWM4/pnumr [21]),
    .b(pnum4[21]),
    .c(pnum4[32]),
    .d(pwm_start_stop[20]),
    .o(\PWM4/n23 [21]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3340 (
    .a(_al_u3339_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcntF[1]),
    .e(pwm_state_read[1]),
    .o(_al_u3340_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*C)*~(D*B))"),
    .INIT(32'h020a22aa))
    _al_u3341 (
    .a(_al_u3340_o),
    .b(\U_AHB/n104_lutinv ),
    .c(\U_AHB/n102 ),
    .d(\U_AHB/h2h_hrdata [1]),
    .e(limit_r_pad[1]),
    .o(_al_u3341_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h33533050))
    _al_u3342 (
    .a(_al_u3337_o),
    .b(_al_u3341_o),
    .c(_al_u3061_o),
    .d(\U_AHB/h2h_haddr [13]),
    .e(\U_AHB/h2h_hrdata [1]),
    .o(\U_AHB/n118 [1]));
  AL_MAP_LUT4 #(
    .EQN("~((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    .INIT(16'h535f))
    _al_u3343 (
    .a(pnumcnt0[0]),
    .b(pnumcnt1[0]),
    .c(\U_AHB/h2h_haddr [2]),
    .d(\U_AHB/h2h_haddr [3]),
    .o(_al_u3343_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3344 (
    .a(_al_u3343_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcnt2[0]),
    .e(pnumcnt3[0]),
    .o(_al_u3344_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3345 (
    .a(_al_u3344_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcnt4[0]),
    .e(pnumcnt5[0]),
    .o(_al_u3345_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3346 (
    .a(_al_u3345_o),
    .b(\U_AHB/n102 ),
    .c(\U_AHB/n99 ),
    .d(pnumcnt6[0]),
    .e(pnumcnt7[0]),
    .o(_al_u3346_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3347 (
    .a(_al_u3346_o),
    .b(\U_AHB/n108 ),
    .c(\U_AHB/n105 ),
    .d(pnumcnt8[0]),
    .e(pnumcnt9[0]),
    .o(_al_u3347_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3348 (
    .a(_al_u3347_o),
    .b(\U_AHB/n113_lutinv ),
    .c(\U_AHB/n111 ),
    .d(pnumcntA[0]),
    .e(\U_AHB/h2h_hrdata [0]),
    .o(_al_u3348_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((E*C)*~(B)*~(D)+(E*C)*B*~(D)+~((E*C))*B*D+(E*C)*B*D))"),
    .INIT(32'h220a22aa))
    _al_u3349 (
    .a(_al_u3061_o),
    .b(pnumcntB[0]),
    .c(pnumcntC[0]),
    .d(\U_AHB/h2h_haddr [2]),
    .e(\U_AHB/h2h_haddr [3]),
    .o(_al_u3349_o));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u335 (
    .a(\PWM4/pnumr [20]),
    .b(pnum4[20]),
    .c(pnum4[32]),
    .d(pwm_start_stop[20]),
    .o(\PWM4/n23 [20]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3350 (
    .a(_al_u3349_o),
    .b(\U_AHB/n90 ),
    .c(\U_AHB/n87 ),
    .d(pnumcntD[0]),
    .e(pnumcntE[0]),
    .o(_al_u3350_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u3351 (
    .a(_al_u3350_o),
    .b(\U_AHB/n96 ),
    .c(\U_AHB/n93 ),
    .d(pnumcntF[0]),
    .e(pwm_state_read[0]),
    .o(_al_u3351_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*C)*~(D*B))"),
    .INIT(32'h020a22aa))
    _al_u3352 (
    .a(_al_u3351_o),
    .b(\U_AHB/n104_lutinv ),
    .c(\U_AHB/n102 ),
    .d(\U_AHB/h2h_hrdata [0]),
    .e(limit_r_pad[0]),
    .o(_al_u3352_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E)"),
    .INIT(32'h33533050))
    _al_u3353 (
    .a(_al_u3348_o),
    .b(_al_u3352_o),
    .c(_al_u3061_o),
    .d(\U_AHB/h2h_haddr [13]),
    .e(\U_AHB/h2h_hrdata [0]),
    .o(\U_AHB/n118 [0]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u336 (
    .a(\PWM4/pnumr [2]),
    .b(pnum4[2]),
    .c(pnum4[32]),
    .d(pwm_start_stop[20]),
    .o(\PWM4/n23 [2]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u337 (
    .a(\PWM4/pnumr [19]),
    .b(pnum4[19]),
    .c(pnum4[32]),
    .d(pwm_start_stop[20]),
    .o(\PWM4/n23 [19]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u338 (
    .a(\PWM4/pnumr [18]),
    .b(pnum4[18]),
    .c(pnum4[32]),
    .d(pwm_start_stop[20]),
    .o(\PWM4/n23 [18]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u339 (
    .a(\PWM4/pnumr [17]),
    .b(pnum4[17]),
    .c(pnum4[32]),
    .d(pwm_start_stop[20]),
    .o(\PWM4/n23 [17]));
  EF2_PHY_SPAD #(
    //.LOCATION("P22"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("16"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u34 (
    .do({open_n966,dir_pad[4]}),
    .ts(1'b1),
    .opad(dir[4]));  // CPLD_SOC_AHB_TOP.v(7)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u340 (
    .a(\PWM4/pnumr [16]),
    .b(pnum4[16]),
    .c(pnum4[32]),
    .d(pwm_start_stop[20]),
    .o(\PWM4/n23 [16]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u341 (
    .a(\PWM4/pnumr [15]),
    .b(pnum4[15]),
    .c(pnum4[32]),
    .d(pwm_start_stop[20]),
    .o(\PWM4/n23 [15]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u342 (
    .a(\PWM4/pnumr [14]),
    .b(pnum4[14]),
    .c(pnum4[32]),
    .d(pwm_start_stop[20]),
    .o(\PWM4/n23 [14]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u343 (
    .a(\PWM4/pnumr [13]),
    .b(pnum4[13]),
    .c(pnum4[32]),
    .d(pwm_start_stop[20]),
    .o(\PWM4/n23 [13]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u344 (
    .a(\PWM4/pnumr [12]),
    .b(pnum4[12]),
    .c(pnum4[32]),
    .d(pwm_start_stop[20]),
    .o(\PWM4/n23 [12]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u345 (
    .a(\PWM4/pnumr [11]),
    .b(pnum4[11]),
    .c(pnum4[32]),
    .d(pwm_start_stop[20]),
    .o(\PWM4/n23 [11]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u346 (
    .a(\PWM4/pnumr [10]),
    .b(pnum4[10]),
    .c(pnum4[32]),
    .d(pwm_start_stop[20]),
    .o(\PWM4/n23 [10]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u347 (
    .a(\PWM4/pnumr [1]),
    .b(pnum4[1]),
    .c(pnum4[32]),
    .d(pwm_start_stop[20]),
    .o(\PWM4/n23 [1]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u348 (
    .a(\PWM4/pnumr [0]),
    .b(pnum4[0]),
    .c(pnum4[32]),
    .d(pwm_start_stop[20]),
    .o(\PWM4/n23 [0]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u349 (
    .a(\PWM5/pnumr [9]),
    .b(pnum5[32]),
    .c(pnum5[9]),
    .d(pwm_start_stop[21]),
    .o(\PWM5/n23 [9]));
  EF2_PHY_PAD #(
    //.LOCATION("P132"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u35 (
    .do({open_n974,open_n975,open_n976,dir_pad[3]}),
    .opad(dir[3]));  // CPLD_SOC_AHB_TOP.v(7)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u350 (
    .a(\PWM5/pnumr [8]),
    .b(pnum5[32]),
    .c(pnum5[8]),
    .d(pwm_start_stop[21]),
    .o(\PWM5/n23 [8]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u351 (
    .a(\PWM5/pnumr [7]),
    .b(pnum5[32]),
    .c(pnum5[7]),
    .d(pwm_start_stop[21]),
    .o(\PWM5/n23 [7]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u352 (
    .a(\PWM5/pnumr [6]),
    .b(pnum5[32]),
    .c(pnum5[6]),
    .d(pwm_start_stop[21]),
    .o(\PWM5/n23 [6]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u353 (
    .a(\PWM5/pnumr [5]),
    .b(pnum5[32]),
    .c(pnum5[5]),
    .d(pwm_start_stop[21]),
    .o(\PWM5/n23 [5]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u354 (
    .a(\PWM5/pnumr [4]),
    .b(pnum5[32]),
    .c(pnum5[4]),
    .d(pwm_start_stop[21]),
    .o(\PWM5/n23 [4]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u355 (
    .a(\PWM5/pnumr [31]),
    .b(pnum5[31]),
    .c(pnum5[32]),
    .d(pwm_start_stop[21]),
    .o(\PWM5/n23 [31]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u356 (
    .a(\PWM5/pnumr [30]),
    .b(pnum5[30]),
    .c(pnum5[32]),
    .d(pwm_start_stop[21]),
    .o(\PWM5/n23 [30]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u357 (
    .a(\PWM5/pnumr [3]),
    .b(pnum5[3]),
    .c(pnum5[32]),
    .d(pwm_start_stop[21]),
    .o(\PWM5/n23 [3]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u358 (
    .a(\PWM5/pnumr [29]),
    .b(pnum5[29]),
    .c(pnum5[32]),
    .d(pwm_start_stop[21]),
    .o(\PWM5/n23 [29]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u359 (
    .a(\PWM5/pnumr [28]),
    .b(pnum5[28]),
    .c(pnum5[32]),
    .d(pwm_start_stop[21]),
    .o(\PWM5/n23 [28]));
  EF2_PHY_PAD #(
    //.LOCATION("P133"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u36 (
    .do({open_n997,open_n998,open_n999,dir_pad[2]}),
    .opad(dir[2]));  // CPLD_SOC_AHB_TOP.v(7)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u360 (
    .a(\PWM5/pnumr [27]),
    .b(pnum5[27]),
    .c(pnum5[32]),
    .d(pwm_start_stop[21]),
    .o(\PWM5/n23 [27]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u361 (
    .a(\PWM5/pnumr [26]),
    .b(pnum5[26]),
    .c(pnum5[32]),
    .d(pwm_start_stop[21]),
    .o(\PWM5/n23 [26]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u362 (
    .a(\PWM5/pnumr [25]),
    .b(pnum5[25]),
    .c(pnum5[32]),
    .d(pwm_start_stop[21]),
    .o(\PWM5/n23 [25]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u363 (
    .a(\PWM5/pnumr [24]),
    .b(pnum5[24]),
    .c(pnum5[32]),
    .d(pwm_start_stop[21]),
    .o(\PWM5/n23 [24]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u364 (
    .a(\PWM5/pnumr [23]),
    .b(pnum5[23]),
    .c(pnum5[32]),
    .d(pwm_start_stop[21]),
    .o(\PWM5/n23 [23]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u365 (
    .a(\PWM5/pnumr [22]),
    .b(pnum5[22]),
    .c(pnum5[32]),
    .d(pwm_start_stop[21]),
    .o(\PWM5/n23 [22]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u366 (
    .a(\PWM5/pnumr [21]),
    .b(pnum5[21]),
    .c(pnum5[32]),
    .d(pwm_start_stop[21]),
    .o(\PWM5/n23 [21]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u367 (
    .a(\PWM5/pnumr [20]),
    .b(pnum5[20]),
    .c(pnum5[32]),
    .d(pwm_start_stop[21]),
    .o(\PWM5/n23 [20]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u368 (
    .a(\PWM5/pnumr [2]),
    .b(pnum5[2]),
    .c(pnum5[32]),
    .d(pwm_start_stop[21]),
    .o(\PWM5/n23 [2]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u369 (
    .a(\PWM5/pnumr [19]),
    .b(pnum5[19]),
    .c(pnum5[32]),
    .d(pwm_start_stop[21]),
    .o(\PWM5/n23 [19]));
  EF2_PHY_SPAD #(
    //.LOCATION("P21"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("16"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u37 (
    .do({open_n1021,dir_pad[1]}),
    .ts(1'b1),
    .opad(dir[1]));  // CPLD_SOC_AHB_TOP.v(7)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u370 (
    .a(\PWM5/pnumr [18]),
    .b(pnum5[18]),
    .c(pnum5[32]),
    .d(pwm_start_stop[21]),
    .o(\PWM5/n23 [18]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u371 (
    .a(\PWM5/pnumr [17]),
    .b(pnum5[17]),
    .c(pnum5[32]),
    .d(pwm_start_stop[21]),
    .o(\PWM5/n23 [17]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u372 (
    .a(\PWM5/pnumr [16]),
    .b(pnum5[16]),
    .c(pnum5[32]),
    .d(pwm_start_stop[21]),
    .o(\PWM5/n23 [16]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u373 (
    .a(\PWM5/pnumr [15]),
    .b(pnum5[15]),
    .c(pnum5[32]),
    .d(pwm_start_stop[21]),
    .o(\PWM5/n23 [15]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u374 (
    .a(\PWM5/pnumr [14]),
    .b(pnum5[14]),
    .c(pnum5[32]),
    .d(pwm_start_stop[21]),
    .o(\PWM5/n23 [14]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u375 (
    .a(\PWM5/pnumr [13]),
    .b(pnum5[13]),
    .c(pnum5[32]),
    .d(pwm_start_stop[21]),
    .o(\PWM5/n23 [13]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u376 (
    .a(\PWM5/pnumr [12]),
    .b(pnum5[12]),
    .c(pnum5[32]),
    .d(pwm_start_stop[21]),
    .o(\PWM5/n23 [12]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u377 (
    .a(\PWM5/pnumr [11]),
    .b(pnum5[11]),
    .c(pnum5[32]),
    .d(pwm_start_stop[21]),
    .o(\PWM5/n23 [11]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u378 (
    .a(\PWM5/pnumr [10]),
    .b(pnum5[10]),
    .c(pnum5[32]),
    .d(pwm_start_stop[21]),
    .o(\PWM5/n23 [10]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u379 (
    .a(\PWM5/pnumr [1]),
    .b(pnum5[1]),
    .c(pnum5[32]),
    .d(pwm_start_stop[21]),
    .o(\PWM5/n23 [1]));
  EF2_PHY_PAD #(
    //.LOCATION("P138"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u38 (
    .do({open_n1029,open_n1030,open_n1031,dir_pad[0]}),
    .opad(dir[0]));  // CPLD_SOC_AHB_TOP.v(7)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u380 (
    .a(\PWM5/pnumr [0]),
    .b(pnum5[0]),
    .c(pnum5[32]),
    .d(pwm_start_stop[21]),
    .o(\PWM5/n23 [0]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u381 (
    .a(\PWM6/pnumr [9]),
    .b(pnum6[32]),
    .c(pnum6[9]),
    .d(pwm_start_stop[22]),
    .o(\PWM6/n23 [9]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u382 (
    .a(\PWM6/pnumr [8]),
    .b(pnum6[32]),
    .c(pnum6[8]),
    .d(pwm_start_stop[22]),
    .o(\PWM6/n23 [8]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u383 (
    .a(\PWM6/pnumr [7]),
    .b(pnum6[32]),
    .c(pnum6[7]),
    .d(pwm_start_stop[22]),
    .o(\PWM6/n23 [7]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u384 (
    .a(\PWM6/pnumr [6]),
    .b(pnum6[32]),
    .c(pnum6[6]),
    .d(pwm_start_stop[22]),
    .o(\PWM6/n23 [6]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u385 (
    .a(\PWM6/pnumr [5]),
    .b(pnum6[32]),
    .c(pnum6[5]),
    .d(pwm_start_stop[22]),
    .o(\PWM6/n23 [5]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u386 (
    .a(\PWM6/pnumr [4]),
    .b(pnum6[32]),
    .c(pnum6[4]),
    .d(pwm_start_stop[22]),
    .o(\PWM6/n23 [4]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u387 (
    .a(\PWM6/pnumr [31]),
    .b(pnum6[31]),
    .c(pnum6[32]),
    .d(pwm_start_stop[22]),
    .o(\PWM6/n23 [31]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u388 (
    .a(\PWM6/pnumr [30]),
    .b(pnum6[30]),
    .c(pnum6[32]),
    .d(pwm_start_stop[22]),
    .o(\PWM6/n23 [30]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u389 (
    .a(\PWM6/pnumr [3]),
    .b(pnum6[3]),
    .c(pnum6[32]),
    .d(pwm_start_stop[22]),
    .o(\PWM6/n23 [3]));
  EF2_PHY_SPAD #(
    //.LOCATION("p10"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u39 (
    .do({open_n1053,gpio_out_pad[31]}),
    .ts(1'b1),
    .opad(gpio_out[31]));  // CPLD_SOC_AHB_TOP.v(8)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u390 (
    .a(\PWM6/pnumr [29]),
    .b(pnum6[29]),
    .c(pnum6[32]),
    .d(pwm_start_stop[22]),
    .o(\PWM6/n23 [29]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u391 (
    .a(\PWM6/pnumr [28]),
    .b(pnum6[28]),
    .c(pnum6[32]),
    .d(pwm_start_stop[22]),
    .o(\PWM6/n23 [28]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u392 (
    .a(\PWM6/pnumr [27]),
    .b(pnum6[27]),
    .c(pnum6[32]),
    .d(pwm_start_stop[22]),
    .o(\PWM6/n23 [27]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u393 (
    .a(\PWM6/pnumr [26]),
    .b(pnum6[26]),
    .c(pnum6[32]),
    .d(pwm_start_stop[22]),
    .o(\PWM6/n23 [26]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u394 (
    .a(\PWM6/pnumr [25]),
    .b(pnum6[25]),
    .c(pnum6[32]),
    .d(pwm_start_stop[22]),
    .o(\PWM6/n23 [25]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u395 (
    .a(\PWM6/pnumr [24]),
    .b(pnum6[24]),
    .c(pnum6[32]),
    .d(pwm_start_stop[22]),
    .o(\PWM6/n23 [24]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u396 (
    .a(\PWM6/pnumr [23]),
    .b(pnum6[23]),
    .c(pnum6[32]),
    .d(pwm_start_stop[22]),
    .o(\PWM6/n23 [23]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u397 (
    .a(\PWM6/pnumr [22]),
    .b(pnum6[22]),
    .c(pnum6[32]),
    .d(pwm_start_stop[22]),
    .o(\PWM6/n23 [22]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u398 (
    .a(\PWM6/pnumr [21]),
    .b(pnum6[21]),
    .c(pnum6[32]),
    .d(pwm_start_stop[22]),
    .o(\PWM6/n23 [21]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u399 (
    .a(\PWM6/pnumr [20]),
    .b(pnum6[20]),
    .c(pnum6[32]),
    .d(pwm_start_stop[22]),
    .o(\PWM6/n23 [20]));
  EF2_PHY_PAD #(
    //.LOCATION("p120"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u40 (
    .do({open_n1061,open_n1062,open_n1063,gpio_out_pad[30]}),
    .opad(gpio_out[30]));  // CPLD_SOC_AHB_TOP.v(8)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u400 (
    .a(\PWM6/pnumr [2]),
    .b(pnum6[2]),
    .c(pnum6[32]),
    .d(pwm_start_stop[22]),
    .o(\PWM6/n23 [2]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u401 (
    .a(\PWM6/pnumr [19]),
    .b(pnum6[19]),
    .c(pnum6[32]),
    .d(pwm_start_stop[22]),
    .o(\PWM6/n23 [19]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u402 (
    .a(\PWM6/pnumr [18]),
    .b(pnum6[18]),
    .c(pnum6[32]),
    .d(pwm_start_stop[22]),
    .o(\PWM6/n23 [18]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u403 (
    .a(\PWM6/pnumr [17]),
    .b(pnum6[17]),
    .c(pnum6[32]),
    .d(pwm_start_stop[22]),
    .o(\PWM6/n23 [17]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u404 (
    .a(\PWM6/pnumr [16]),
    .b(pnum6[16]),
    .c(pnum6[32]),
    .d(pwm_start_stop[22]),
    .o(\PWM6/n23 [16]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u405 (
    .a(\PWM6/pnumr [15]),
    .b(pnum6[15]),
    .c(pnum6[32]),
    .d(pwm_start_stop[22]),
    .o(\PWM6/n23 [15]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u406 (
    .a(\PWM6/pnumr [14]),
    .b(pnum6[14]),
    .c(pnum6[32]),
    .d(pwm_start_stop[22]),
    .o(\PWM6/n23 [14]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u407 (
    .a(\PWM6/pnumr [13]),
    .b(pnum6[13]),
    .c(pnum6[32]),
    .d(pwm_start_stop[22]),
    .o(\PWM6/n23 [13]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u408 (
    .a(\PWM6/pnumr [12]),
    .b(pnum6[12]),
    .c(pnum6[32]),
    .d(pwm_start_stop[22]),
    .o(\PWM6/n23 [12]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u409 (
    .a(\PWM6/pnumr [11]),
    .b(pnum6[11]),
    .c(pnum6[32]),
    .d(pwm_start_stop[22]),
    .o(\PWM6/n23 [11]));
  EF2_PHY_SPAD #(
    //.LOCATION("p19"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u41 (
    .do({open_n1085,gpio_out_pad[29]}),
    .ts(1'b1),
    .opad(gpio_out[29]));  // CPLD_SOC_AHB_TOP.v(8)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u410 (
    .a(\PWM6/pnumr [10]),
    .b(pnum6[10]),
    .c(pnum6[32]),
    .d(pwm_start_stop[22]),
    .o(\PWM6/n23 [10]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u411 (
    .a(\PWM6/pnumr [1]),
    .b(pnum6[1]),
    .c(pnum6[32]),
    .d(pwm_start_stop[22]),
    .o(\PWM6/n23 [1]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u412 (
    .a(\PWM6/pnumr [0]),
    .b(pnum6[0]),
    .c(pnum6[32]),
    .d(pwm_start_stop[22]),
    .o(\PWM6/n23 [0]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u413 (
    .a(\PWM7/pnumr [9]),
    .b(pnum7[32]),
    .c(pnum7[9]),
    .d(pwm_start_stop[23]),
    .o(\PWM7/n23 [9]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u414 (
    .a(\PWM7/pnumr [8]),
    .b(pnum7[32]),
    .c(pnum7[8]),
    .d(pwm_start_stop[23]),
    .o(\PWM7/n23 [8]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u415 (
    .a(\PWM7/pnumr [7]),
    .b(pnum7[32]),
    .c(pnum7[7]),
    .d(pwm_start_stop[23]),
    .o(\PWM7/n23 [7]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u416 (
    .a(\PWM7/pnumr [6]),
    .b(pnum7[32]),
    .c(pnum7[6]),
    .d(pwm_start_stop[23]),
    .o(\PWM7/n23 [6]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u417 (
    .a(\PWM7/pnumr [5]),
    .b(pnum7[32]),
    .c(pnum7[5]),
    .d(pwm_start_stop[23]),
    .o(\PWM7/n23 [5]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u418 (
    .a(\PWM7/pnumr [4]),
    .b(pnum7[32]),
    .c(pnum7[4]),
    .d(pwm_start_stop[23]),
    .o(\PWM7/n23 [4]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u419 (
    .a(\PWM7/pnumr [31]),
    .b(pnum7[31]),
    .c(pnum7[32]),
    .d(pwm_start_stop[23]),
    .o(\PWM7/n23 [31]));
  EF2_PHY_PAD #(
    //.LOCATION("p61"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u42 (
    .do({open_n1093,open_n1094,open_n1095,gpio_out_pad[28]}),
    .opad(gpio_out[28]));  // CPLD_SOC_AHB_TOP.v(8)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u420 (
    .a(\PWM7/pnumr [30]),
    .b(pnum7[30]),
    .c(pnum7[32]),
    .d(pwm_start_stop[23]),
    .o(\PWM7/n23 [30]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u421 (
    .a(\PWM7/pnumr [3]),
    .b(pnum7[3]),
    .c(pnum7[32]),
    .d(pwm_start_stop[23]),
    .o(\PWM7/n23 [3]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u422 (
    .a(\PWM7/pnumr [29]),
    .b(pnum7[29]),
    .c(pnum7[32]),
    .d(pwm_start_stop[23]),
    .o(\PWM7/n23 [29]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u423 (
    .a(\PWM7/pnumr [28]),
    .b(pnum7[28]),
    .c(pnum7[32]),
    .d(pwm_start_stop[23]),
    .o(\PWM7/n23 [28]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u424 (
    .a(\PWM7/pnumr [27]),
    .b(pnum7[27]),
    .c(pnum7[32]),
    .d(pwm_start_stop[23]),
    .o(\PWM7/n23 [27]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u425 (
    .a(\PWM7/pnumr [26]),
    .b(pnum7[26]),
    .c(pnum7[32]),
    .d(pwm_start_stop[23]),
    .o(\PWM7/n23 [26]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u426 (
    .a(\PWM7/pnumr [25]),
    .b(pnum7[25]),
    .c(pnum7[32]),
    .d(pwm_start_stop[23]),
    .o(\PWM7/n23 [25]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u427 (
    .a(\PWM7/pnumr [24]),
    .b(pnum7[24]),
    .c(pnum7[32]),
    .d(pwm_start_stop[23]),
    .o(\PWM7/n23 [24]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u428 (
    .a(\PWM7/pnumr [23]),
    .b(pnum7[23]),
    .c(pnum7[32]),
    .d(pwm_start_stop[23]),
    .o(\PWM7/n23 [23]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u429 (
    .a(\PWM7/pnumr [22]),
    .b(pnum7[22]),
    .c(pnum7[32]),
    .d(pwm_start_stop[23]),
    .o(\PWM7/n23 [22]));
  EF2_PHY_PAD #(
    //.LOCATION("p62"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u43 (
    .do({open_n1116,open_n1117,open_n1118,gpio_out_pad[27]}),
    .opad(gpio_out[27]));  // CPLD_SOC_AHB_TOP.v(8)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u430 (
    .a(\PWM7/pnumr [21]),
    .b(pnum7[21]),
    .c(pnum7[32]),
    .d(pwm_start_stop[23]),
    .o(\PWM7/n23 [21]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u431 (
    .a(\PWM7/pnumr [20]),
    .b(pnum7[20]),
    .c(pnum7[32]),
    .d(pwm_start_stop[23]),
    .o(\PWM7/n23 [20]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u432 (
    .a(\PWM7/pnumr [2]),
    .b(pnum7[2]),
    .c(pnum7[32]),
    .d(pwm_start_stop[23]),
    .o(\PWM7/n23 [2]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u433 (
    .a(\PWM7/pnumr [19]),
    .b(pnum7[19]),
    .c(pnum7[32]),
    .d(pwm_start_stop[23]),
    .o(\PWM7/n23 [19]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u434 (
    .a(\PWM7/pnumr [18]),
    .b(pnum7[18]),
    .c(pnum7[32]),
    .d(pwm_start_stop[23]),
    .o(\PWM7/n23 [18]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u435 (
    .a(\PWM7/pnumr [17]),
    .b(pnum7[17]),
    .c(pnum7[32]),
    .d(pwm_start_stop[23]),
    .o(\PWM7/n23 [17]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u436 (
    .a(\PWM7/pnumr [16]),
    .b(pnum7[16]),
    .c(pnum7[32]),
    .d(pwm_start_stop[23]),
    .o(\PWM7/n23 [16]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u437 (
    .a(\PWM7/pnumr [15]),
    .b(pnum7[15]),
    .c(pnum7[32]),
    .d(pwm_start_stop[23]),
    .o(\PWM7/n23 [15]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u438 (
    .a(\PWM7/pnumr [14]),
    .b(pnum7[14]),
    .c(pnum7[32]),
    .d(pwm_start_stop[23]),
    .o(\PWM7/n23 [14]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u439 (
    .a(\PWM7/pnumr [13]),
    .b(pnum7[13]),
    .c(pnum7[32]),
    .d(pwm_start_stop[23]),
    .o(\PWM7/n23 [13]));
  EF2_PHY_SPAD #(
    //.LOCATION("p91"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u44 (
    .do({open_n1140,gpio_out_pad[26]}),
    .ts(1'b1),
    .opad(gpio_out[26]));  // CPLD_SOC_AHB_TOP.v(8)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u440 (
    .a(\PWM7/pnumr [12]),
    .b(pnum7[12]),
    .c(pnum7[32]),
    .d(pwm_start_stop[23]),
    .o(\PWM7/n23 [12]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u441 (
    .a(\PWM7/pnumr [11]),
    .b(pnum7[11]),
    .c(pnum7[32]),
    .d(pwm_start_stop[23]),
    .o(\PWM7/n23 [11]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u442 (
    .a(\PWM7/pnumr [10]),
    .b(pnum7[10]),
    .c(pnum7[32]),
    .d(pwm_start_stop[23]),
    .o(\PWM7/n23 [10]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u443 (
    .a(\PWM7/pnumr [1]),
    .b(pnum7[1]),
    .c(pnum7[32]),
    .d(pwm_start_stop[23]),
    .o(\PWM7/n23 [1]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u444 (
    .a(\PWM7/pnumr [0]),
    .b(pnum7[0]),
    .c(pnum7[32]),
    .d(pwm_start_stop[23]),
    .o(\PWM7/n23 [0]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u445 (
    .a(\PWM8/pnumr [9]),
    .b(pnum8[32]),
    .c(pnum8[9]),
    .d(pwm_start_stop[24]),
    .o(\PWM8/n23 [9]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u446 (
    .a(\PWM8/pnumr [8]),
    .b(pnum8[32]),
    .c(pnum8[8]),
    .d(pwm_start_stop[24]),
    .o(\PWM8/n23 [8]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u447 (
    .a(\PWM8/pnumr [7]),
    .b(pnum8[32]),
    .c(pnum8[7]),
    .d(pwm_start_stop[24]),
    .o(\PWM8/n23 [7]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u448 (
    .a(\PWM8/pnumr [6]),
    .b(pnum8[32]),
    .c(pnum8[6]),
    .d(pwm_start_stop[24]),
    .o(\PWM8/n23 [6]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u449 (
    .a(\PWM8/pnumr [5]),
    .b(pnum8[32]),
    .c(pnum8[5]),
    .d(pwm_start_stop[24]),
    .o(\PWM8/n23 [5]));
  EF2_PHY_PAD #(
    //.LOCATION("p109"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u45 (
    .do({open_n1148,open_n1149,open_n1150,gpio_out_pad[25]}),
    .opad(gpio_out[25]));  // CPLD_SOC_AHB_TOP.v(8)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u450 (
    .a(\PWM8/pnumr [4]),
    .b(pnum8[32]),
    .c(pnum8[4]),
    .d(pwm_start_stop[24]),
    .o(\PWM8/n23 [4]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u451 (
    .a(\PWM8/pnumr [31]),
    .b(pnum8[31]),
    .c(pnum8[32]),
    .d(pwm_start_stop[24]),
    .o(\PWM8/n23 [31]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u452 (
    .a(\PWM8/pnumr [30]),
    .b(pnum8[30]),
    .c(pnum8[32]),
    .d(pwm_start_stop[24]),
    .o(\PWM8/n23 [30]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u453 (
    .a(\PWM8/pnumr [3]),
    .b(pnum8[3]),
    .c(pnum8[32]),
    .d(pwm_start_stop[24]),
    .o(\PWM8/n23 [3]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u454 (
    .a(\PWM8/pnumr [29]),
    .b(pnum8[29]),
    .c(pnum8[32]),
    .d(pwm_start_stop[24]),
    .o(\PWM8/n23 [29]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u455 (
    .a(\PWM8/pnumr [28]),
    .b(pnum8[28]),
    .c(pnum8[32]),
    .d(pwm_start_stop[24]),
    .o(\PWM8/n23 [28]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u456 (
    .a(\PWM8/pnumr [27]),
    .b(pnum8[27]),
    .c(pnum8[32]),
    .d(pwm_start_stop[24]),
    .o(\PWM8/n23 [27]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u457 (
    .a(\PWM8/pnumr [26]),
    .b(pnum8[26]),
    .c(pnum8[32]),
    .d(pwm_start_stop[24]),
    .o(\PWM8/n23 [26]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u458 (
    .a(\PWM8/pnumr [25]),
    .b(pnum8[25]),
    .c(pnum8[32]),
    .d(pwm_start_stop[24]),
    .o(\PWM8/n23 [25]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u459 (
    .a(\PWM8/pnumr [24]),
    .b(pnum8[24]),
    .c(pnum8[32]),
    .d(pwm_start_stop[24]),
    .o(\PWM8/n23 [24]));
  EF2_PHY_PAD #(
    //.LOCATION("p143"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u46 (
    .do({open_n1171,open_n1172,open_n1173,gpio_out_pad[24]}),
    .opad(gpio_out[24]));  // CPLD_SOC_AHB_TOP.v(8)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u460 (
    .a(\PWM8/pnumr [23]),
    .b(pnum8[23]),
    .c(pnum8[32]),
    .d(pwm_start_stop[24]),
    .o(\PWM8/n23 [23]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u461 (
    .a(\PWM8/pnumr [22]),
    .b(pnum8[22]),
    .c(pnum8[32]),
    .d(pwm_start_stop[24]),
    .o(\PWM8/n23 [22]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u462 (
    .a(\PWM8/pnumr [21]),
    .b(pnum8[21]),
    .c(pnum8[32]),
    .d(pwm_start_stop[24]),
    .o(\PWM8/n23 [21]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u463 (
    .a(\PWM8/pnumr [20]),
    .b(pnum8[20]),
    .c(pnum8[32]),
    .d(pwm_start_stop[24]),
    .o(\PWM8/n23 [20]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u464 (
    .a(\PWM8/pnumr [2]),
    .b(pnum8[2]),
    .c(pnum8[32]),
    .d(pwm_start_stop[24]),
    .o(\PWM8/n23 [2]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u465 (
    .a(\PWM8/pnumr [19]),
    .b(pnum8[19]),
    .c(pnum8[32]),
    .d(pwm_start_stop[24]),
    .o(\PWM8/n23 [19]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u466 (
    .a(\PWM8/pnumr [18]),
    .b(pnum8[18]),
    .c(pnum8[32]),
    .d(pwm_start_stop[24]),
    .o(\PWM8/n23 [18]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u467 (
    .a(\PWM8/pnumr [17]),
    .b(pnum8[17]),
    .c(pnum8[32]),
    .d(pwm_start_stop[24]),
    .o(\PWM8/n23 [17]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u468 (
    .a(\PWM8/pnumr [16]),
    .b(pnum8[16]),
    .c(pnum8[32]),
    .d(pwm_start_stop[24]),
    .o(\PWM8/n23 [16]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u469 (
    .a(\PWM8/pnumr [15]),
    .b(pnum8[15]),
    .c(pnum8[32]),
    .d(pwm_start_stop[24]),
    .o(\PWM8/n23 [15]));
  EF2_PHY_PAD #(
    //.LOCATION("p71"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u47 (
    .do({open_n1194,open_n1195,open_n1196,gpio_out_pad[23]}),
    .opad(gpio_out[23]));  // CPLD_SOC_AHB_TOP.v(8)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u470 (
    .a(\PWM8/pnumr [14]),
    .b(pnum8[14]),
    .c(pnum8[32]),
    .d(pwm_start_stop[24]),
    .o(\PWM8/n23 [14]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u471 (
    .a(\PWM8/pnumr [13]),
    .b(pnum8[13]),
    .c(pnum8[32]),
    .d(pwm_start_stop[24]),
    .o(\PWM8/n23 [13]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u472 (
    .a(\PWM8/pnumr [12]),
    .b(pnum8[12]),
    .c(pnum8[32]),
    .d(pwm_start_stop[24]),
    .o(\PWM8/n23 [12]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u473 (
    .a(\PWM8/pnumr [11]),
    .b(pnum8[11]),
    .c(pnum8[32]),
    .d(pwm_start_stop[24]),
    .o(\PWM8/n23 [11]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u474 (
    .a(\PWM8/pnumr [10]),
    .b(pnum8[10]),
    .c(pnum8[32]),
    .d(pwm_start_stop[24]),
    .o(\PWM8/n23 [10]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u475 (
    .a(\PWM8/pnumr [1]),
    .b(pnum8[1]),
    .c(pnum8[32]),
    .d(pwm_start_stop[24]),
    .o(\PWM8/n23 [1]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u476 (
    .a(\PWM8/pnumr [0]),
    .b(pnum8[0]),
    .c(pnum8[32]),
    .d(pwm_start_stop[24]),
    .o(\PWM8/n23 [0]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u477 (
    .a(\PWM9/pnumr [9]),
    .b(pnum9[32]),
    .c(pnum9[9]),
    .d(pwm_start_stop[25]),
    .o(\PWM9/n23 [9]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u478 (
    .a(\PWM9/pnumr [8]),
    .b(pnum9[32]),
    .c(pnum9[8]),
    .d(pwm_start_stop[25]),
    .o(\PWM9/n23 [8]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u479 (
    .a(\PWM9/pnumr [7]),
    .b(pnum9[32]),
    .c(pnum9[7]),
    .d(pwm_start_stop[25]),
    .o(\PWM9/n23 [7]));
  EF2_PHY_SPAD #(
    //.LOCATION("p73"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u48 (
    .do({open_n1218,gpio_out_pad[22]}),
    .ts(1'b1),
    .opad(gpio_out[22]));  // CPLD_SOC_AHB_TOP.v(8)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u480 (
    .a(\PWM9/pnumr [6]),
    .b(pnum9[32]),
    .c(pnum9[6]),
    .d(pwm_start_stop[25]),
    .o(\PWM9/n23 [6]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u481 (
    .a(\PWM9/pnumr [5]),
    .b(pnum9[32]),
    .c(pnum9[5]),
    .d(pwm_start_stop[25]),
    .o(\PWM9/n23 [5]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u482 (
    .a(\PWM9/pnumr [4]),
    .b(pnum9[32]),
    .c(pnum9[4]),
    .d(pwm_start_stop[25]),
    .o(\PWM9/n23 [4]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u483 (
    .a(\PWM9/pnumr [31]),
    .b(pnum9[31]),
    .c(pnum9[32]),
    .d(pwm_start_stop[25]),
    .o(\PWM9/n23 [31]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u484 (
    .a(\PWM9/pnumr [30]),
    .b(pnum9[30]),
    .c(pnum9[32]),
    .d(pwm_start_stop[25]),
    .o(\PWM9/n23 [30]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u485 (
    .a(\PWM9/pnumr [3]),
    .b(pnum9[3]),
    .c(pnum9[32]),
    .d(pwm_start_stop[25]),
    .o(\PWM9/n23 [3]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u486 (
    .a(\PWM9/pnumr [29]),
    .b(pnum9[29]),
    .c(pnum9[32]),
    .d(pwm_start_stop[25]),
    .o(\PWM9/n23 [29]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u487 (
    .a(\PWM9/pnumr [28]),
    .b(pnum9[28]),
    .c(pnum9[32]),
    .d(pwm_start_stop[25]),
    .o(\PWM9/n23 [28]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u488 (
    .a(\PWM9/pnumr [27]),
    .b(pnum9[27]),
    .c(pnum9[32]),
    .d(pwm_start_stop[25]),
    .o(\PWM9/n23 [27]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u489 (
    .a(\PWM9/pnumr [26]),
    .b(pnum9[26]),
    .c(pnum9[32]),
    .d(pwm_start_stop[25]),
    .o(\PWM9/n23 [26]));
  EF2_PHY_SPAD #(
    //.LOCATION("p11"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u49 (
    .do({open_n1227,gpio_out_pad[21]}),
    .ts(1'b1),
    .opad(gpio_out[21]));  // CPLD_SOC_AHB_TOP.v(8)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u490 (
    .a(\PWM9/pnumr [25]),
    .b(pnum9[25]),
    .c(pnum9[32]),
    .d(pwm_start_stop[25]),
    .o(\PWM9/n23 [25]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u491 (
    .a(\PWM9/pnumr [24]),
    .b(pnum9[24]),
    .c(pnum9[32]),
    .d(pwm_start_stop[25]),
    .o(\PWM9/n23 [24]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u492 (
    .a(\PWM9/pnumr [23]),
    .b(pnum9[23]),
    .c(pnum9[32]),
    .d(pwm_start_stop[25]),
    .o(\PWM9/n23 [23]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u493 (
    .a(\PWM9/pnumr [22]),
    .b(pnum9[22]),
    .c(pnum9[32]),
    .d(pwm_start_stop[25]),
    .o(\PWM9/n23 [22]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u494 (
    .a(\PWM9/pnumr [21]),
    .b(pnum9[21]),
    .c(pnum9[32]),
    .d(pwm_start_stop[25]),
    .o(\PWM9/n23 [21]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u495 (
    .a(\PWM9/pnumr [20]),
    .b(pnum9[20]),
    .c(pnum9[32]),
    .d(pwm_start_stop[25]),
    .o(\PWM9/n23 [20]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u496 (
    .a(\PWM9/pnumr [2]),
    .b(pnum9[2]),
    .c(pnum9[32]),
    .d(pwm_start_stop[25]),
    .o(\PWM9/n23 [2]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u497 (
    .a(\PWM9/pnumr [19]),
    .b(pnum9[19]),
    .c(pnum9[32]),
    .d(pwm_start_stop[25]),
    .o(\PWM9/n23 [19]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u498 (
    .a(\PWM9/pnumr [18]),
    .b(pnum9[18]),
    .c(pnum9[32]),
    .d(pwm_start_stop[25]),
    .o(\PWM9/n23 [18]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u499 (
    .a(\PWM9/pnumr [17]),
    .b(pnum9[17]),
    .c(pnum9[32]),
    .d(pwm_start_stop[25]),
    .o(\PWM9/n23 [17]));
  EF2_PHY_SPAD #(
    //.LOCATION("p13"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u50 (
    .do({open_n1236,gpio_out_pad[20]}),
    .ts(1'b1),
    .opad(gpio_out[20]));  // CPLD_SOC_AHB_TOP.v(8)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u500 (
    .a(\PWM9/pnumr [16]),
    .b(pnum9[16]),
    .c(pnum9[32]),
    .d(pwm_start_stop[25]),
    .o(\PWM9/n23 [16]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u501 (
    .a(\PWM9/pnumr [15]),
    .b(pnum9[15]),
    .c(pnum9[32]),
    .d(pwm_start_stop[25]),
    .o(\PWM9/n23 [15]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u502 (
    .a(\PWM9/pnumr [14]),
    .b(pnum9[14]),
    .c(pnum9[32]),
    .d(pwm_start_stop[25]),
    .o(\PWM9/n23 [14]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u503 (
    .a(\PWM9/pnumr [13]),
    .b(pnum9[13]),
    .c(pnum9[32]),
    .d(pwm_start_stop[25]),
    .o(\PWM9/n23 [13]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u504 (
    .a(\PWM9/pnumr [12]),
    .b(pnum9[12]),
    .c(pnum9[32]),
    .d(pwm_start_stop[25]),
    .o(\PWM9/n23 [12]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u505 (
    .a(\PWM9/pnumr [11]),
    .b(pnum9[11]),
    .c(pnum9[32]),
    .d(pwm_start_stop[25]),
    .o(\PWM9/n23 [11]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u506 (
    .a(\PWM9/pnumr [10]),
    .b(pnum9[10]),
    .c(pnum9[32]),
    .d(pwm_start_stop[25]),
    .o(\PWM9/n23 [10]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u507 (
    .a(\PWM9/pnumr [1]),
    .b(pnum9[1]),
    .c(pnum9[32]),
    .d(pwm_start_stop[25]),
    .o(\PWM9/n23 [1]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u508 (
    .a(\PWM9/pnumr [0]),
    .b(pnum9[0]),
    .c(pnum9[32]),
    .d(pwm_start_stop[25]),
    .o(\PWM9/n23 [0]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u509 (
    .a(\PWMA/pnumr [9]),
    .b(pnumA[32]),
    .c(pnumA[9]),
    .d(pwm_start_stop[26]),
    .o(\PWMA/n23 [9]));
  EF2_PHY_PAD #(
    //.LOCATION("p39"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u51 (
    .do({open_n1244,open_n1245,open_n1246,gpio_out_pad[19]}),
    .opad(gpio_out[19]));  // CPLD_SOC_AHB_TOP.v(8)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u510 (
    .a(\PWMA/pnumr [8]),
    .b(pnumA[32]),
    .c(pnumA[8]),
    .d(pwm_start_stop[26]),
    .o(\PWMA/n23 [8]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u511 (
    .a(\PWMA/pnumr [7]),
    .b(pnumA[32]),
    .c(pnumA[7]),
    .d(pwm_start_stop[26]),
    .o(\PWMA/n23 [7]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u512 (
    .a(\PWMA/pnumr [6]),
    .b(pnumA[32]),
    .c(pnumA[6]),
    .d(pwm_start_stop[26]),
    .o(\PWMA/n23 [6]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u513 (
    .a(\PWMA/pnumr [5]),
    .b(pnumA[32]),
    .c(pnumA[5]),
    .d(pwm_start_stop[26]),
    .o(\PWMA/n23 [5]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u514 (
    .a(\PWMA/pnumr [4]),
    .b(pnumA[32]),
    .c(pnumA[4]),
    .d(pwm_start_stop[26]),
    .o(\PWMA/n23 [4]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u515 (
    .a(\PWMA/pnumr [31]),
    .b(pnumA[31]),
    .c(pnumA[32]),
    .d(pwm_start_stop[26]),
    .o(\PWMA/n23 [31]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u516 (
    .a(\PWMA/pnumr [30]),
    .b(pnumA[30]),
    .c(pnumA[32]),
    .d(pwm_start_stop[26]),
    .o(\PWMA/n23 [30]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u517 (
    .a(\PWMA/pnumr [3]),
    .b(pnumA[3]),
    .c(pnumA[32]),
    .d(pwm_start_stop[26]),
    .o(\PWMA/n23 [3]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u518 (
    .a(\PWMA/pnumr [29]),
    .b(pnumA[29]),
    .c(pnumA[32]),
    .d(pwm_start_stop[26]),
    .o(\PWMA/n23 [29]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u519 (
    .a(\PWMA/pnumr [28]),
    .b(pnumA[28]),
    .c(pnumA[32]),
    .d(pwm_start_stop[26]),
    .o(\PWMA/n23 [28]));
  EF2_PHY_SPAD #(
    //.LOCATION("p74"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u52 (
    .do({open_n1268,gpio_out_pad[18]}),
    .ts(1'b1),
    .opad(gpio_out[18]));  // CPLD_SOC_AHB_TOP.v(8)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u520 (
    .a(\PWMA/pnumr [27]),
    .b(pnumA[27]),
    .c(pnumA[32]),
    .d(pwm_start_stop[26]),
    .o(\PWMA/n23 [27]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u521 (
    .a(\PWMA/pnumr [26]),
    .b(pnumA[26]),
    .c(pnumA[32]),
    .d(pwm_start_stop[26]),
    .o(\PWMA/n23 [26]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u522 (
    .a(\PWMA/pnumr [25]),
    .b(pnumA[25]),
    .c(pnumA[32]),
    .d(pwm_start_stop[26]),
    .o(\PWMA/n23 [25]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u523 (
    .a(\PWMA/pnumr [24]),
    .b(pnumA[24]),
    .c(pnumA[32]),
    .d(pwm_start_stop[26]),
    .o(\PWMA/n23 [24]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u524 (
    .a(\PWMA/pnumr [23]),
    .b(pnumA[23]),
    .c(pnumA[32]),
    .d(pwm_start_stop[26]),
    .o(\PWMA/n23 [23]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u525 (
    .a(\PWMA/pnumr [22]),
    .b(pnumA[22]),
    .c(pnumA[32]),
    .d(pwm_start_stop[26]),
    .o(\PWMA/n23 [22]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u526 (
    .a(\PWMA/pnumr [21]),
    .b(pnumA[21]),
    .c(pnumA[32]),
    .d(pwm_start_stop[26]),
    .o(\PWMA/n23 [21]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u527 (
    .a(\PWMA/pnumr [20]),
    .b(pnumA[20]),
    .c(pnumA[32]),
    .d(pwm_start_stop[26]),
    .o(\PWMA/n23 [20]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u528 (
    .a(\PWMA/pnumr [2]),
    .b(pnumA[2]),
    .c(pnumA[32]),
    .d(pwm_start_stop[26]),
    .o(\PWMA/n23 [2]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u529 (
    .a(\PWMA/pnumr [19]),
    .b(pnumA[19]),
    .c(pnumA[32]),
    .d(pwm_start_stop[26]),
    .o(\PWMA/n23 [19]));
  EF2_PHY_PAD #(
    //.LOCATION("p110"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u53 (
    .do({open_n1276,open_n1277,open_n1278,gpio_out_pad[17]}),
    .opad(gpio_out[17]));  // CPLD_SOC_AHB_TOP.v(8)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u530 (
    .a(\PWMA/pnumr [18]),
    .b(pnumA[18]),
    .c(pnumA[32]),
    .d(pwm_start_stop[26]),
    .o(\PWMA/n23 [18]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u531 (
    .a(\PWMA/pnumr [17]),
    .b(pnumA[17]),
    .c(pnumA[32]),
    .d(pwm_start_stop[26]),
    .o(\PWMA/n23 [17]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u532 (
    .a(\PWMA/pnumr [16]),
    .b(pnumA[16]),
    .c(pnumA[32]),
    .d(pwm_start_stop[26]),
    .o(\PWMA/n23 [16]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u533 (
    .a(\PWMA/pnumr [15]),
    .b(pnumA[15]),
    .c(pnumA[32]),
    .d(pwm_start_stop[26]),
    .o(\PWMA/n23 [15]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u534 (
    .a(\PWMA/pnumr [14]),
    .b(pnumA[14]),
    .c(pnumA[32]),
    .d(pwm_start_stop[26]),
    .o(\PWMA/n23 [14]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u535 (
    .a(\PWMA/pnumr [13]),
    .b(pnumA[13]),
    .c(pnumA[32]),
    .d(pwm_start_stop[26]),
    .o(\PWMA/n23 [13]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u536 (
    .a(\PWMA/pnumr [12]),
    .b(pnumA[12]),
    .c(pnumA[32]),
    .d(pwm_start_stop[26]),
    .o(\PWMA/n23 [12]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u537 (
    .a(\PWMA/pnumr [11]),
    .b(pnumA[11]),
    .c(pnumA[32]),
    .d(pwm_start_stop[26]),
    .o(\PWMA/n23 [11]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u538 (
    .a(\PWMA/pnumr [10]),
    .b(pnumA[10]),
    .c(pnumA[32]),
    .d(pwm_start_stop[26]),
    .o(\PWMA/n23 [10]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u539 (
    .a(\PWMA/pnumr [1]),
    .b(pnumA[1]),
    .c(pnumA[32]),
    .d(pwm_start_stop[26]),
    .o(\PWMA/n23 [1]));
  EF2_PHY_PAD #(
    //.LOCATION("p140"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u54 (
    .do({open_n1299,open_n1300,open_n1301,gpio_out_pad[16]}),
    .opad(gpio_out[16]));  // CPLD_SOC_AHB_TOP.v(8)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u540 (
    .a(\PWMA/pnumr [0]),
    .b(pnumA[0]),
    .c(pnumA[32]),
    .d(pwm_start_stop[26]),
    .o(\PWMA/n23 [0]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u541 (
    .a(\PWMB/pnumr [9]),
    .b(pnumB[32]),
    .c(pnumB[9]),
    .d(pwm_start_stop[27]),
    .o(\PWMB/n23 [9]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u542 (
    .a(\PWMB/pnumr [8]),
    .b(pnumB[32]),
    .c(pnumB[8]),
    .d(pwm_start_stop[27]),
    .o(\PWMB/n23 [8]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u543 (
    .a(\PWMB/pnumr [7]),
    .b(pnumB[32]),
    .c(pnumB[7]),
    .d(pwm_start_stop[27]),
    .o(\PWMB/n23 [7]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u544 (
    .a(\PWMB/pnumr [6]),
    .b(pnumB[32]),
    .c(pnumB[6]),
    .d(pwm_start_stop[27]),
    .o(\PWMB/n23 [6]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u545 (
    .a(\PWMB/pnumr [5]),
    .b(pnumB[32]),
    .c(pnumB[5]),
    .d(pwm_start_stop[27]),
    .o(\PWMB/n23 [5]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u546 (
    .a(\PWMB/pnumr [4]),
    .b(pnumB[32]),
    .c(pnumB[4]),
    .d(pwm_start_stop[27]),
    .o(\PWMB/n23 [4]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u547 (
    .a(\PWMB/pnumr [31]),
    .b(pnumB[31]),
    .c(pnumB[32]),
    .d(pwm_start_stop[27]),
    .o(\PWMB/n23 [31]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u548 (
    .a(\PWMB/pnumr [30]),
    .b(pnumB[30]),
    .c(pnumB[32]),
    .d(pwm_start_stop[27]),
    .o(\PWMB/n23 [30]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u549 (
    .a(\PWMB/pnumr [3]),
    .b(pnumB[3]),
    .c(pnumB[32]),
    .d(pwm_start_stop[27]),
    .o(\PWMB/n23 [3]));
  EF2_PHY_SPAD #(
    //.LOCATION("p75"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u55 (
    .do({open_n1323,gpio_out_pad[15]}),
    .ts(1'b1),
    .opad(gpio_out[15]));  // CPLD_SOC_AHB_TOP.v(8)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u550 (
    .a(\PWMB/pnumr [29]),
    .b(pnumB[29]),
    .c(pnumB[32]),
    .d(pwm_start_stop[27]),
    .o(\PWMB/n23 [29]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u551 (
    .a(\PWMB/pnumr [28]),
    .b(pnumB[28]),
    .c(pnumB[32]),
    .d(pwm_start_stop[27]),
    .o(\PWMB/n23 [28]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u552 (
    .a(\PWMB/pnumr [27]),
    .b(pnumB[27]),
    .c(pnumB[32]),
    .d(pwm_start_stop[27]),
    .o(\PWMB/n23 [27]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u553 (
    .a(\PWMB/pnumr [26]),
    .b(pnumB[26]),
    .c(pnumB[32]),
    .d(pwm_start_stop[27]),
    .o(\PWMB/n23 [26]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u554 (
    .a(\PWMB/pnumr [25]),
    .b(pnumB[25]),
    .c(pnumB[32]),
    .d(pwm_start_stop[27]),
    .o(\PWMB/n23 [25]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u555 (
    .a(\PWMB/pnumr [24]),
    .b(pnumB[24]),
    .c(pnumB[32]),
    .d(pwm_start_stop[27]),
    .o(\PWMB/n23 [24]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u556 (
    .a(\PWMB/pnumr [23]),
    .b(pnumB[23]),
    .c(pnumB[32]),
    .d(pwm_start_stop[27]),
    .o(\PWMB/n23 [23]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u557 (
    .a(\PWMB/pnumr [22]),
    .b(pnumB[22]),
    .c(pnumB[32]),
    .d(pwm_start_stop[27]),
    .o(\PWMB/n23 [22]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u558 (
    .a(\PWMB/pnumr [21]),
    .b(pnumB[21]),
    .c(pnumB[32]),
    .d(pwm_start_stop[27]),
    .o(\PWMB/n23 [21]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u559 (
    .a(\PWMB/pnumr [20]),
    .b(pnumB[20]),
    .c(pnumB[32]),
    .d(pwm_start_stop[27]),
    .o(\PWMB/n23 [20]));
  EF2_PHY_SPAD #(
    //.LOCATION("p9"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u56 (
    .do({open_n1332,gpio_out_pad[14]}),
    .ts(1'b1),
    .opad(gpio_out[14]));  // CPLD_SOC_AHB_TOP.v(8)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u560 (
    .a(\PWMB/pnumr [2]),
    .b(pnumB[2]),
    .c(pnumB[32]),
    .d(pwm_start_stop[27]),
    .o(\PWMB/n23 [2]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u561 (
    .a(\PWMB/pnumr [19]),
    .b(pnumB[19]),
    .c(pnumB[32]),
    .d(pwm_start_stop[27]),
    .o(\PWMB/n23 [19]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u562 (
    .a(\PWMB/pnumr [18]),
    .b(pnumB[18]),
    .c(pnumB[32]),
    .d(pwm_start_stop[27]),
    .o(\PWMB/n23 [18]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u563 (
    .a(\PWMB/pnumr [17]),
    .b(pnumB[17]),
    .c(pnumB[32]),
    .d(pwm_start_stop[27]),
    .o(\PWMB/n23 [17]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u564 (
    .a(\PWMB/pnumr [16]),
    .b(pnumB[16]),
    .c(pnumB[32]),
    .d(pwm_start_stop[27]),
    .o(\PWMB/n23 [16]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u565 (
    .a(\PWMB/pnumr [15]),
    .b(pnumB[15]),
    .c(pnumB[32]),
    .d(pwm_start_stop[27]),
    .o(\PWMB/n23 [15]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u566 (
    .a(\PWMB/pnumr [14]),
    .b(pnumB[14]),
    .c(pnumB[32]),
    .d(pwm_start_stop[27]),
    .o(\PWMB/n23 [14]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u567 (
    .a(\PWMB/pnumr [13]),
    .b(pnumB[13]),
    .c(pnumB[32]),
    .d(pwm_start_stop[27]),
    .o(\PWMB/n23 [13]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u568 (
    .a(\PWMB/pnumr [12]),
    .b(pnumB[12]),
    .c(pnumB[32]),
    .d(pwm_start_stop[27]),
    .o(\PWMB/n23 [12]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u569 (
    .a(\PWMB/pnumr [11]),
    .b(pnumB[11]),
    .c(pnumB[32]),
    .d(pwm_start_stop[27]),
    .o(\PWMB/n23 [11]));
  EF2_PHY_PAD #(
    //.LOCATION("p139"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u57 (
    .do({open_n1340,open_n1341,open_n1342,gpio_out_pad[13]}),
    .opad(gpio_out[13]));  // CPLD_SOC_AHB_TOP.v(8)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u570 (
    .a(\PWMB/pnumr [10]),
    .b(pnumB[10]),
    .c(pnumB[32]),
    .d(pwm_start_stop[27]),
    .o(\PWMB/n23 [10]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u571 (
    .a(\PWMB/pnumr [1]),
    .b(pnumB[1]),
    .c(pnumB[32]),
    .d(pwm_start_stop[27]),
    .o(\PWMB/n23 [1]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u572 (
    .a(\PWMB/pnumr [0]),
    .b(pnumB[0]),
    .c(pnumB[32]),
    .d(pwm_start_stop[27]),
    .o(\PWMB/n23 [0]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u573 (
    .a(\PWMC/pnumr [9]),
    .b(pnumC[32]),
    .c(pnumC[9]),
    .d(pwm_start_stop[28]),
    .o(\PWMC/n23 [9]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u574 (
    .a(\PWMC/pnumr [8]),
    .b(pnumC[32]),
    .c(pnumC[8]),
    .d(pwm_start_stop[28]),
    .o(\PWMC/n23 [8]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u575 (
    .a(\PWMC/pnumr [7]),
    .b(pnumC[32]),
    .c(pnumC[7]),
    .d(pwm_start_stop[28]),
    .o(\PWMC/n23 [7]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u576 (
    .a(\PWMC/pnumr [6]),
    .b(pnumC[32]),
    .c(pnumC[6]),
    .d(pwm_start_stop[28]),
    .o(\PWMC/n23 [6]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u577 (
    .a(\PWMC/pnumr [5]),
    .b(pnumC[32]),
    .c(pnumC[5]),
    .d(pwm_start_stop[28]),
    .o(\PWMC/n23 [5]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u578 (
    .a(\PWMC/pnumr [4]),
    .b(pnumC[32]),
    .c(pnumC[4]),
    .d(pwm_start_stop[28]),
    .o(\PWMC/n23 [4]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u579 (
    .a(\PWMC/pnumr [31]),
    .b(pnumC[31]),
    .c(pnumC[32]),
    .d(pwm_start_stop[28]),
    .o(\PWMC/n23 [31]));
  EF2_PHY_SPAD #(
    //.LOCATION("p76"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u58 (
    .do({open_n1364,gpio_out_pad[12]}),
    .ts(1'b1),
    .opad(gpio_out[12]));  // CPLD_SOC_AHB_TOP.v(8)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u580 (
    .a(\PWMC/pnumr [30]),
    .b(pnumC[30]),
    .c(pnumC[32]),
    .d(pwm_start_stop[28]),
    .o(\PWMC/n23 [30]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u581 (
    .a(\PWMC/pnumr [3]),
    .b(pnumC[3]),
    .c(pnumC[32]),
    .d(pwm_start_stop[28]),
    .o(\PWMC/n23 [3]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u582 (
    .a(\PWMC/pnumr [29]),
    .b(pnumC[29]),
    .c(pnumC[32]),
    .d(pwm_start_stop[28]),
    .o(\PWMC/n23 [29]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u583 (
    .a(\PWMC/pnumr [28]),
    .b(pnumC[28]),
    .c(pnumC[32]),
    .d(pwm_start_stop[28]),
    .o(\PWMC/n23 [28]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u584 (
    .a(\PWMC/pnumr [27]),
    .b(pnumC[27]),
    .c(pnumC[32]),
    .d(pwm_start_stop[28]),
    .o(\PWMC/n23 [27]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u585 (
    .a(\PWMC/pnumr [26]),
    .b(pnumC[26]),
    .c(pnumC[32]),
    .d(pwm_start_stop[28]),
    .o(\PWMC/n23 [26]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u586 (
    .a(\PWMC/pnumr [25]),
    .b(pnumC[25]),
    .c(pnumC[32]),
    .d(pwm_start_stop[28]),
    .o(\PWMC/n23 [25]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u587 (
    .a(\PWMC/pnumr [24]),
    .b(pnumC[24]),
    .c(pnumC[32]),
    .d(pwm_start_stop[28]),
    .o(\PWMC/n23 [24]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u588 (
    .a(\PWMC/pnumr [23]),
    .b(pnumC[23]),
    .c(pnumC[32]),
    .d(pwm_start_stop[28]),
    .o(\PWMC/n23 [23]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u589 (
    .a(\PWMC/pnumr [22]),
    .b(pnumC[22]),
    .c(pnumC[32]),
    .d(pwm_start_stop[28]),
    .o(\PWMC/n23 [22]));
  EF2_PHY_SPAD #(
    //.LOCATION("p83"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u59 (
    .do({open_n1373,gpio_out_pad[11]}),
    .ts(1'b1),
    .opad(gpio_out[11]));  // CPLD_SOC_AHB_TOP.v(8)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u590 (
    .a(\PWMC/pnumr [21]),
    .b(pnumC[21]),
    .c(pnumC[32]),
    .d(pwm_start_stop[28]),
    .o(\PWMC/n23 [21]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u591 (
    .a(\PWMC/pnumr [20]),
    .b(pnumC[20]),
    .c(pnumC[32]),
    .d(pwm_start_stop[28]),
    .o(\PWMC/n23 [20]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u592 (
    .a(\PWMC/pnumr [2]),
    .b(pnumC[2]),
    .c(pnumC[32]),
    .d(pwm_start_stop[28]),
    .o(\PWMC/n23 [2]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u593 (
    .a(\PWMC/pnumr [19]),
    .b(pnumC[19]),
    .c(pnumC[32]),
    .d(pwm_start_stop[28]),
    .o(\PWMC/n23 [19]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u594 (
    .a(\PWMC/pnumr [18]),
    .b(pnumC[18]),
    .c(pnumC[32]),
    .d(pwm_start_stop[28]),
    .o(\PWMC/n23 [18]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u595 (
    .a(\PWMC/pnumr [17]),
    .b(pnumC[17]),
    .c(pnumC[32]),
    .d(pwm_start_stop[28]),
    .o(\PWMC/n23 [17]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u596 (
    .a(\PWMC/pnumr [16]),
    .b(pnumC[16]),
    .c(pnumC[32]),
    .d(pwm_start_stop[28]),
    .o(\PWMC/n23 [16]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u597 (
    .a(\PWMC/pnumr [15]),
    .b(pnumC[15]),
    .c(pnumC[32]),
    .d(pwm_start_stop[28]),
    .o(\PWMC/n23 [15]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u598 (
    .a(\PWMC/pnumr [14]),
    .b(pnumC[14]),
    .c(pnumC[32]),
    .d(pwm_start_stop[28]),
    .o(\PWMC/n23 [14]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u599 (
    .a(\PWMC/pnumr [13]),
    .b(pnumC[13]),
    .c(pnumC[32]),
    .d(pwm_start_stop[28]),
    .o(\PWMC/n23 [13]));
  EF2_PHY_SPAD #(
    //.LOCATION("p12"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u60 (
    .do({open_n1382,gpio_out_pad[10]}),
    .ts(1'b1),
    .opad(gpio_out[10]));  // CPLD_SOC_AHB_TOP.v(8)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u600 (
    .a(\PWMC/pnumr [12]),
    .b(pnumC[12]),
    .c(pnumC[32]),
    .d(pwm_start_stop[28]),
    .o(\PWMC/n23 [12]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u601 (
    .a(\PWMC/pnumr [11]),
    .b(pnumC[11]),
    .c(pnumC[32]),
    .d(pwm_start_stop[28]),
    .o(\PWMC/n23 [11]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u602 (
    .a(\PWMC/pnumr [10]),
    .b(pnumC[10]),
    .c(pnumC[32]),
    .d(pwm_start_stop[28]),
    .o(\PWMC/n23 [10]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u603 (
    .a(\PWMC/pnumr [1]),
    .b(pnumC[1]),
    .c(pnumC[32]),
    .d(pwm_start_stop[28]),
    .o(\PWMC/n23 [1]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u604 (
    .a(\PWMC/pnumr [0]),
    .b(pnumC[0]),
    .c(pnumC[32]),
    .d(pwm_start_stop[28]),
    .o(\PWMC/n23 [0]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u605 (
    .a(\PWMD/pnumr [9]),
    .b(pnumD[32]),
    .c(pnumD[9]),
    .d(pwm_start_stop[29]),
    .o(\PWMD/n23 [9]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u606 (
    .a(\PWMD/pnumr [8]),
    .b(pnumD[32]),
    .c(pnumD[8]),
    .d(pwm_start_stop[29]),
    .o(\PWMD/n23 [8]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u607 (
    .a(\PWMD/pnumr [7]),
    .b(pnumD[32]),
    .c(pnumD[7]),
    .d(pwm_start_stop[29]),
    .o(\PWMD/n23 [7]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u608 (
    .a(\PWMD/pnumr [6]),
    .b(pnumD[32]),
    .c(pnumD[6]),
    .d(pwm_start_stop[29]),
    .o(\PWMD/n23 [6]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u609 (
    .a(\PWMD/pnumr [5]),
    .b(pnumD[32]),
    .c(pnumD[5]),
    .d(pwm_start_stop[29]),
    .o(\PWMD/n23 [5]));
  EF2_PHY_SPAD #(
    //.LOCATION("p77"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u61 (
    .do({open_n1391,gpio_out_pad[9]}),
    .ts(1'b1),
    .opad(gpio_out[9]));  // CPLD_SOC_AHB_TOP.v(8)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u610 (
    .a(\PWMD/pnumr [4]),
    .b(pnumD[32]),
    .c(pnumD[4]),
    .d(pwm_start_stop[29]),
    .o(\PWMD/n23 [4]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u611 (
    .a(\PWMD/pnumr [31]),
    .b(pnumD[31]),
    .c(pnumD[32]),
    .d(pwm_start_stop[29]),
    .o(\PWMD/n23 [31]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u612 (
    .a(\PWMD/pnumr [30]),
    .b(pnumD[30]),
    .c(pnumD[32]),
    .d(pwm_start_stop[29]),
    .o(\PWMD/n23 [30]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u613 (
    .a(\PWMD/pnumr [3]),
    .b(pnumD[3]),
    .c(pnumD[32]),
    .d(pwm_start_stop[29]),
    .o(\PWMD/n23 [3]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u614 (
    .a(\PWMD/pnumr [29]),
    .b(pnumD[29]),
    .c(pnumD[32]),
    .d(pwm_start_stop[29]),
    .o(\PWMD/n23 [29]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u615 (
    .a(\PWMD/pnumr [28]),
    .b(pnumD[28]),
    .c(pnumD[32]),
    .d(pwm_start_stop[29]),
    .o(\PWMD/n23 [28]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u616 (
    .a(\PWMD/pnumr [27]),
    .b(pnumD[27]),
    .c(pnumD[32]),
    .d(pwm_start_stop[29]),
    .o(\PWMD/n23 [27]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u617 (
    .a(\PWMD/pnumr [26]),
    .b(pnumD[26]),
    .c(pnumD[32]),
    .d(pwm_start_stop[29]),
    .o(\PWMD/n23 [26]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u618 (
    .a(\PWMD/pnumr [25]),
    .b(pnumD[25]),
    .c(pnumD[32]),
    .d(pwm_start_stop[29]),
    .o(\PWMD/n23 [25]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u619 (
    .a(\PWMD/pnumr [24]),
    .b(pnumD[24]),
    .c(pnumD[32]),
    .d(pwm_start_stop[29]),
    .o(\PWMD/n23 [24]));
  EF2_PHY_SPAD #(
    //.LOCATION("p84"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u62 (
    .do({open_n1400,gpio_out_pad[8]}),
    .ts(1'b1),
    .opad(gpio_out[8]));  // CPLD_SOC_AHB_TOP.v(8)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u620 (
    .a(\PWMD/pnumr [23]),
    .b(pnumD[23]),
    .c(pnumD[32]),
    .d(pwm_start_stop[29]),
    .o(\PWMD/n23 [23]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u621 (
    .a(\PWMD/pnumr [22]),
    .b(pnumD[22]),
    .c(pnumD[32]),
    .d(pwm_start_stop[29]),
    .o(\PWMD/n23 [22]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u622 (
    .a(\PWMD/pnumr [21]),
    .b(pnumD[21]),
    .c(pnumD[32]),
    .d(pwm_start_stop[29]),
    .o(\PWMD/n23 [21]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u623 (
    .a(\PWMD/pnumr [20]),
    .b(pnumD[20]),
    .c(pnumD[32]),
    .d(pwm_start_stop[29]),
    .o(\PWMD/n23 [20]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u624 (
    .a(\PWMD/pnumr [2]),
    .b(pnumD[2]),
    .c(pnumD[32]),
    .d(pwm_start_stop[29]),
    .o(\PWMD/n23 [2]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u625 (
    .a(\PWMD/pnumr [19]),
    .b(pnumD[19]),
    .c(pnumD[32]),
    .d(pwm_start_stop[29]),
    .o(\PWMD/n23 [19]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u626 (
    .a(\PWMD/pnumr [18]),
    .b(pnumD[18]),
    .c(pnumD[32]),
    .d(pwm_start_stop[29]),
    .o(\PWMD/n23 [18]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u627 (
    .a(\PWMD/pnumr [17]),
    .b(pnumD[17]),
    .c(pnumD[32]),
    .d(pwm_start_stop[29]),
    .o(\PWMD/n23 [17]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u628 (
    .a(\PWMD/pnumr [16]),
    .b(pnumD[16]),
    .c(pnumD[32]),
    .d(pwm_start_stop[29]),
    .o(\PWMD/n23 [16]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u629 (
    .a(\PWMD/pnumr [15]),
    .b(pnumD[15]),
    .c(pnumD[32]),
    .d(pwm_start_stop[29]),
    .o(\PWMD/n23 [15]));
  EF2_PHY_SPAD #(
    //.LOCATION("p14"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u63 (
    .do({open_n1409,gpio_out_pad[7]}),
    .ts(1'b1),
    .opad(gpio_out[7]));  // CPLD_SOC_AHB_TOP.v(8)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u630 (
    .a(\PWMD/pnumr [14]),
    .b(pnumD[14]),
    .c(pnumD[32]),
    .d(pwm_start_stop[29]),
    .o(\PWMD/n23 [14]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u631 (
    .a(\PWMD/pnumr [13]),
    .b(pnumD[13]),
    .c(pnumD[32]),
    .d(pwm_start_stop[29]),
    .o(\PWMD/n23 [13]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u632 (
    .a(\PWMD/pnumr [12]),
    .b(pnumD[12]),
    .c(pnumD[32]),
    .d(pwm_start_stop[29]),
    .o(\PWMD/n23 [12]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u633 (
    .a(\PWMD/pnumr [11]),
    .b(pnumD[11]),
    .c(pnumD[32]),
    .d(pwm_start_stop[29]),
    .o(\PWMD/n23 [11]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u634 (
    .a(\PWMD/pnumr [10]),
    .b(pnumD[10]),
    .c(pnumD[32]),
    .d(pwm_start_stop[29]),
    .o(\PWMD/n23 [10]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u635 (
    .a(\PWMD/pnumr [1]),
    .b(pnumD[1]),
    .c(pnumD[32]),
    .d(pwm_start_stop[29]),
    .o(\PWMD/n23 [1]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u636 (
    .a(\PWMD/pnumr [0]),
    .b(pnumD[0]),
    .c(pnumD[32]),
    .d(pwm_start_stop[29]),
    .o(\PWMD/n23 [0]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u637 (
    .a(\PWME/pnumr [9]),
    .b(pnumE[32]),
    .c(pnumE[9]),
    .d(pwm_start_stop[30]),
    .o(\PWME/n23 [9]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u638 (
    .a(\PWME/pnumr [8]),
    .b(pnumE[32]),
    .c(pnumE[8]),
    .d(pwm_start_stop[30]),
    .o(\PWME/n23 [8]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u639 (
    .a(\PWME/pnumr [7]),
    .b(pnumE[32]),
    .c(pnumE[7]),
    .d(pwm_start_stop[30]),
    .o(\PWME/n23 [7]));
  EF2_PHY_SPAD #(
    //.LOCATION("p78"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u64 (
    .do({open_n1418,gpio_out_pad[6]}),
    .ts(1'b1),
    .opad(gpio_out[6]));  // CPLD_SOC_AHB_TOP.v(8)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u640 (
    .a(\PWME/pnumr [6]),
    .b(pnumE[32]),
    .c(pnumE[6]),
    .d(pwm_start_stop[30]),
    .o(\PWME/n23 [6]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u641 (
    .a(\PWME/pnumr [5]),
    .b(pnumE[32]),
    .c(pnumE[5]),
    .d(pwm_start_stop[30]),
    .o(\PWME/n23 [5]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u642 (
    .a(\PWME/pnumr [4]),
    .b(pnumE[32]),
    .c(pnumE[4]),
    .d(pwm_start_stop[30]),
    .o(\PWME/n23 [4]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u643 (
    .a(\PWME/pnumr [31]),
    .b(pnumE[31]),
    .c(pnumE[32]),
    .d(pwm_start_stop[30]),
    .o(\PWME/n23 [31]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u644 (
    .a(\PWME/pnumr [30]),
    .b(pnumE[30]),
    .c(pnumE[32]),
    .d(pwm_start_stop[30]),
    .o(\PWME/n23 [30]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u645 (
    .a(\PWME/pnumr [3]),
    .b(pnumE[3]),
    .c(pnumE[32]),
    .d(pwm_start_stop[30]),
    .o(\PWME/n23 [3]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u646 (
    .a(\PWME/pnumr [29]),
    .b(pnumE[29]),
    .c(pnumE[32]),
    .d(pwm_start_stop[30]),
    .o(\PWME/n23 [29]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u647 (
    .a(\PWME/pnumr [28]),
    .b(pnumE[28]),
    .c(pnumE[32]),
    .d(pwm_start_stop[30]),
    .o(\PWME/n23 [28]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u648 (
    .a(\PWME/pnumr [27]),
    .b(pnumE[27]),
    .c(pnumE[32]),
    .d(pwm_start_stop[30]),
    .o(\PWME/n23 [27]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u649 (
    .a(\PWME/pnumr [26]),
    .b(pnumE[26]),
    .c(pnumE[32]),
    .d(pwm_start_stop[30]),
    .o(\PWME/n23 [26]));
  EF2_PHY_SPAD #(
    //.LOCATION("p97"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u65 (
    .do({open_n1427,gpio_out_pad[5]}),
    .ts(1'b1),
    .opad(gpio_out[5]));  // CPLD_SOC_AHB_TOP.v(8)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u650 (
    .a(\PWME/pnumr [25]),
    .b(pnumE[25]),
    .c(pnumE[32]),
    .d(pwm_start_stop[30]),
    .o(\PWME/n23 [25]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u651 (
    .a(\PWME/pnumr [24]),
    .b(pnumE[24]),
    .c(pnumE[32]),
    .d(pwm_start_stop[30]),
    .o(\PWME/n23 [24]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u652 (
    .a(\PWME/pnumr [23]),
    .b(pnumE[23]),
    .c(pnumE[32]),
    .d(pwm_start_stop[30]),
    .o(\PWME/n23 [23]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u653 (
    .a(\PWME/pnumr [22]),
    .b(pnumE[22]),
    .c(pnumE[32]),
    .d(pwm_start_stop[30]),
    .o(\PWME/n23 [22]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u654 (
    .a(\PWME/pnumr [21]),
    .b(pnumE[21]),
    .c(pnumE[32]),
    .d(pwm_start_stop[30]),
    .o(\PWME/n23 [21]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u655 (
    .a(\PWME/pnumr [20]),
    .b(pnumE[20]),
    .c(pnumE[32]),
    .d(pwm_start_stop[30]),
    .o(\PWME/n23 [20]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u656 (
    .a(\PWME/pnumr [2]),
    .b(pnumE[2]),
    .c(pnumE[32]),
    .d(pwm_start_stop[30]),
    .o(\PWME/n23 [2]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u657 (
    .a(\PWME/pnumr [19]),
    .b(pnumE[19]),
    .c(pnumE[32]),
    .d(pwm_start_stop[30]),
    .o(\PWME/n23 [19]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u658 (
    .a(\PWME/pnumr [18]),
    .b(pnumE[18]),
    .c(pnumE[32]),
    .d(pwm_start_stop[30]),
    .o(\PWME/n23 [18]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u659 (
    .a(\PWME/pnumr [17]),
    .b(pnumE[17]),
    .c(pnumE[32]),
    .d(pwm_start_stop[30]),
    .o(\PWME/n23 [17]));
  EF2_PHY_SPAD #(
    //.LOCATION("p15"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u66 (
    .do({open_n1436,gpio_out_pad[4]}),
    .ts(1'b1),
    .opad(gpio_out[4]));  // CPLD_SOC_AHB_TOP.v(8)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u660 (
    .a(\PWME/pnumr [16]),
    .b(pnumE[16]),
    .c(pnumE[32]),
    .d(pwm_start_stop[30]),
    .o(\PWME/n23 [16]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u661 (
    .a(\PWME/pnumr [15]),
    .b(pnumE[15]),
    .c(pnumE[32]),
    .d(pwm_start_stop[30]),
    .o(\PWME/n23 [15]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u662 (
    .a(\PWME/pnumr [14]),
    .b(pnumE[14]),
    .c(pnumE[32]),
    .d(pwm_start_stop[30]),
    .o(\PWME/n23 [14]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u663 (
    .a(\PWME/pnumr [13]),
    .b(pnumE[13]),
    .c(pnumE[32]),
    .d(pwm_start_stop[30]),
    .o(\PWME/n23 [13]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u664 (
    .a(\PWME/pnumr [12]),
    .b(pnumE[12]),
    .c(pnumE[32]),
    .d(pwm_start_stop[30]),
    .o(\PWME/n23 [12]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u665 (
    .a(\PWME/pnumr [11]),
    .b(pnumE[11]),
    .c(pnumE[32]),
    .d(pwm_start_stop[30]),
    .o(\PWME/n23 [11]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u666 (
    .a(\PWME/pnumr [10]),
    .b(pnumE[10]),
    .c(pnumE[32]),
    .d(pwm_start_stop[30]),
    .o(\PWME/n23 [10]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u667 (
    .a(\PWME/pnumr [1]),
    .b(pnumE[1]),
    .c(pnumE[32]),
    .d(pwm_start_stop[30]),
    .o(\PWME/n23 [1]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u668 (
    .a(\PWME/pnumr [0]),
    .b(pnumE[0]),
    .c(pnumE[32]),
    .d(pwm_start_stop[30]),
    .o(\PWME/n23 [0]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u669 (
    .a(\PWMF/pnumr [9]),
    .b(pnumF[32]),
    .c(pnumF[9]),
    .d(pwm_start_stop[31]),
    .o(\PWMF/n23 [9]));
  EF2_PHY_SPAD #(
    //.LOCATION("p92"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u67 (
    .do({open_n1445,gpio_out_pad[3]}),
    .ts(1'b1),
    .opad(gpio_out[3]));  // CPLD_SOC_AHB_TOP.v(8)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u670 (
    .a(\PWMF/pnumr [8]),
    .b(pnumF[32]),
    .c(pnumF[8]),
    .d(pwm_start_stop[31]),
    .o(\PWMF/n23 [8]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u671 (
    .a(\PWMF/pnumr [7]),
    .b(pnumF[32]),
    .c(pnumF[7]),
    .d(pwm_start_stop[31]),
    .o(\PWMF/n23 [7]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u672 (
    .a(\PWMF/pnumr [6]),
    .b(pnumF[32]),
    .c(pnumF[6]),
    .d(pwm_start_stop[31]),
    .o(\PWMF/n23 [6]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u673 (
    .a(\PWMF/pnumr [5]),
    .b(pnumF[32]),
    .c(pnumF[5]),
    .d(pwm_start_stop[31]),
    .o(\PWMF/n23 [5]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(C)*~(B)+(~D*A)*C*~(B)+~((~D*A))*C*B+(~D*A)*C*B)"),
    .INIT(16'hc0e2))
    _al_u674 (
    .a(\PWMF/pnumr [4]),
    .b(pnumF[32]),
    .c(pnumF[4]),
    .d(pwm_start_stop[31]),
    .o(\PWMF/n23 [4]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u675 (
    .a(\PWMF/pnumr [31]),
    .b(pnumF[31]),
    .c(pnumF[32]),
    .d(pwm_start_stop[31]),
    .o(\PWMF/n23 [31]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u676 (
    .a(\PWMF/pnumr [30]),
    .b(pnumF[30]),
    .c(pnumF[32]),
    .d(pwm_start_stop[31]),
    .o(\PWMF/n23 [30]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u677 (
    .a(\PWMF/pnumr [3]),
    .b(pnumF[3]),
    .c(pnumF[32]),
    .d(pwm_start_stop[31]),
    .o(\PWMF/n23 [3]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u678 (
    .a(\PWMF/pnumr [29]),
    .b(pnumF[29]),
    .c(pnumF[32]),
    .d(pwm_start_stop[31]),
    .o(\PWMF/n23 [29]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u679 (
    .a(\PWMF/pnumr [28]),
    .b(pnumF[28]),
    .c(pnumF[32]),
    .d(pwm_start_stop[31]),
    .o(\PWMF/n23 [28]));
  EF2_PHY_SPAD #(
    //.LOCATION("p17"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u68 (
    .do({open_n1454,gpio_out_pad[2]}),
    .ts(1'b1),
    .opad(gpio_out[2]));  // CPLD_SOC_AHB_TOP.v(8)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u680 (
    .a(\PWMF/pnumr [27]),
    .b(pnumF[27]),
    .c(pnumF[32]),
    .d(pwm_start_stop[31]),
    .o(\PWMF/n23 [27]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u681 (
    .a(\PWMF/pnumr [26]),
    .b(pnumF[26]),
    .c(pnumF[32]),
    .d(pwm_start_stop[31]),
    .o(\PWMF/n23 [26]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u682 (
    .a(\PWMF/pnumr [25]),
    .b(pnumF[25]),
    .c(pnumF[32]),
    .d(pwm_start_stop[31]),
    .o(\PWMF/n23 [25]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u683 (
    .a(\PWMF/pnumr [24]),
    .b(pnumF[24]),
    .c(pnumF[32]),
    .d(pwm_start_stop[31]),
    .o(\PWMF/n23 [24]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u684 (
    .a(\PWMF/pnumr [23]),
    .b(pnumF[23]),
    .c(pnumF[32]),
    .d(pwm_start_stop[31]),
    .o(\PWMF/n23 [23]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u685 (
    .a(\PWMF/pnumr [22]),
    .b(pnumF[22]),
    .c(pnumF[32]),
    .d(pwm_start_stop[31]),
    .o(\PWMF/n23 [22]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u686 (
    .a(\PWMF/pnumr [21]),
    .b(pnumF[21]),
    .c(pnumF[32]),
    .d(pwm_start_stop[31]),
    .o(\PWMF/n23 [21]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u687 (
    .a(\PWMF/pnumr [20]),
    .b(pnumF[20]),
    .c(pnumF[32]),
    .d(pwm_start_stop[31]),
    .o(\PWMF/n23 [20]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u688 (
    .a(\PWMF/pnumr [2]),
    .b(pnumF[2]),
    .c(pnumF[32]),
    .d(pwm_start_stop[31]),
    .o(\PWMF/n23 [2]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u689 (
    .a(\PWMF/pnumr [19]),
    .b(pnumF[19]),
    .c(pnumF[32]),
    .d(pwm_start_stop[31]),
    .o(\PWMF/n23 [19]));
  EF2_PHY_SPAD #(
    //.LOCATION("p93"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u69 (
    .do({open_n1463,gpio_out_pad[1]}),
    .ts(1'b1),
    .opad(gpio_out[1]));  // CPLD_SOC_AHB_TOP.v(8)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u690 (
    .a(\PWMF/pnumr [18]),
    .b(pnumF[18]),
    .c(pnumF[32]),
    .d(pwm_start_stop[31]),
    .o(\PWMF/n23 [18]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u691 (
    .a(\PWMF/pnumr [17]),
    .b(pnumF[17]),
    .c(pnumF[32]),
    .d(pwm_start_stop[31]),
    .o(\PWMF/n23 [17]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u692 (
    .a(\PWMF/pnumr [16]),
    .b(pnumF[16]),
    .c(pnumF[32]),
    .d(pwm_start_stop[31]),
    .o(\PWMF/n23 [16]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u693 (
    .a(\PWMF/pnumr [15]),
    .b(pnumF[15]),
    .c(pnumF[32]),
    .d(pwm_start_stop[31]),
    .o(\PWMF/n23 [15]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u694 (
    .a(\PWMF/pnumr [14]),
    .b(pnumF[14]),
    .c(pnumF[32]),
    .d(pwm_start_stop[31]),
    .o(\PWMF/n23 [14]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u695 (
    .a(\PWMF/pnumr [13]),
    .b(pnumF[13]),
    .c(pnumF[32]),
    .d(pwm_start_stop[31]),
    .o(\PWMF/n23 [13]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u696 (
    .a(\PWMF/pnumr [12]),
    .b(pnumF[12]),
    .c(pnumF[32]),
    .d(pwm_start_stop[31]),
    .o(\PWMF/n23 [12]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u697 (
    .a(\PWMF/pnumr [11]),
    .b(pnumF[11]),
    .c(pnumF[32]),
    .d(pwm_start_stop[31]),
    .o(\PWMF/n23 [11]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u698 (
    .a(\PWMF/pnumr [10]),
    .b(pnumF[10]),
    .c(pnumF[32]),
    .d(pwm_start_stop[31]),
    .o(\PWMF/n23 [10]));
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u699 (
    .a(\PWMF/pnumr [1]),
    .b(pnumF[1]),
    .c(pnumF[32]),
    .d(pwm_start_stop[31]),
    .o(\PWMF/n23 [1]));
  EF2_PHY_SPAD #(
    //.LOCATION("p98"),
    //.PCICLAMP("ON"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u70 (
    .do({open_n1472,gpio_out_pad[0]}),
    .ts(1'b1),
    .opad(gpio_out[0]));  // CPLD_SOC_AHB_TOP.v(8)
  AL_MAP_LUT4 #(
    .EQN("((~D*A)*~(B)*~(C)+(~D*A)*B*~(C)+~((~D*A))*B*C+(~D*A)*B*C)"),
    .INIT(16'hc0ca))
    _al_u700 (
    .a(\PWMF/pnumr [0]),
    .b(pnumF[0]),
    .c(pnumF[32]),
    .d(pwm_start_stop[31]),
    .o(\PWMF/n23 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u701 (
    .a(\U_AHB/h2h_hwrite ),
    .b(\U_AHB/h2h_haddr [2]),
    .c(\U_AHB/h2h_haddr [13]),
    .d(\U_AHB/h2h_haddr [14]),
    .o(\U_AHB/n8 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u702 (
    .a(\U_AHB/h2h_hwrite ),
    .b(\U_AHB/h2h_haddr [12]),
    .c(\U_AHB/h2h_haddr [13]),
    .d(\U_AHB/h2h_haddr [14]),
    .o(\U_AHB/n28 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    _al_u703 (
    .a(\U_AHB/h2h_hwrite ),
    .b(\U_AHB/h2h_haddr [13]),
    .c(\U_AHB/h2h_haddr [14]),
    .d(\U_AHB/h2h_haddr [11]),
    .o(\U_AHB/n26 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    _al_u704 (
    .a(\U_AHB/h2h_hwrite ),
    .b(\U_AHB/h2h_haddr [13]),
    .c(\U_AHB/h2h_haddr [14]),
    .d(\U_AHB/h2h_haddr [10]),
    .o(\U_AHB/n24 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    _al_u705 (
    .a(\U_AHB/h2h_hwrite ),
    .b(\U_AHB/h2h_haddr [13]),
    .c(\U_AHB/h2h_haddr [14]),
    .d(\U_AHB/h2h_haddr [9]),
    .o(\U_AHB/n22 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    _al_u706 (
    .a(\U_AHB/h2h_hwrite ),
    .b(\U_AHB/h2h_haddr [13]),
    .c(\U_AHB/h2h_haddr [14]),
    .d(\U_AHB/h2h_haddr [8]),
    .o(\U_AHB/n20 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    _al_u707 (
    .a(\U_AHB/h2h_hwrite ),
    .b(\U_AHB/h2h_haddr [13]),
    .c(\U_AHB/h2h_haddr [14]),
    .d(\U_AHB/h2h_haddr [7]),
    .o(\U_AHB/n18 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    _al_u708 (
    .a(\U_AHB/h2h_hwrite ),
    .b(\U_AHB/h2h_haddr [13]),
    .c(\U_AHB/h2h_haddr [14]),
    .d(\U_AHB/h2h_haddr [6]),
    .o(\U_AHB/n16 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    _al_u709 (
    .a(\U_AHB/h2h_hwrite ),
    .b(\U_AHB/h2h_haddr [13]),
    .c(\U_AHB/h2h_haddr [14]),
    .d(\U_AHB/h2h_haddr [5]),
    .o(\U_AHB/n14 ));
  EF2_PHY_SPAD #(
    //.LOCATION("P100"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("16"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u71 (
    .do({open_n1481,ledout_pad[3]}),
    .ts(1'b1),
    .opad(ledout[3]));  // CPLD_SOC_AHB_TOP.v(10)
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    _al_u710 (
    .a(\U_AHB/h2h_hwrite ),
    .b(\U_AHB/h2h_haddr [13]),
    .c(\U_AHB/h2h_haddr [14]),
    .d(\U_AHB/h2h_haddr [4]),
    .o(\U_AHB/n12 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u711 (
    .a(\U_AHB/h2h_hwrite ),
    .b(\U_AHB/h2h_haddr [3]),
    .c(\U_AHB/h2h_haddr [13]),
    .d(\U_AHB/h2h_haddr [14]),
    .o(\U_AHB/n10 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u712 (
    .a(\U_AHB/h2h_hwrite ),
    .b(\U_AHB/h2h_haddr [13]),
    .c(\U_AHB/h2h_haddr [14]),
    .d(\U_AHB/h2h_haddr [6]),
    .o(\U_AHB/n4 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u713 (
    .a(\U_AHB/h2h_hwrite ),
    .b(\U_AHB/h2h_haddr [13]),
    .c(\U_AHB/h2h_haddr [14]),
    .d(\U_AHB/h2h_haddr [4]),
    .o(\U_AHB/n34 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u714 (
    .a(\U_AHB/h2h_hwrite ),
    .b(\U_AHB/h2h_haddr [3]),
    .c(\U_AHB/h2h_haddr [13]),
    .d(\U_AHB/h2h_haddr [14]),
    .o(\U_AHB/n32 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u715 (
    .a(\U_AHB/h2h_hwrite ),
    .b(\U_AHB/h2h_haddr [2]),
    .c(\U_AHB/h2h_haddr [13]),
    .d(\U_AHB/h2h_haddr [14]),
    .o(\U_AHB/n30 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u716 (
    .a(\U_AHB/h2h_hwrite ),
    .b(\U_AHB/h2h_haddr [13]),
    .c(\U_AHB/h2h_haddr [14]),
    .d(\U_AHB/h2h_haddr [5]),
    .o(\U_AHB/n2 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u717 (
    .a(\U_AHB/h2h_hwrite ),
    .b(\U_AHB/h2h_haddr [12]),
    .c(\U_AHB/h2h_haddr [13]),
    .d(\U_AHB/h2h_haddr [14]),
    .o(\U_AHB/n71 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u718 (
    .a(\U_AHB/h2h_hwrite ),
    .b(\U_AHB/h2h_haddr [13]),
    .c(\U_AHB/h2h_haddr [14]),
    .d(\U_AHB/h2h_haddr [11]),
    .o(\U_AHB/n69 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u719 (
    .a(\U_AHB/h2h_hwrite ),
    .b(\U_AHB/h2h_haddr [13]),
    .c(\U_AHB/h2h_haddr [14]),
    .d(\U_AHB/h2h_haddr [10]),
    .o(\U_AHB/n67 ));
  EF2_PHY_SPAD #(
    //.LOCATION("P103"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("16"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u72 (
    .do({open_n1490,ledout_pad[2]}),
    .ts(1'b1),
    .opad(ledout[2]));  // CPLD_SOC_AHB_TOP.v(10)
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u720 (
    .a(\U_AHB/h2h_hwrite ),
    .b(\U_AHB/h2h_haddr [13]),
    .c(\U_AHB/h2h_haddr [14]),
    .d(\U_AHB/h2h_haddr [9]),
    .o(\U_AHB/n65 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u721 (
    .a(\U_AHB/h2h_hwrite ),
    .b(\U_AHB/h2h_haddr [13]),
    .c(\U_AHB/h2h_haddr [14]),
    .d(\U_AHB/h2h_haddr [8]),
    .o(\U_AHB/n63 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u722 (
    .a(\U_AHB/h2h_hwrite ),
    .b(\U_AHB/h2h_haddr [13]),
    .c(\U_AHB/h2h_haddr [14]),
    .d(\U_AHB/h2h_haddr [7]),
    .o(\U_AHB/n61 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u723 (
    .a(\U_AHB/h2h_hwrite ),
    .b(\U_AHB/h2h_haddr [13]),
    .c(\U_AHB/h2h_haddr [14]),
    .d(\U_AHB/h2h_haddr [6]),
    .o(\U_AHB/n59 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u724 (
    .a(\U_AHB/h2h_hwrite ),
    .b(\U_AHB/h2h_haddr [13]),
    .c(\U_AHB/h2h_haddr [14]),
    .d(\U_AHB/h2h_haddr [5]),
    .o(\U_AHB/n57 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u725 (
    .a(\U_AHB/h2h_hwrite ),
    .b(\U_AHB/h2h_haddr [13]),
    .c(\U_AHB/h2h_haddr [14]),
    .d(\U_AHB/h2h_haddr [4]),
    .o(\U_AHB/n55 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u726 (
    .a(\U_AHB/h2h_hwrite ),
    .b(\U_AHB/h2h_haddr [3]),
    .c(\U_AHB/h2h_haddr [13]),
    .d(\U_AHB/h2h_haddr [14]),
    .o(\U_AHB/n53 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u727 (
    .a(\U_AHB/h2h_hwrite ),
    .b(\U_AHB/h2h_haddr [2]),
    .c(\U_AHB/h2h_haddr [13]),
    .d(\U_AHB/h2h_haddr [14]),
    .o(\U_AHB/n51 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u728 (
    .a(\U_AHB/h2h_hwrite ),
    .b(\U_AHB/h2h_haddr [3]),
    .c(\U_AHB/h2h_haddr [13]),
    .d(\U_AHB/h2h_haddr [14]),
    .o(\U_AHB/n75 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u729 (
    .a(\U_AHB/h2h_hwrite ),
    .b(\U_AHB/h2h_haddr [2]),
    .c(\U_AHB/h2h_haddr [13]),
    .d(\U_AHB/h2h_haddr [14]),
    .o(\U_AHB/n73 ));
  EF2_PHY_SPAD #(
    //.LOCATION("P104"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DRIVE("16"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("INV"))
    _al_u73 (
    .do({open_n1499,ledout_pad[1]}),
    .ts(1'b1),
    .opad(ledout[1]));  // CPLD_SOC_AHB_TOP.v(10)
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u730 (
    .a(\U_AHB/h2h_hwrite ),
    .b(\U_AHB/h2h_haddr [13]),
    .c(\U_AHB/h2h_haddr [14]),
    .d(\U_AHB/h2h_haddr [6]),
    .o(\U_AHB/n47 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u731 (
    .a(\U_AHB/h2h_hwrite ),
    .b(\U_AHB/h2h_haddr [13]),
    .c(\U_AHB/h2h_haddr [14]),
    .d(\U_AHB/h2h_haddr [5]),
    .o(\U_AHB/n45 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u732 (
    .a(\U_AHB/h2h_hwrite ),
    .b(\U_AHB/h2h_haddr [13]),
    .c(\U_AHB/h2h_haddr [14]),
    .d(\U_AHB/h2h_haddr [7]),
    .o(\U_AHB/n79 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u733 (
    .a(\U_AHB/h2h_hwrite ),
    .b(\U_AHB/h2h_haddr [13]),
    .c(\U_AHB/h2h_haddr [14]),
    .d(\U_AHB/h2h_haddr [4]),
    .o(\U_AHB/n77 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u734 (
    .a(\PWM0/FreCnt [23]),
    .b(\PWM0/FreCnt [24]),
    .c(\PWM0/FreCnt [25]),
    .d(\PWM0/FreCnt [26]),
    .o(_al_u734_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u735 (
    .a(_al_u734_o),
    .b(\PWM0/FreCnt [3]),
    .c(\PWM0/FreCnt [4]),
    .d(\PWM0/FreCnt [5]),
    .e(\PWM0/FreCnt [6]),
    .o(_al_u735_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u736 (
    .a(_al_u735_o),
    .b(\PWM0/FreCnt [7]),
    .c(\PWM0/FreCnt [8]),
    .d(\PWM0/FreCnt [9]),
    .o(_al_u736_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u737 (
    .a(\PWM0/FreCnt [0]),
    .b(\PWM0/FreCnt [1]),
    .c(\PWM0/FreCnt [10]),
    .d(\PWM0/FreCnt [11]),
    .o(_al_u737_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u738 (
    .a(_al_u737_o),
    .b(\PWM0/FreCnt [12]),
    .c(\PWM0/FreCnt [13]),
    .d(\PWM0/FreCnt [14]),
    .e(\PWM0/FreCnt [15]),
    .o(_al_u738_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u739 (
    .a(\PWM0/FreCnt [16]),
    .b(\PWM0/FreCnt [17]),
    .c(\PWM0/FreCnt [18]),
    .d(\PWM0/FreCnt [19]),
    .o(_al_u739_o));
  EF2_PHY_SPAD #(
    //.LOCATION("P87"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u74 (
    .ipad(limit_l[15]),
    .ts(1'b1),
    .di(limit_l_pad[15]));  // CPLD_SOC_AHB_TOP.v(5)
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u740 (
    .a(_al_u739_o),
    .b(\PWM0/FreCnt [2]),
    .c(\PWM0/FreCnt [20]),
    .d(\PWM0/FreCnt [21]),
    .e(\PWM0/FreCnt [22]),
    .o(_al_u740_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u741 (
    .a(_al_u736_o),
    .b(_al_u738_o),
    .c(_al_u740_o),
    .o(\PWM0/n0_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u742 (
    .a(\PWM0/n0_lutinv ),
    .b(\PWM0/stopreq ),
    .o(\PWM0/n1 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u743 (
    .a(\PWM0/n0_lutinv ),
    .b(\PWM0/n11 ),
    .o(\PWM0/mux3_b0_sel_is_3_o ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u744 (
    .a(\PWM0/n0_lutinv ),
    .b(\PWM0/n12 [9]),
    .c(freq0[9]),
    .o(\PWM0/n13 [9]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u745 (
    .a(\PWM0/n0_lutinv ),
    .b(\PWM0/n12 [8]),
    .c(freq0[8]),
    .o(\PWM0/n13 [8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u746 (
    .a(\PWM0/n0_lutinv ),
    .b(\PWM0/n12 [7]),
    .c(freq0[7]),
    .o(\PWM0/n13 [7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u747 (
    .a(\PWM0/n0_lutinv ),
    .b(\PWM0/n12 [6]),
    .c(freq0[6]),
    .o(\PWM0/n13 [6]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u748 (
    .a(\PWM0/n0_lutinv ),
    .b(\PWM0/n12 [5]),
    .c(freq0[5]),
    .o(\PWM0/n13 [5]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u749 (
    .a(\PWM0/n0_lutinv ),
    .b(\PWM0/n12 [4]),
    .c(freq0[4]),
    .o(\PWM0/n13 [4]));
  EF2_PHY_SPAD #(
    //.LOCATION("P85"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u75 (
    .ipad(limit_l[14]),
    .ts(1'b1),
    .di(limit_l_pad[14]));  // CPLD_SOC_AHB_TOP.v(5)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u750 (
    .a(\PWM0/n0_lutinv ),
    .b(\PWM0/n12 [3]),
    .c(freq0[3]),
    .o(\PWM0/n13 [3]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u751 (
    .a(\PWM0/n0_lutinv ),
    .b(\PWM0/n12 [26]),
    .c(freq0[26]),
    .o(\PWM0/n13 [26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u752 (
    .a(\PWM0/n0_lutinv ),
    .b(\PWM0/n12 [25]),
    .c(freq0[25]),
    .o(\PWM0/n13 [25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u753 (
    .a(\PWM0/n0_lutinv ),
    .b(\PWM0/n12 [24]),
    .c(freq0[24]),
    .o(\PWM0/n13 [24]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u754 (
    .a(\PWM0/n0_lutinv ),
    .b(\PWM0/n12 [23]),
    .c(freq0[23]),
    .o(\PWM0/n13 [23]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u755 (
    .a(\PWM0/n0_lutinv ),
    .b(\PWM0/n12 [22]),
    .c(freq0[22]),
    .o(\PWM0/n13 [22]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u756 (
    .a(\PWM0/n0_lutinv ),
    .b(\PWM0/n12 [21]),
    .c(freq0[21]),
    .o(\PWM0/n13 [21]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u757 (
    .a(\PWM0/n0_lutinv ),
    .b(\PWM0/n12 [20]),
    .c(freq0[20]),
    .o(\PWM0/n13 [20]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u758 (
    .a(\PWM0/n0_lutinv ),
    .b(\PWM0/n12 [2]),
    .c(freq0[2]),
    .o(\PWM0/n13 [2]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u759 (
    .a(\PWM0/n0_lutinv ),
    .b(\PWM0/n12 [19]),
    .c(freq0[19]),
    .o(\PWM0/n13 [19]));
  EF2_PHY_SPAD #(
    //.LOCATION("P1"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u76 (
    .ipad(limit_l[13]),
    .ts(1'b1),
    .di(limit_l_pad[13]));  // CPLD_SOC_AHB_TOP.v(5)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u760 (
    .a(\PWM0/n0_lutinv ),
    .b(\PWM0/n12 [18]),
    .c(freq0[18]),
    .o(\PWM0/n13 [18]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u761 (
    .a(\PWM0/n0_lutinv ),
    .b(\PWM0/n12 [17]),
    .c(freq0[17]),
    .o(\PWM0/n13 [17]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u762 (
    .a(\PWM0/n0_lutinv ),
    .b(\PWM0/n12 [16]),
    .c(freq0[16]),
    .o(\PWM0/n13 [16]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u763 (
    .a(\PWM0/n0_lutinv ),
    .b(\PWM0/n12 [15]),
    .c(freq0[15]),
    .o(\PWM0/n13 [15]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u764 (
    .a(\PWM0/n0_lutinv ),
    .b(\PWM0/n12 [14]),
    .c(freq0[14]),
    .o(\PWM0/n13 [14]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u765 (
    .a(\PWM0/n0_lutinv ),
    .b(\PWM0/n12 [13]),
    .c(freq0[13]),
    .o(\PWM0/n13 [13]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u766 (
    .a(\PWM0/n0_lutinv ),
    .b(\PWM0/n12 [12]),
    .c(freq0[12]),
    .o(\PWM0/n13 [12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u767 (
    .a(\PWM0/n0_lutinv ),
    .b(\PWM0/n12 [11]),
    .c(freq0[11]),
    .o(\PWM0/n13 [11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u768 (
    .a(\PWM0/n0_lutinv ),
    .b(\PWM0/n12 [10]),
    .c(freq0[10]),
    .o(\PWM0/n13 [10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u769 (
    .a(\PWM0/n0_lutinv ),
    .b(\PWM0/n12 [1]),
    .c(freq0[1]),
    .o(\PWM0/n13 [1]));
  EF2_PHY_PAD #(
    //.LOCATION("P69"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u77 (
    .ipad(limit_l[12]),
    .di(limit_l_pad[12]));  // CPLD_SOC_AHB_TOP.v(5)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u770 (
    .a(\PWM0/n0_lutinv ),
    .b(\PWM0/n12 [0]),
    .c(freq0[0]),
    .o(\PWM0/n13 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u771 (
    .a(\PWM1/FreCnt [23]),
    .b(\PWM1/FreCnt [24]),
    .c(\PWM1/FreCnt [25]),
    .d(\PWM1/FreCnt [26]),
    .o(_al_u771_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u772 (
    .a(_al_u771_o),
    .b(\PWM1/FreCnt [3]),
    .c(\PWM1/FreCnt [4]),
    .d(\PWM1/FreCnt [5]),
    .e(\PWM1/FreCnt [6]),
    .o(_al_u772_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u773 (
    .a(_al_u772_o),
    .b(\PWM1/FreCnt [7]),
    .c(\PWM1/FreCnt [8]),
    .d(\PWM1/FreCnt [9]),
    .o(_al_u773_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u774 (
    .a(\PWM1/FreCnt [0]),
    .b(\PWM1/FreCnt [1]),
    .c(\PWM1/FreCnt [10]),
    .d(\PWM1/FreCnt [11]),
    .o(_al_u774_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u775 (
    .a(_al_u774_o),
    .b(\PWM1/FreCnt [12]),
    .c(\PWM1/FreCnt [13]),
    .d(\PWM1/FreCnt [14]),
    .e(\PWM1/FreCnt [15]),
    .o(_al_u775_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u776 (
    .a(\PWM1/FreCnt [16]),
    .b(\PWM1/FreCnt [17]),
    .c(\PWM1/FreCnt [18]),
    .d(\PWM1/FreCnt [19]),
    .o(_al_u776_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u777 (
    .a(_al_u776_o),
    .b(\PWM1/FreCnt [2]),
    .c(\PWM1/FreCnt [20]),
    .d(\PWM1/FreCnt [21]),
    .e(\PWM1/FreCnt [22]),
    .o(_al_u777_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u778 (
    .a(_al_u773_o),
    .b(_al_u775_o),
    .c(_al_u777_o),
    .o(\PWM1/n0_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u779 (
    .a(\PWM1/n0_lutinv ),
    .b(\PWM1/stopreq ),
    .o(\PWM1/n1 ));
  EF2_PHY_PAD #(
    //.LOCATION("P67"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u78 (
    .ipad(limit_l[11]),
    .di(limit_l_pad[11]));  // CPLD_SOC_AHB_TOP.v(5)
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u780 (
    .a(\PWM1/n0_lutinv ),
    .b(\PWM1/n11 ),
    .o(\PWM1/mux3_b0_sel_is_3_o ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u781 (
    .a(\PWM1/n0_lutinv ),
    .b(\PWM1/n12 [9]),
    .c(freq1[9]),
    .o(\PWM1/n13 [9]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u782 (
    .a(\PWM1/n0_lutinv ),
    .b(\PWM1/n12 [8]),
    .c(freq1[8]),
    .o(\PWM1/n13 [8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u783 (
    .a(\PWM1/n0_lutinv ),
    .b(\PWM1/n12 [7]),
    .c(freq1[7]),
    .o(\PWM1/n13 [7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u784 (
    .a(\PWM1/n0_lutinv ),
    .b(\PWM1/n12 [6]),
    .c(freq1[6]),
    .o(\PWM1/n13 [6]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u785 (
    .a(\PWM1/n0_lutinv ),
    .b(\PWM1/n12 [5]),
    .c(freq1[5]),
    .o(\PWM1/n13 [5]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u786 (
    .a(\PWM1/n0_lutinv ),
    .b(\PWM1/n12 [4]),
    .c(freq1[4]),
    .o(\PWM1/n13 [4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u787 (
    .a(\PWM1/n0_lutinv ),
    .b(\PWM1/n12 [3]),
    .c(freq1[3]),
    .o(\PWM1/n13 [3]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u788 (
    .a(\PWM1/n0_lutinv ),
    .b(\PWM1/n12 [26]),
    .c(freq1[26]),
    .o(\PWM1/n13 [26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u789 (
    .a(\PWM1/n0_lutinv ),
    .b(\PWM1/n12 [25]),
    .c(freq1[25]),
    .o(\PWM1/n13 [25]));
  EF2_PHY_PAD #(
    //.LOCATION("P65"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u79 (
    .ipad(limit_l[10]),
    .di(limit_l_pad[10]));  // CPLD_SOC_AHB_TOP.v(5)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u790 (
    .a(\PWM1/n0_lutinv ),
    .b(\PWM1/n12 [24]),
    .c(freq1[24]),
    .o(\PWM1/n13 [24]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u791 (
    .a(\PWM1/n0_lutinv ),
    .b(\PWM1/n12 [23]),
    .c(freq1[23]),
    .o(\PWM1/n13 [23]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u792 (
    .a(\PWM1/n0_lutinv ),
    .b(\PWM1/n12 [22]),
    .c(freq1[22]),
    .o(\PWM1/n13 [22]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u793 (
    .a(\PWM1/n0_lutinv ),
    .b(\PWM1/n12 [21]),
    .c(freq1[21]),
    .o(\PWM1/n13 [21]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u794 (
    .a(\PWM1/n0_lutinv ),
    .b(\PWM1/n12 [20]),
    .c(freq1[20]),
    .o(\PWM1/n13 [20]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u795 (
    .a(\PWM1/n0_lutinv ),
    .b(\PWM1/n12 [2]),
    .c(freq1[2]),
    .o(\PWM1/n13 [2]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u796 (
    .a(\PWM1/n0_lutinv ),
    .b(\PWM1/n12 [19]),
    .c(freq1[19]),
    .o(\PWM1/n13 [19]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u797 (
    .a(\PWM1/n0_lutinv ),
    .b(\PWM1/n12 [18]),
    .c(freq1[18]),
    .o(\PWM1/n13 [18]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u798 (
    .a(\PWM1/n0_lutinv ),
    .b(\PWM1/n12 [17]),
    .c(freq1[17]),
    .o(\PWM1/n13 [17]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u799 (
    .a(\PWM1/n0_lutinv ),
    .b(\PWM1/n12 [16]),
    .c(freq1[16]),
    .o(\PWM1/n13 [16]));
  EF2_PHY_SPAD #(
    //.LOCATION("P34"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u80 (
    .ipad(limit_l[9]),
    .ts(1'b1),
    .di(limit_l_pad[9]));  // CPLD_SOC_AHB_TOP.v(5)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u800 (
    .a(\PWM1/n0_lutinv ),
    .b(\PWM1/n12 [15]),
    .c(freq1[15]),
    .o(\PWM1/n13 [15]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u801 (
    .a(\PWM1/n0_lutinv ),
    .b(\PWM1/n12 [14]),
    .c(freq1[14]),
    .o(\PWM1/n13 [14]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u802 (
    .a(\PWM1/n0_lutinv ),
    .b(\PWM1/n12 [13]),
    .c(freq1[13]),
    .o(\PWM1/n13 [13]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u803 (
    .a(\PWM1/n0_lutinv ),
    .b(\PWM1/n12 [12]),
    .c(freq1[12]),
    .o(\PWM1/n13 [12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u804 (
    .a(\PWM1/n0_lutinv ),
    .b(\PWM1/n12 [11]),
    .c(freq1[11]),
    .o(\PWM1/n13 [11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u805 (
    .a(\PWM1/n0_lutinv ),
    .b(\PWM1/n12 [10]),
    .c(freq1[10]),
    .o(\PWM1/n13 [10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u806 (
    .a(\PWM1/n0_lutinv ),
    .b(\PWM1/n12 [1]),
    .c(freq1[1]),
    .o(\PWM1/n13 [1]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u807 (
    .a(\PWM1/n0_lutinv ),
    .b(\PWM1/n12 [0]),
    .c(freq1[0]),
    .o(\PWM1/n13 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u808 (
    .a(\PWM2/FreCnt [23]),
    .b(\PWM2/FreCnt [24]),
    .c(\PWM2/FreCnt [25]),
    .d(\PWM2/FreCnt [26]),
    .o(_al_u808_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u809 (
    .a(_al_u808_o),
    .b(\PWM2/FreCnt [3]),
    .c(\PWM2/FreCnt [4]),
    .d(\PWM2/FreCnt [5]),
    .e(\PWM2/FreCnt [6]),
    .o(_al_u809_o));
  EF2_PHY_SPAD #(
    //.LOCATION("P33"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u81 (
    .ipad(limit_l[8]),
    .ts(1'b1),
    .di(limit_l_pad[8]));  // CPLD_SOC_AHB_TOP.v(5)
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u810 (
    .a(_al_u809_o),
    .b(\PWM2/FreCnt [7]),
    .c(\PWM2/FreCnt [8]),
    .d(\PWM2/FreCnt [9]),
    .o(_al_u810_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u811 (
    .a(\PWM2/FreCnt [0]),
    .b(\PWM2/FreCnt [1]),
    .c(\PWM2/FreCnt [10]),
    .d(\PWM2/FreCnt [11]),
    .o(_al_u811_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u812 (
    .a(_al_u811_o),
    .b(\PWM2/FreCnt [12]),
    .c(\PWM2/FreCnt [13]),
    .d(\PWM2/FreCnt [14]),
    .e(\PWM2/FreCnt [15]),
    .o(_al_u812_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u813 (
    .a(\PWM2/FreCnt [16]),
    .b(\PWM2/FreCnt [17]),
    .c(\PWM2/FreCnt [18]),
    .d(\PWM2/FreCnt [19]),
    .o(_al_u813_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u814 (
    .a(_al_u813_o),
    .b(\PWM2/FreCnt [2]),
    .c(\PWM2/FreCnt [20]),
    .d(\PWM2/FreCnt [21]),
    .e(\PWM2/FreCnt [22]),
    .o(_al_u814_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u815 (
    .a(_al_u810_o),
    .b(_al_u812_o),
    .c(_al_u814_o),
    .o(\PWM2/n0_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u816 (
    .a(\PWM2/n0_lutinv ),
    .b(\PWM2/stopreq ),
    .o(\PWM2/n1 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u817 (
    .a(\PWM2/n0_lutinv ),
    .b(\PWM2/n11 ),
    .o(\PWM2/mux3_b0_sel_is_3_o ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u818 (
    .a(\PWM2/n0_lutinv ),
    .b(\PWM2/n12 [9]),
    .c(freq2[9]),
    .o(\PWM2/n13 [9]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u819 (
    .a(\PWM2/n0_lutinv ),
    .b(\PWM2/n12 [8]),
    .c(freq2[8]),
    .o(\PWM2/n13 [8]));
  EF2_PHY_SPAD #(
    //.LOCATION("P89"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u82 (
    .ipad(limit_l[7]),
    .ts(1'b1),
    .di(limit_l_pad[7]));  // CPLD_SOC_AHB_TOP.v(5)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u820 (
    .a(\PWM2/n0_lutinv ),
    .b(\PWM2/n12 [7]),
    .c(freq2[7]),
    .o(\PWM2/n13 [7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u821 (
    .a(\PWM2/n0_lutinv ),
    .b(\PWM2/n12 [6]),
    .c(freq2[6]),
    .o(\PWM2/n13 [6]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u822 (
    .a(\PWM2/n0_lutinv ),
    .b(\PWM2/n12 [5]),
    .c(freq2[5]),
    .o(\PWM2/n13 [5]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u823 (
    .a(\PWM2/n0_lutinv ),
    .b(\PWM2/n12 [4]),
    .c(freq2[4]),
    .o(\PWM2/n13 [4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u824 (
    .a(\PWM2/n0_lutinv ),
    .b(\PWM2/n12 [3]),
    .c(freq2[3]),
    .o(\PWM2/n13 [3]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u825 (
    .a(\PWM2/n0_lutinv ),
    .b(\PWM2/n12 [26]),
    .c(freq2[26]),
    .o(\PWM2/n13 [26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u826 (
    .a(\PWM2/n0_lutinv ),
    .b(\PWM2/n12 [25]),
    .c(freq2[25]),
    .o(\PWM2/n13 [25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u827 (
    .a(\PWM2/n0_lutinv ),
    .b(\PWM2/n12 [24]),
    .c(freq2[24]),
    .o(\PWM2/n13 [24]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u828 (
    .a(\PWM2/n0_lutinv ),
    .b(\PWM2/n12 [23]),
    .c(freq2[23]),
    .o(\PWM2/n13 [23]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u829 (
    .a(\PWM2/n0_lutinv ),
    .b(\PWM2/n12 [22]),
    .c(freq2[22]),
    .o(\PWM2/n13 [22]));
  EF2_PHY_SPAD #(
    //.LOCATION("P2"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u83 (
    .ipad(limit_l[6]),
    .ts(1'b1),
    .di(limit_l_pad[6]));  // CPLD_SOC_AHB_TOP.v(5)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u830 (
    .a(\PWM2/n0_lutinv ),
    .b(\PWM2/n12 [21]),
    .c(freq2[21]),
    .o(\PWM2/n13 [21]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u831 (
    .a(\PWM2/n0_lutinv ),
    .b(\PWM2/n12 [20]),
    .c(freq2[20]),
    .o(\PWM2/n13 [20]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u832 (
    .a(\PWM2/n0_lutinv ),
    .b(\PWM2/n12 [2]),
    .c(freq2[2]),
    .o(\PWM2/n13 [2]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u833 (
    .a(\PWM2/n0_lutinv ),
    .b(\PWM2/n12 [19]),
    .c(freq2[19]),
    .o(\PWM2/n13 [19]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u834 (
    .a(\PWM2/n0_lutinv ),
    .b(\PWM2/n12 [18]),
    .c(freq2[18]),
    .o(\PWM2/n13 [18]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u835 (
    .a(\PWM2/n0_lutinv ),
    .b(\PWM2/n12 [17]),
    .c(freq2[17]),
    .o(\PWM2/n13 [17]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u836 (
    .a(\PWM2/n0_lutinv ),
    .b(\PWM2/n12 [16]),
    .c(freq2[16]),
    .o(\PWM2/n13 [16]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u837 (
    .a(\PWM2/n0_lutinv ),
    .b(\PWM2/n12 [15]),
    .c(freq2[15]),
    .o(\PWM2/n13 [15]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u838 (
    .a(\PWM2/n0_lutinv ),
    .b(\PWM2/n12 [14]),
    .c(freq2[14]),
    .o(\PWM2/n13 [14]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u839 (
    .a(\PWM2/n0_lutinv ),
    .b(\PWM2/n12 [13]),
    .c(freq2[13]),
    .o(\PWM2/n13 [13]));
  EF2_PHY_SPAD #(
    //.LOCATION("P6"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u84 (
    .ipad(limit_l[5]),
    .ts(1'b1),
    .di(limit_l_pad[5]));  // CPLD_SOC_AHB_TOP.v(5)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u840 (
    .a(\PWM2/n0_lutinv ),
    .b(\PWM2/n12 [12]),
    .c(freq2[12]),
    .o(\PWM2/n13 [12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u841 (
    .a(\PWM2/n0_lutinv ),
    .b(\PWM2/n12 [11]),
    .c(freq2[11]),
    .o(\PWM2/n13 [11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u842 (
    .a(\PWM2/n0_lutinv ),
    .b(\PWM2/n12 [10]),
    .c(freq2[10]),
    .o(\PWM2/n13 [10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u843 (
    .a(\PWM2/n0_lutinv ),
    .b(\PWM2/n12 [1]),
    .c(freq2[1]),
    .o(\PWM2/n13 [1]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u844 (
    .a(\PWM2/n0_lutinv ),
    .b(\PWM2/n12 [0]),
    .c(freq2[0]),
    .o(\PWM2/n13 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u845 (
    .a(\PWM3/FreCnt [23]),
    .b(\PWM3/FreCnt [24]),
    .c(\PWM3/FreCnt [25]),
    .d(\PWM3/FreCnt [26]),
    .o(_al_u845_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u846 (
    .a(_al_u845_o),
    .b(\PWM3/FreCnt [3]),
    .c(\PWM3/FreCnt [4]),
    .d(\PWM3/FreCnt [5]),
    .e(\PWM3/FreCnt [6]),
    .o(_al_u846_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u847 (
    .a(_al_u846_o),
    .b(\PWM3/FreCnt [7]),
    .c(\PWM3/FreCnt [8]),
    .d(\PWM3/FreCnt [9]),
    .o(_al_u847_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u848 (
    .a(\PWM3/FreCnt [0]),
    .b(\PWM3/FreCnt [1]),
    .c(\PWM3/FreCnt [10]),
    .d(\PWM3/FreCnt [11]),
    .o(_al_u848_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u849 (
    .a(_al_u848_o),
    .b(\PWM3/FreCnt [12]),
    .c(\PWM3/FreCnt [13]),
    .d(\PWM3/FreCnt [14]),
    .e(\PWM3/FreCnt [15]),
    .o(_al_u849_o));
  EF2_PHY_PAD #(
    //.LOCATION("P60"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u85 (
    .ipad(limit_l[4]),
    .di(limit_l_pad[4]));  // CPLD_SOC_AHB_TOP.v(5)
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u850 (
    .a(\PWM3/FreCnt [16]),
    .b(\PWM3/FreCnt [17]),
    .c(\PWM3/FreCnt [18]),
    .d(\PWM3/FreCnt [19]),
    .o(_al_u850_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u851 (
    .a(_al_u850_o),
    .b(\PWM3/FreCnt [2]),
    .c(\PWM3/FreCnt [20]),
    .d(\PWM3/FreCnt [21]),
    .e(\PWM3/FreCnt [22]),
    .o(_al_u851_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u852 (
    .a(_al_u847_o),
    .b(_al_u849_o),
    .c(_al_u851_o),
    .o(\PWM3/n0_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u853 (
    .a(\PWM3/n0_lutinv ),
    .b(\PWM3/stopreq ),
    .o(\PWM3/n1 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u854 (
    .a(\PWM3/n0_lutinv ),
    .b(\PWM3/n11 ),
    .o(\PWM3/mux3_b0_sel_is_3_o ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u855 (
    .a(\PWM3/n0_lutinv ),
    .b(\PWM3/n12 [9]),
    .c(freq3[9]),
    .o(\PWM3/n13 [9]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u856 (
    .a(\PWM3/n0_lutinv ),
    .b(\PWM3/n12 [8]),
    .c(freq3[8]),
    .o(\PWM3/n13 [8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u857 (
    .a(\PWM3/n0_lutinv ),
    .b(\PWM3/n12 [7]),
    .c(freq3[7]),
    .o(\PWM3/n13 [7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u858 (
    .a(\PWM3/n0_lutinv ),
    .b(\PWM3/n12 [6]),
    .c(freq3[6]),
    .o(\PWM3/n13 [6]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u859 (
    .a(\PWM3/n0_lutinv ),
    .b(\PWM3/n12 [5]),
    .c(freq3[5]),
    .o(\PWM3/n13 [5]));
  EF2_PHY_PAD #(
    //.LOCATION("P58"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u86 (
    .ipad(limit_l[3]),
    .di(limit_l_pad[3]));  // CPLD_SOC_AHB_TOP.v(5)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u860 (
    .a(\PWM3/n0_lutinv ),
    .b(\PWM3/n12 [4]),
    .c(freq3[4]),
    .o(\PWM3/n13 [4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u861 (
    .a(\PWM3/n0_lutinv ),
    .b(\PWM3/n12 [3]),
    .c(freq3[3]),
    .o(\PWM3/n13 [3]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u862 (
    .a(\PWM3/n0_lutinv ),
    .b(\PWM3/n12 [26]),
    .c(freq3[26]),
    .o(\PWM3/n13 [26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u863 (
    .a(\PWM3/n0_lutinv ),
    .b(\PWM3/n12 [25]),
    .c(freq3[25]),
    .o(\PWM3/n13 [25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u864 (
    .a(\PWM3/n0_lutinv ),
    .b(\PWM3/n12 [24]),
    .c(freq3[24]),
    .o(\PWM3/n13 [24]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u865 (
    .a(\PWM3/n0_lutinv ),
    .b(\PWM3/n12 [23]),
    .c(freq3[23]),
    .o(\PWM3/n13 [23]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u866 (
    .a(\PWM3/n0_lutinv ),
    .b(\PWM3/n12 [22]),
    .c(freq3[22]),
    .o(\PWM3/n13 [22]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u867 (
    .a(\PWM3/n0_lutinv ),
    .b(\PWM3/n12 [21]),
    .c(freq3[21]),
    .o(\PWM3/n13 [21]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u868 (
    .a(\PWM3/n0_lutinv ),
    .b(\PWM3/n12 [20]),
    .c(freq3[20]),
    .o(\PWM3/n13 [20]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u869 (
    .a(\PWM3/n0_lutinv ),
    .b(\PWM3/n12 [2]),
    .c(freq3[2]),
    .o(\PWM3/n13 [2]));
  EF2_PHY_PAD #(
    //.LOCATION("P56"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u87 (
    .ipad(limit_l[2]),
    .di(limit_l_pad[2]));  // CPLD_SOC_AHB_TOP.v(5)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u870 (
    .a(\PWM3/n0_lutinv ),
    .b(\PWM3/n12 [19]),
    .c(freq3[19]),
    .o(\PWM3/n13 [19]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u871 (
    .a(\PWM3/n0_lutinv ),
    .b(\PWM3/n12 [18]),
    .c(freq3[18]),
    .o(\PWM3/n13 [18]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u872 (
    .a(\PWM3/n0_lutinv ),
    .b(\PWM3/n12 [17]),
    .c(freq3[17]),
    .o(\PWM3/n13 [17]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u873 (
    .a(\PWM3/n0_lutinv ),
    .b(\PWM3/n12 [16]),
    .c(freq3[16]),
    .o(\PWM3/n13 [16]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u874 (
    .a(\PWM3/n0_lutinv ),
    .b(\PWM3/n12 [15]),
    .c(freq3[15]),
    .o(\PWM3/n13 [15]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u875 (
    .a(\PWM3/n0_lutinv ),
    .b(\PWM3/n12 [14]),
    .c(freq3[14]),
    .o(\PWM3/n13 [14]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u876 (
    .a(\PWM3/n0_lutinv ),
    .b(\PWM3/n12 [13]),
    .c(freq3[13]),
    .o(\PWM3/n13 [13]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u877 (
    .a(\PWM3/n0_lutinv ),
    .b(\PWM3/n12 [12]),
    .c(freq3[12]),
    .o(\PWM3/n13 [12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u878 (
    .a(\PWM3/n0_lutinv ),
    .b(\PWM3/n12 [11]),
    .c(freq3[11]),
    .o(\PWM3/n13 [11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u879 (
    .a(\PWM3/n0_lutinv ),
    .b(\PWM3/n12 [10]),
    .c(freq3[10]),
    .o(\PWM3/n13 [10]));
  EF2_PHY_PAD #(
    //.LOCATION("P50"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u88 (
    .ipad(limit_l[1]),
    .di(limit_l_pad[1]));  // CPLD_SOC_AHB_TOP.v(5)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u880 (
    .a(\PWM3/n0_lutinv ),
    .b(\PWM3/n12 [1]),
    .c(freq3[1]),
    .o(\PWM3/n13 [1]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u881 (
    .a(\PWM3/n0_lutinv ),
    .b(\PWM3/n12 [0]),
    .c(freq3[0]),
    .o(\PWM3/n13 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u882 (
    .a(\PWM4/FreCnt [23]),
    .b(\PWM4/FreCnt [24]),
    .c(\PWM4/FreCnt [25]),
    .d(\PWM4/FreCnt [26]),
    .o(_al_u882_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u883 (
    .a(_al_u882_o),
    .b(\PWM4/FreCnt [3]),
    .c(\PWM4/FreCnt [4]),
    .d(\PWM4/FreCnt [5]),
    .e(\PWM4/FreCnt [6]),
    .o(_al_u883_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u884 (
    .a(_al_u883_o),
    .b(\PWM4/FreCnt [7]),
    .c(\PWM4/FreCnt [8]),
    .d(\PWM4/FreCnt [9]),
    .o(_al_u884_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u885 (
    .a(\PWM4/FreCnt [0]),
    .b(\PWM4/FreCnt [1]),
    .c(\PWM4/FreCnt [10]),
    .d(\PWM4/FreCnt [11]),
    .o(_al_u885_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u886 (
    .a(_al_u885_o),
    .b(\PWM4/FreCnt [12]),
    .c(\PWM4/FreCnt [13]),
    .d(\PWM4/FreCnt [14]),
    .e(\PWM4/FreCnt [15]),
    .o(_al_u886_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u887 (
    .a(\PWM4/FreCnt [16]),
    .b(\PWM4/FreCnt [17]),
    .c(\PWM4/FreCnt [18]),
    .d(\PWM4/FreCnt [19]),
    .o(_al_u887_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u888 (
    .a(_al_u887_o),
    .b(\PWM4/FreCnt [2]),
    .c(\PWM4/FreCnt [20]),
    .d(\PWM4/FreCnt [21]),
    .e(\PWM4/FreCnt [22]),
    .o(_al_u888_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u889 (
    .a(_al_u884_o),
    .b(_al_u886_o),
    .c(_al_u888_o),
    .o(\PWM4/n0_lutinv ));
  EF2_PHY_PAD #(
    //.LOCATION("P41"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u89 (
    .ipad(limit_l[0]),
    .di(limit_l_pad[0]));  // CPLD_SOC_AHB_TOP.v(5)
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u890 (
    .a(\PWM4/n0_lutinv ),
    .b(\PWM4/stopreq ),
    .o(\PWM4/n1 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u891 (
    .a(\PWM4/n0_lutinv ),
    .b(\PWM4/n11 ),
    .o(\PWM4/mux3_b0_sel_is_3_o ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u892 (
    .a(\PWM4/n0_lutinv ),
    .b(\PWM4/n12 [9]),
    .c(freq4[9]),
    .o(\PWM4/n13 [9]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u893 (
    .a(\PWM4/n0_lutinv ),
    .b(\PWM4/n12 [8]),
    .c(freq4[8]),
    .o(\PWM4/n13 [8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u894 (
    .a(\PWM4/n0_lutinv ),
    .b(\PWM4/n12 [7]),
    .c(freq4[7]),
    .o(\PWM4/n13 [7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u895 (
    .a(\PWM4/n0_lutinv ),
    .b(\PWM4/n12 [6]),
    .c(freq4[6]),
    .o(\PWM4/n13 [6]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u896 (
    .a(\PWM4/n0_lutinv ),
    .b(\PWM4/n12 [5]),
    .c(freq4[5]),
    .o(\PWM4/n13 [5]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u897 (
    .a(\PWM4/n0_lutinv ),
    .b(\PWM4/n12 [4]),
    .c(freq4[4]),
    .o(\PWM4/n13 [4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u898 (
    .a(\PWM4/n0_lutinv ),
    .b(\PWM4/n12 [3]),
    .c(freq4[3]),
    .o(\PWM4/n13 [3]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u899 (
    .a(\PWM4/n0_lutinv ),
    .b(\PWM4/n12 [26]),
    .c(freq4[26]),
    .o(\PWM4/n13 [26]));
  EF2_PHY_SPAD #(
    //.LOCATION("P95"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u90 (
    .ipad(limit_r[15]),
    .ts(1'b1),
    .di(limit_r_pad[15]));  // CPLD_SOC_AHB_TOP.v(6)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u900 (
    .a(\PWM4/n0_lutinv ),
    .b(\PWM4/n12 [25]),
    .c(freq4[25]),
    .o(\PWM4/n13 [25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u901 (
    .a(\PWM4/n0_lutinv ),
    .b(\PWM4/n12 [24]),
    .c(freq4[24]),
    .o(\PWM4/n13 [24]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u902 (
    .a(\PWM4/n0_lutinv ),
    .b(\PWM4/n12 [23]),
    .c(freq4[23]),
    .o(\PWM4/n13 [23]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u903 (
    .a(\PWM4/n0_lutinv ),
    .b(\PWM4/n12 [22]),
    .c(freq4[22]),
    .o(\PWM4/n13 [22]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u904 (
    .a(\PWM4/n0_lutinv ),
    .b(\PWM4/n12 [21]),
    .c(freq4[21]),
    .o(\PWM4/n13 [21]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u905 (
    .a(\PWM4/n0_lutinv ),
    .b(\PWM4/n12 [20]),
    .c(freq4[20]),
    .o(\PWM4/n13 [20]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u906 (
    .a(\PWM4/n0_lutinv ),
    .b(\PWM4/n12 [2]),
    .c(freq4[2]),
    .o(\PWM4/n13 [2]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u907 (
    .a(\PWM4/n0_lutinv ),
    .b(\PWM4/n12 [19]),
    .c(freq4[19]),
    .o(\PWM4/n13 [19]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u908 (
    .a(\PWM4/n0_lutinv ),
    .b(\PWM4/n12 [18]),
    .c(freq4[18]),
    .o(\PWM4/n13 [18]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u909 (
    .a(\PWM4/n0_lutinv ),
    .b(\PWM4/n12 [17]),
    .c(freq4[17]),
    .o(\PWM4/n13 [17]));
  EF2_PHY_SPAD #(
    //.LOCATION("P81"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u91 (
    .ipad(limit_r[14]),
    .ts(1'b1),
    .di(limit_r_pad[14]));  // CPLD_SOC_AHB_TOP.v(6)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u910 (
    .a(\PWM4/n0_lutinv ),
    .b(\PWM4/n12 [16]),
    .c(freq4[16]),
    .o(\PWM4/n13 [16]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u911 (
    .a(\PWM4/n0_lutinv ),
    .b(\PWM4/n12 [15]),
    .c(freq4[15]),
    .o(\PWM4/n13 [15]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u912 (
    .a(\PWM4/n0_lutinv ),
    .b(\PWM4/n12 [14]),
    .c(freq4[14]),
    .o(\PWM4/n13 [14]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u913 (
    .a(\PWM4/n0_lutinv ),
    .b(\PWM4/n12 [13]),
    .c(freq4[13]),
    .o(\PWM4/n13 [13]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u914 (
    .a(\PWM4/n0_lutinv ),
    .b(\PWM4/n12 [12]),
    .c(freq4[12]),
    .o(\PWM4/n13 [12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u915 (
    .a(\PWM4/n0_lutinv ),
    .b(\PWM4/n12 [11]),
    .c(freq4[11]),
    .o(\PWM4/n13 [11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u916 (
    .a(\PWM4/n0_lutinv ),
    .b(\PWM4/n12 [10]),
    .c(freq4[10]),
    .o(\PWM4/n13 [10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u917 (
    .a(\PWM4/n0_lutinv ),
    .b(\PWM4/n12 [1]),
    .c(freq4[1]),
    .o(\PWM4/n13 [1]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u918 (
    .a(\PWM4/n0_lutinv ),
    .b(\PWM4/n12 [0]),
    .c(freq4[0]),
    .o(\PWM4/n13 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u919 (
    .a(\PWM5/FreCnt [23]),
    .b(\PWM5/FreCnt [24]),
    .c(\PWM5/FreCnt [25]),
    .d(\PWM5/FreCnt [26]),
    .o(_al_u919_o));
  EF2_PHY_SPAD #(
    //.LOCATION("P3"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u92 (
    .ipad(limit_r[13]),
    .ts(1'b1),
    .di(limit_r_pad[13]));  // CPLD_SOC_AHB_TOP.v(6)
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u920 (
    .a(_al_u919_o),
    .b(\PWM5/FreCnt [3]),
    .c(\PWM5/FreCnt [4]),
    .d(\PWM5/FreCnt [5]),
    .e(\PWM5/FreCnt [6]),
    .o(_al_u920_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u921 (
    .a(_al_u920_o),
    .b(\PWM5/FreCnt [7]),
    .c(\PWM5/FreCnt [8]),
    .d(\PWM5/FreCnt [9]),
    .o(_al_u921_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u922 (
    .a(\PWM5/FreCnt [0]),
    .b(\PWM5/FreCnt [1]),
    .c(\PWM5/FreCnt [10]),
    .d(\PWM5/FreCnt [11]),
    .o(_al_u922_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u923 (
    .a(_al_u922_o),
    .b(\PWM5/FreCnt [12]),
    .c(\PWM5/FreCnt [13]),
    .d(\PWM5/FreCnt [14]),
    .e(\PWM5/FreCnt [15]),
    .o(_al_u923_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u924 (
    .a(\PWM5/FreCnt [16]),
    .b(\PWM5/FreCnt [17]),
    .c(\PWM5/FreCnt [18]),
    .d(\PWM5/FreCnt [19]),
    .o(_al_u924_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u925 (
    .a(_al_u924_o),
    .b(\PWM5/FreCnt [2]),
    .c(\PWM5/FreCnt [20]),
    .d(\PWM5/FreCnt [21]),
    .e(\PWM5/FreCnt [22]),
    .o(_al_u925_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u926 (
    .a(_al_u921_o),
    .b(_al_u923_o),
    .c(_al_u925_o),
    .o(\PWM5/n0_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u927 (
    .a(\PWM5/n0_lutinv ),
    .b(\PWM5/stopreq ),
    .o(\PWM5/n1 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u928 (
    .a(\PWM5/n0_lutinv ),
    .b(\PWM5/n11 ),
    .o(\PWM5/mux3_b0_sel_is_3_o ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u929 (
    .a(\PWM5/n0_lutinv ),
    .b(\PWM5/n12 [9]),
    .c(freq5[9]),
    .o(\PWM5/n13 [9]));
  EF2_PHY_SPAD #(
    //.LOCATION("P5"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u93 (
    .ipad(limit_r[12]),
    .ts(1'b1),
    .di(limit_r_pad[12]));  // CPLD_SOC_AHB_TOP.v(6)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u930 (
    .a(\PWM5/n0_lutinv ),
    .b(\PWM5/n12 [8]),
    .c(freq5[8]),
    .o(\PWM5/n13 [8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u931 (
    .a(\PWM5/n0_lutinv ),
    .b(\PWM5/n12 [7]),
    .c(freq5[7]),
    .o(\PWM5/n13 [7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u932 (
    .a(\PWM5/n0_lutinv ),
    .b(\PWM5/n12 [6]),
    .c(freq5[6]),
    .o(\PWM5/n13 [6]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u933 (
    .a(\PWM5/n0_lutinv ),
    .b(\PWM5/n12 [5]),
    .c(freq5[5]),
    .o(\PWM5/n13 [5]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u934 (
    .a(\PWM5/n0_lutinv ),
    .b(\PWM5/n12 [4]),
    .c(freq5[4]),
    .o(\PWM5/n13 [4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u935 (
    .a(\PWM5/n0_lutinv ),
    .b(\PWM5/n12 [3]),
    .c(freq5[3]),
    .o(\PWM5/n13 [3]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u936 (
    .a(\PWM5/n0_lutinv ),
    .b(\PWM5/n12 [26]),
    .c(freq5[26]),
    .o(\PWM5/n13 [26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u937 (
    .a(\PWM5/n0_lutinv ),
    .b(\PWM5/n12 [25]),
    .c(freq5[25]),
    .o(\PWM5/n13 [25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u938 (
    .a(\PWM5/n0_lutinv ),
    .b(\PWM5/n12 [24]),
    .c(freq5[24]),
    .o(\PWM5/n13 [24]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u939 (
    .a(\PWM5/n0_lutinv ),
    .b(\PWM5/n12 [23]),
    .c(freq5[23]),
    .o(\PWM5/n13 [23]));
  EF2_PHY_PAD #(
    //.LOCATION("P68"),
    //.PCICLAMP("ON"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u94 (
    .ipad(limit_r[11]),
    .di(limit_r_pad[11]));  // CPLD_SOC_AHB_TOP.v(6)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u940 (
    .a(\PWM5/n0_lutinv ),
    .b(\PWM5/n12 [22]),
    .c(freq5[22]),
    .o(\PWM5/n13 [22]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u941 (
    .a(\PWM5/n0_lutinv ),
    .b(\PWM5/n12 [21]),
    .c(freq5[21]),
    .o(\PWM5/n13 [21]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u942 (
    .a(\PWM5/n0_lutinv ),
    .b(\PWM5/n12 [20]),
    .c(freq5[20]),
    .o(\PWM5/n13 [20]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u943 (
    .a(\PWM5/n0_lutinv ),
    .b(\PWM5/n12 [2]),
    .c(freq5[2]),
    .o(\PWM5/n13 [2]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u944 (
    .a(\PWM5/n0_lutinv ),
    .b(\PWM5/n12 [19]),
    .c(freq5[19]),
    .o(\PWM5/n13 [19]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u945 (
    .a(\PWM5/n0_lutinv ),
    .b(\PWM5/n12 [18]),
    .c(freq5[18]),
    .o(\PWM5/n13 [18]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u946 (
    .a(\PWM5/n0_lutinv ),
    .b(\PWM5/n12 [17]),
    .c(freq5[17]),
    .o(\PWM5/n13 [17]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u947 (
    .a(\PWM5/n0_lutinv ),
    .b(\PWM5/n12 [16]),
    .c(freq5[16]),
    .o(\PWM5/n13 [16]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u948 (
    .a(\PWM5/n0_lutinv ),
    .b(\PWM5/n12 [15]),
    .c(freq5[15]),
    .o(\PWM5/n13 [15]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u949 (
    .a(\PWM5/n0_lutinv ),
    .b(\PWM5/n12 [14]),
    .c(freq5[14]),
    .o(\PWM5/n13 [14]));
  EF2_PHY_SPAD #(
    //.LOCATION("P35"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u95 (
    .ipad(limit_r[10]),
    .ts(1'b1),
    .di(limit_r_pad[10]));  // CPLD_SOC_AHB_TOP.v(6)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u950 (
    .a(\PWM5/n0_lutinv ),
    .b(\PWM5/n12 [13]),
    .c(freq5[13]),
    .o(\PWM5/n13 [13]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u951 (
    .a(\PWM5/n0_lutinv ),
    .b(\PWM5/n12 [12]),
    .c(freq5[12]),
    .o(\PWM5/n13 [12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u952 (
    .a(\PWM5/n0_lutinv ),
    .b(\PWM5/n12 [11]),
    .c(freq5[11]),
    .o(\PWM5/n13 [11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u953 (
    .a(\PWM5/n0_lutinv ),
    .b(\PWM5/n12 [10]),
    .c(freq5[10]),
    .o(\PWM5/n13 [10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u954 (
    .a(\PWM5/n0_lutinv ),
    .b(\PWM5/n12 [1]),
    .c(freq5[1]),
    .o(\PWM5/n13 [1]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u955 (
    .a(\PWM5/n0_lutinv ),
    .b(\PWM5/n12 [0]),
    .c(freq5[0]),
    .o(\PWM5/n13 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u956 (
    .a(\PWM6/FreCnt [23]),
    .b(\PWM6/FreCnt [24]),
    .c(\PWM6/FreCnt [25]),
    .d(\PWM6/FreCnt [26]),
    .o(_al_u956_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u957 (
    .a(_al_u956_o),
    .b(\PWM6/FreCnt [3]),
    .c(\PWM6/FreCnt [4]),
    .d(\PWM6/FreCnt [5]),
    .e(\PWM6/FreCnt [6]),
    .o(_al_u957_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u958 (
    .a(_al_u957_o),
    .b(\PWM6/FreCnt [7]),
    .c(\PWM6/FreCnt [8]),
    .d(\PWM6/FreCnt [9]),
    .o(_al_u958_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u959 (
    .a(\PWM6/FreCnt [0]),
    .b(\PWM6/FreCnt [1]),
    .c(\PWM6/FreCnt [10]),
    .d(\PWM6/FreCnt [11]),
    .o(_al_u959_o));
  EF2_PHY_SPAD #(
    //.LOCATION("P94"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u96 (
    .ipad(limit_r[9]),
    .ts(1'b1),
    .di(limit_r_pad[9]));  // CPLD_SOC_AHB_TOP.v(6)
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u960 (
    .a(_al_u959_o),
    .b(\PWM6/FreCnt [12]),
    .c(\PWM6/FreCnt [13]),
    .d(\PWM6/FreCnt [14]),
    .e(\PWM6/FreCnt [15]),
    .o(_al_u960_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u961 (
    .a(\PWM6/FreCnt [16]),
    .b(\PWM6/FreCnt [17]),
    .c(\PWM6/FreCnt [18]),
    .d(\PWM6/FreCnt [19]),
    .o(_al_u961_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u962 (
    .a(_al_u961_o),
    .b(\PWM6/FreCnt [2]),
    .c(\PWM6/FreCnt [20]),
    .d(\PWM6/FreCnt [21]),
    .e(\PWM6/FreCnt [22]),
    .o(_al_u962_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u963 (
    .a(_al_u958_o),
    .b(_al_u960_o),
    .c(_al_u962_o),
    .o(\PWM6/n0_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u964 (
    .a(\PWM6/n0_lutinv ),
    .b(\PWM6/stopreq ),
    .o(\PWM6/n1 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u965 (
    .a(\PWM6/n0_lutinv ),
    .b(\PWM6/n11 ),
    .o(\PWM6/mux3_b0_sel_is_3_o ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u966 (
    .a(\PWM6/n0_lutinv ),
    .b(\PWM6/n12 [9]),
    .c(freq6[9]),
    .o(\PWM6/n13 [9]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u967 (
    .a(\PWM6/n0_lutinv ),
    .b(\PWM6/n12 [8]),
    .c(freq6[8]),
    .o(\PWM6/n13 [8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u968 (
    .a(\PWM6/n0_lutinv ),
    .b(\PWM6/n12 [7]),
    .c(freq6[7]),
    .o(\PWM6/n13 [7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u969 (
    .a(\PWM6/n0_lutinv ),
    .b(\PWM6/n12 [6]),
    .c(freq6[6]),
    .o(\PWM6/n13 [6]));
  EF2_PHY_SPAD #(
    //.LOCATION("P86"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u97 (
    .ipad(limit_r[8]),
    .ts(1'b1),
    .di(limit_r_pad[8]));  // CPLD_SOC_AHB_TOP.v(6)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u970 (
    .a(\PWM6/n0_lutinv ),
    .b(\PWM6/n12 [5]),
    .c(freq6[5]),
    .o(\PWM6/n13 [5]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u971 (
    .a(\PWM6/n0_lutinv ),
    .b(\PWM6/n12 [4]),
    .c(freq6[4]),
    .o(\PWM6/n13 [4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u972 (
    .a(\PWM6/n0_lutinv ),
    .b(\PWM6/n12 [3]),
    .c(freq6[3]),
    .o(\PWM6/n13 [3]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u973 (
    .a(\PWM6/n0_lutinv ),
    .b(\PWM6/n12 [26]),
    .c(freq6[26]),
    .o(\PWM6/n13 [26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u974 (
    .a(\PWM6/n0_lutinv ),
    .b(\PWM6/n12 [25]),
    .c(freq6[25]),
    .o(\PWM6/n13 [25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u975 (
    .a(\PWM6/n0_lutinv ),
    .b(\PWM6/n12 [24]),
    .c(freq6[24]),
    .o(\PWM6/n13 [24]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u976 (
    .a(\PWM6/n0_lutinv ),
    .b(\PWM6/n12 [23]),
    .c(freq6[23]),
    .o(\PWM6/n13 [23]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u977 (
    .a(\PWM6/n0_lutinv ),
    .b(\PWM6/n12 [22]),
    .c(freq6[22]),
    .o(\PWM6/n13 [22]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u978 (
    .a(\PWM6/n0_lutinv ),
    .b(\PWM6/n12 [21]),
    .c(freq6[21]),
    .o(\PWM6/n13 [21]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u979 (
    .a(\PWM6/n0_lutinv ),
    .b(\PWM6/n12 [20]),
    .c(freq6[20]),
    .o(\PWM6/n13 [20]));
  EF2_PHY_SPAD #(
    //.LOCATION("P82"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u98 (
    .ipad(limit_r[7]),
    .ts(1'b1),
    .di(limit_r_pad[7]));  // CPLD_SOC_AHB_TOP.v(6)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u980 (
    .a(\PWM6/n0_lutinv ),
    .b(\PWM6/n12 [2]),
    .c(freq6[2]),
    .o(\PWM6/n13 [2]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u981 (
    .a(\PWM6/n0_lutinv ),
    .b(\PWM6/n12 [19]),
    .c(freq6[19]),
    .o(\PWM6/n13 [19]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u982 (
    .a(\PWM6/n0_lutinv ),
    .b(\PWM6/n12 [18]),
    .c(freq6[18]),
    .o(\PWM6/n13 [18]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u983 (
    .a(\PWM6/n0_lutinv ),
    .b(\PWM6/n12 [17]),
    .c(freq6[17]),
    .o(\PWM6/n13 [17]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u984 (
    .a(\PWM6/n0_lutinv ),
    .b(\PWM6/n12 [16]),
    .c(freq6[16]),
    .o(\PWM6/n13 [16]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u985 (
    .a(\PWM6/n0_lutinv ),
    .b(\PWM6/n12 [15]),
    .c(freq6[15]),
    .o(\PWM6/n13 [15]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u986 (
    .a(\PWM6/n0_lutinv ),
    .b(\PWM6/n12 [14]),
    .c(freq6[14]),
    .o(\PWM6/n13 [14]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u987 (
    .a(\PWM6/n0_lutinv ),
    .b(\PWM6/n12 [13]),
    .c(freq6[13]),
    .o(\PWM6/n13 [13]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u988 (
    .a(\PWM6/n0_lutinv ),
    .b(\PWM6/n12 [12]),
    .c(freq6[12]),
    .o(\PWM6/n13 [12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u989 (
    .a(\PWM6/n0_lutinv ),
    .b(\PWM6/n12 [11]),
    .c(freq6[11]),
    .o(\PWM6/n13 [11]));
  EF2_PHY_SPAD #(
    //.LOCATION("P4"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("TS"))
    _al_u99 (
    .ipad(limit_r[6]),
    .ts(1'b1),
    .di(limit_r_pad[6]));  // CPLD_SOC_AHB_TOP.v(6)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u990 (
    .a(\PWM6/n0_lutinv ),
    .b(\PWM6/n12 [10]),
    .c(freq6[10]),
    .o(\PWM6/n13 [10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u991 (
    .a(\PWM6/n0_lutinv ),
    .b(\PWM6/n12 [1]),
    .c(freq6[1]),
    .o(\PWM6/n13 [1]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u992 (
    .a(\PWM6/n0_lutinv ),
    .b(\PWM6/n12 [0]),
    .c(freq6[0]),
    .o(\PWM6/n13 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u993 (
    .a(\PWM7/FreCnt [23]),
    .b(\PWM7/FreCnt [24]),
    .c(\PWM7/FreCnt [25]),
    .d(\PWM7/FreCnt [26]),
    .o(_al_u993_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u994 (
    .a(_al_u993_o),
    .b(\PWM7/FreCnt [3]),
    .c(\PWM7/FreCnt [4]),
    .d(\PWM7/FreCnt [5]),
    .e(\PWM7/FreCnt [6]),
    .o(_al_u994_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u995 (
    .a(_al_u994_o),
    .b(\PWM7/FreCnt [7]),
    .c(\PWM7/FreCnt [8]),
    .d(\PWM7/FreCnt [9]),
    .o(_al_u995_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u996 (
    .a(\PWM7/FreCnt [0]),
    .b(\PWM7/FreCnt [1]),
    .c(\PWM7/FreCnt [10]),
    .d(\PWM7/FreCnt [11]),
    .o(_al_u996_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u997 (
    .a(_al_u996_o),
    .b(\PWM7/FreCnt [12]),
    .c(\PWM7/FreCnt [13]),
    .d(\PWM7/FreCnt [14]),
    .e(\PWM7/FreCnt [15]),
    .o(_al_u997_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u998 (
    .a(\PWM7/FreCnt [16]),
    .b(\PWM7/FreCnt [17]),
    .c(\PWM7/FreCnt [18]),
    .d(\PWM7/FreCnt [19]),
    .o(_al_u998_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u999 (
    .a(_al_u998_o),
    .b(\PWM7/FreCnt [2]),
    .c(\PWM7/FreCnt [20]),
    .d(\PWM7/FreCnt [21]),
    .e(\PWM7/FreCnt [22]),
    .o(_al_u999_o));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    _bufkeep_clk100m (
    .i(clk100m_keep),
    .o(clk100m));  // CPLD_SOC_AHB_TOP.v(13)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u0  (
    .a(timer[0]),
    .b(1'b1),
    .c(\add0/c0 ),
    .o({\add0/c1 ,n2[0]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u1  (
    .a(timer[1]),
    .b(1'b0),
    .c(\add0/c1 ),
    .o({\add0/c2 ,n2[1]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u10  (
    .a(timer[10]),
    .b(1'b0),
    .c(\add0/c10 ),
    .o({\add0/c11 ,n2[10]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u11  (
    .a(timer[11]),
    .b(1'b0),
    .c(\add0/c11 ),
    .o({\add0/c12 ,n2[11]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u12  (
    .a(timer[12]),
    .b(1'b0),
    .c(\add0/c12 ),
    .o({\add0/c13 ,n2[12]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u13  (
    .a(timer[13]),
    .b(1'b0),
    .c(\add0/c13 ),
    .o({\add0/c14 ,n2[13]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u14  (
    .a(timer[14]),
    .b(1'b0),
    .c(\add0/c14 ),
    .o({\add0/c15 ,n2[14]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u15  (
    .a(timer[15]),
    .b(1'b0),
    .c(\add0/c15 ),
    .o({\add0/c16 ,n2[15]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u16  (
    .a(timer[16]),
    .b(1'b0),
    .c(\add0/c16 ),
    .o({\add0/c17 ,n2[16]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u17  (
    .a(timer[17]),
    .b(1'b0),
    .c(\add0/c17 ),
    .o({\add0/c18 ,n2[17]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u18  (
    .a(timer[18]),
    .b(1'b0),
    .c(\add0/c18 ),
    .o({\add0/c19 ,n2[18]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u19  (
    .a(timer[19]),
    .b(1'b0),
    .c(\add0/c19 ),
    .o({\add0/c20 ,n2[19]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u2  (
    .a(timer[2]),
    .b(1'b0),
    .c(\add0/c2 ),
    .o({\add0/c3 ,n2[2]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u20  (
    .a(timer[20]),
    .b(1'b0),
    .c(\add0/c20 ),
    .o({\add0/c21 ,n2[20]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u21  (
    .a(timer[21]),
    .b(1'b0),
    .c(\add0/c21 ),
    .o({\add0/c22 ,n2[21]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u22  (
    .a(timer[22]),
    .b(1'b0),
    .c(\add0/c22 ),
    .o({\add0/c23 ,n2[22]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u23  (
    .a(timer[23]),
    .b(1'b0),
    .c(\add0/c23 ),
    .o({\add0/c24 ,n2[23]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u24  (
    .a(timer[24]),
    .b(1'b0),
    .c(\add0/c24 ),
    .o({\add0/c25 ,n2[24]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u25  (
    .a(timer[25]),
    .b(1'b0),
    .c(\add0/c25 ),
    .o({\add0/c26 ,n2[25]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u26  (
    .a(timer[26]),
    .b(1'b0),
    .c(\add0/c26 ),
    .o({\add0/c27 ,n2[26]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u27  (
    .a(timer[27]),
    .b(1'b0),
    .c(\add0/c27 ),
    .o({\add0/c28 ,n2[27]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u28  (
    .a(timer[28]),
    .b(1'b0),
    .c(\add0/c28 ),
    .o({\add0/c29 ,n2[28]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u29  (
    .a(timer[29]),
    .b(1'b0),
    .c(\add0/c29 ),
    .o({\add0/c30 ,n2[29]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u3  (
    .a(timer[3]),
    .b(1'b0),
    .c(\add0/c3 ),
    .o({\add0/c4 ,n2[3]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u30  (
    .a(timer[30]),
    .b(1'b0),
    .c(\add0/c30 ),
    .o({\add0/c31 ,n2[30]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u31  (
    .a(timer[31]),
    .b(1'b0),
    .c(\add0/c31 ),
    .o({open_n1866,n2[31]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u4  (
    .a(timer[4]),
    .b(1'b0),
    .c(\add0/c4 ),
    .o({\add0/c5 ,n2[4]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u5  (
    .a(timer[5]),
    .b(1'b0),
    .c(\add0/c5 ),
    .o({\add0/c6 ,n2[5]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u6  (
    .a(timer[6]),
    .b(1'b0),
    .c(\add0/c6 ),
    .o({\add0/c7 ,n2[6]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u7  (
    .a(timer[7]),
    .b(1'b0),
    .c(\add0/c7 ),
    .o({\add0/c8 ,n2[7]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u8  (
    .a(timer[8]),
    .b(1'b0),
    .c(\add0/c8 ),
    .o({\add0/c9 ,n2[8]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \add0/u9  (
    .a(timer[9]),
    .b(1'b0),
    .c(\add0/c9 ),
    .o({\add0/c10 ,n2[9]}));
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \add0/ucin  (
    .a(1'b0),
    .o({\add0/c0 ,open_n1869}));
  EF2_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  reg_ar_as_w1 reg0_b0 (
    .clk(clk25m),
    .d(n3[0]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(timer[0]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b1 (
    .clk(clk25m),
    .d(n3[1]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(timer[1]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b10 (
    .clk(clk25m),
    .d(n3[10]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(timer[10]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b11 (
    .clk(clk25m),
    .d(n3[11]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(timer[11]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b12 (
    .clk(clk25m),
    .d(n3[12]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(timer[12]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b13 (
    .clk(clk25m),
    .d(n3[13]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(timer[13]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b14 (
    .clk(clk25m),
    .d(n3[14]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(timer[14]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b15 (
    .clk(clk25m),
    .d(n3[15]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(timer[15]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b16 (
    .clk(clk25m),
    .d(n3[16]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(timer[16]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b17 (
    .clk(clk25m),
    .d(n3[17]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(timer[17]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b18 (
    .clk(clk25m),
    .d(n3[18]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(timer[18]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b19 (
    .clk(clk25m),
    .d(n3[19]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(timer[19]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b2 (
    .clk(clk25m),
    .d(n3[2]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(timer[2]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b20 (
    .clk(clk25m),
    .d(n3[20]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(timer[20]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b21 (
    .clk(clk25m),
    .d(n3[21]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(timer[21]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b22 (
    .clk(clk25m),
    .d(n3[22]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(timer[22]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b23 (
    .clk(clk25m),
    .d(n3[23]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(timer[23]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b24 (
    .clk(clk25m),
    .d(n3[24]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(timer[24]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b25 (
    .clk(clk25m),
    .d(n3[25]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(timer[25]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b26 (
    .clk(clk25m),
    .d(n3[26]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(timer[26]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b27 (
    .clk(clk25m),
    .d(n3[27]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(timer[27]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b28 (
    .clk(clk25m),
    .d(n3[28]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(timer[28]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b29 (
    .clk(clk25m),
    .d(n3[29]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(timer[29]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b3 (
    .clk(clk25m),
    .d(n3[3]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(timer[3]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b30 (
    .clk(clk25m),
    .d(n3[30]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(timer[30]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b31 (
    .clk(clk25m),
    .d(n3[31]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(timer[31]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b4 (
    .clk(clk25m),
    .d(n3[4]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(timer[4]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b5 (
    .clk(clk25m),
    .d(n3[5]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(timer[5]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b6 (
    .clk(clk25m),
    .d(n3[6]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(timer[6]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b7 (
    .clk(clk25m),
    .d(n3[7]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(timer[7]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b8 (
    .clk(clk25m),
    .d(n3[8]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(timer[8]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b9 (
    .clk(clk25m),
    .d(n3[9]),
    .en(1'b1),
    .reset(~rst_n_pad),
    .set(1'b0),
    .q(timer[9]));  // CPLD_SOC_AHB_TOP.v(35)
  EF2_PHY_SPAD #(
    //.CLKSRC("CLK"),
    //.LOCATION("P105"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("FAST"),
    .DO_DFFMODE("FF"),
    .DO_REGSET("SET"),
    .DRIVE("16"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .OUTCEMUX("CE"),
    .OUTCLKMUX("CLK"),
    .OUTRSTMUX("INV"),
    .SRMODE("ASYNC"),
    .TSMUX("INV"))
    reg1_b0_DO (
    .ce(_al_n1_en),
    .clk(clk25m),
    .do({open_n1917,n4_neg}),
    .rst(rst_n_pad),
    .ts(1'b1),
    .opad(ledout[0]));  // CPLD_SOC_AHB_TOP.v(49)
  reg_ar_as_w1 reg1_b1 (
    .clk(clk25m),
    .d(n10[1]),
    .en(1'b1),
    .reset(1'b0),
    .set(~rst_n_pad),
    .q(ledout_pad[1]));  // CPLD_SOC_AHB_TOP.v(49)
  reg_ar_as_w1 reg1_b2 (
    .clk(clk25m),
    .d(n10[2]),
    .en(1'b1),
    .reset(1'b0),
    .set(~rst_n_pad),
    .q(ledout_pad[2]));  // CPLD_SOC_AHB_TOP.v(49)
  reg_ar_as_w1 reg1_b3 (
    .clk(clk25m),
    .d(n10[3]),
    .en(1'b1),
    .reset(1'b0),
    .set(~rst_n_pad),
    .q(ledout_pad[3]));  // CPLD_SOC_AHB_TOP.v(49)

endmodule 

module reg_ar_as_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  parameter REGSET = "RESET";
  wire enout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_DFF #(
    .INI((REGSET == "SET") ? 1'b1 : 1'b0))
    u_seq0 (
    .clk(clk),
    .d(enout),
    .reset(reset),
    .set(set),
    .q(q));

endmodule 

module AL_BUFKEEP
  (
  i,
  o
  );

  input i;
  output o;

  parameter KEEP = "OUT";

  buf u1 (o, i);

endmodule 

module reg_sr_as_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  parameter REGSET = "RESET";
  wire enout;
  wire resetout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_MUX u_reset0 (
    .i0(enout),
    .i1(1'b0),
    .sel(reset),
    .o(resetout));
  AL_DFF #(
    .INI((REGSET == "SET") ? 1'b1 : 1'b0))
    u_seq0 (
    .clk(clk),
    .d(resetout),
    .reset(1'b0),
    .set(set),
    .q(q));

endmodule 

module reg_ar_ss_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  parameter REGSET = "RESET";
  wire enout;
  wire setout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_DFF #(
    .INI((REGSET == "SET") ? 1'b1 : 1'b0))
    u_seq0 (
    .clk(clk),
    .d(setout),
    .reset(reset),
    .set(1'b0),
    .q(q));
  AL_MUX u_set0 (
    .i0(enout),
    .i1(1'b1),
    .sel(set),
    .o(setout));

endmodule 

module AL_MUX
  (
  input i0,
  input i1,
  input sel,
  output o
  );

  wire not_sel, sel_i0, sel_i1;
  not u0 (not_sel, sel);
  and u1 (sel_i1, sel, i1);
  and u2 (sel_i0, not_sel, i0);
  or u3 (o, sel_i1, sel_i0);

endmodule

module AL_DFF
  (
  input reset,
  input set,
  input clk,
  input d,
  output reg q
  );

  parameter INI = 1'b0;

  always @(posedge reset or posedge set or posedge clk)
  begin
    if (reset)
      q <= 1'b0;
    else if (set)
      q <= 1'b1;
    else
      q <= d;
  end

endmodule

