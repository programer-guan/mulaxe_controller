// Verilog netlist created by TD v4.5.12562
// Thu Dec 19 17:41:47 2019

`timescale 1ns / 1ps
module CPLD_SOC_AHB_TOP  // CPLD_SOC_AHB_TOP.v(1)
  (
  clkin,
  limit_l,
  limit_r,
  rst_n,
  dir,
  gpio_out,
  ledout,
  pwm
  );

  input clkin;  // CPLD_SOC_AHB_TOP.v(3)
  input [15:0] limit_l;  // CPLD_SOC_AHB_TOP.v(5)
  input [15:0] limit_r;  // CPLD_SOC_AHB_TOP.v(6)
  input rst_n;  // CPLD_SOC_AHB_TOP.v(4)
  output [15:0] dir;  // CPLD_SOC_AHB_TOP.v(7)
  output [31:0] gpio_out;  // CPLD_SOC_AHB_TOP.v(8)
  output [3:0] ledout;  // CPLD_SOC_AHB_TOP.v(10)
  output [15:0] pwm;  // CPLD_SOC_AHB_TOP.v(7)

  wire [26:0] \PWM0/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWM0/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWM0/n12 ;
  wire [26:0] \PWM0/n13 ;
  wire [31:0] \PWM0/n22 ;
  wire [31:0] \PWM0/n23 ;
  wire [24:0] \PWM0/n26 ;
  wire [23:0] \PWM0/n27 ;
  wire [23:0] \PWM0/n29 ;
  wire [23:0] \PWM0/n31 ;
  wire [31:0] \PWM0/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWM1/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWM1/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWM1/n12 ;
  wire [26:0] \PWM1/n13 ;
  wire [31:0] \PWM1/n22 ;
  wire [31:0] \PWM1/n23 ;
  wire [24:0] \PWM1/n26 ;
  wire [23:0] \PWM1/n27 ;
  wire [23:0] \PWM1/n29 ;
  wire [23:0] \PWM1/n31 ;
  wire [31:0] \PWM1/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWM2/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWM2/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWM2/n12 ;
  wire [26:0] \PWM2/n13 ;
  wire [31:0] \PWM2/n22 ;
  wire [31:0] \PWM2/n23 ;
  wire [24:0] \PWM2/n26 ;
  wire [23:0] \PWM2/n27 ;
  wire [23:0] \PWM2/n29 ;
  wire [23:0] \PWM2/n31 ;
  wire [31:0] \PWM2/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWM3/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWM3/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWM3/n12 ;
  wire [26:0] \PWM3/n13 ;
  wire [31:0] \PWM3/n22 ;
  wire [31:0] \PWM3/n23 ;
  wire [24:0] \PWM3/n26 ;
  wire [23:0] \PWM3/n27 ;
  wire [23:0] \PWM3/n29 ;
  wire [23:0] \PWM3/n31 ;
  wire [31:0] \PWM3/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWM4/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWM4/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWM4/n12 ;
  wire [26:0] \PWM4/n13 ;
  wire [31:0] \PWM4/n22 ;
  wire [31:0] \PWM4/n23 ;
  wire [24:0] \PWM4/n26 ;
  wire [23:0] \PWM4/n27 ;
  wire [23:0] \PWM4/n29 ;
  wire [23:0] \PWM4/n31 ;
  wire [31:0] \PWM4/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWM5/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWM5/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWM5/n12 ;
  wire [26:0] \PWM5/n13 ;
  wire [31:0] \PWM5/n22 ;
  wire [31:0] \PWM5/n23 ;
  wire [24:0] \PWM5/n26 ;
  wire [23:0] \PWM5/n27 ;
  wire [23:0] \PWM5/n29 ;
  wire [23:0] \PWM5/n31 ;
  wire [31:0] \PWM5/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWM6/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWM6/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWM6/n12 ;
  wire [26:0] \PWM6/n13 ;
  wire [31:0] \PWM6/n22 ;
  wire [31:0] \PWM6/n23 ;
  wire [24:0] \PWM6/n26 ;
  wire [23:0] \PWM6/n27 ;
  wire [23:0] \PWM6/n29 ;
  wire [23:0] \PWM6/n31 ;
  wire [31:0] \PWM6/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWM7/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWM7/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWM7/n12 ;
  wire [26:0] \PWM7/n13 ;
  wire [31:0] \PWM7/n22 ;
  wire [31:0] \PWM7/n23 ;
  wire [24:0] \PWM7/n26 ;
  wire [23:0] \PWM7/n27 ;
  wire [23:0] \PWM7/n29 ;
  wire [23:0] \PWM7/n31 ;
  wire [31:0] \PWM7/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWM8/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWM8/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWM8/n12 ;
  wire [26:0] \PWM8/n13 ;
  wire [31:0] \PWM8/n22 ;
  wire [31:0] \PWM8/n23 ;
  wire [24:0] \PWM8/n26 ;
  wire [23:0] \PWM8/n27 ;
  wire [23:0] \PWM8/n29 ;
  wire [23:0] \PWM8/n31 ;
  wire [31:0] \PWM8/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWM9/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWM9/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWM9/n12 ;
  wire [26:0] \PWM9/n13 ;
  wire [31:0] \PWM9/n22 ;
  wire [31:0] \PWM9/n23 ;
  wire [24:0] \PWM9/n26 ;
  wire [23:0] \PWM9/n27 ;
  wire [23:0] \PWM9/n29 ;
  wire [23:0] \PWM9/n31 ;
  wire [31:0] \PWM9/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWMA/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWMA/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWMA/n12 ;
  wire [26:0] \PWMA/n13 ;
  wire [31:0] \PWMA/n22 ;
  wire [31:0] \PWMA/n23 ;
  wire [24:0] \PWMA/n26 ;
  wire [23:0] \PWMA/n27 ;
  wire [23:0] \PWMA/n29 ;
  wire [23:0] \PWMA/n31 ;
  wire [31:0] \PWMA/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWMB/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWMB/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWMB/n12 ;
  wire [26:0] \PWMB/n13 ;
  wire [31:0] \PWMB/n22 ;
  wire [31:0] \PWMB/n23 ;
  wire [24:0] \PWMB/n26 ;
  wire [23:0] \PWMB/n27 ;
  wire [23:0] \PWMB/n29 ;
  wire [23:0] \PWMB/n31 ;
  wire [31:0] \PWMB/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWMC/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWMC/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWMC/n12 ;
  wire [26:0] \PWMC/n13 ;
  wire [31:0] \PWMC/n22 ;
  wire [31:0] \PWMC/n23 ;
  wire [24:0] \PWMC/n26 ;
  wire [23:0] \PWMC/n27 ;
  wire [23:0] \PWMC/n29 ;
  wire [23:0] \PWMC/n31 ;
  wire [31:0] \PWMC/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWMD/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWMD/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWMD/n12 ;
  wire [26:0] \PWMD/n13 ;
  wire [31:0] \PWMD/n22 ;
  wire [31:0] \PWMD/n23 ;
  wire [24:0] \PWMD/n26 ;
  wire [23:0] \PWMD/n27 ;
  wire [23:0] \PWMD/n29 ;
  wire [23:0] \PWMD/n31 ;
  wire [31:0] \PWMD/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWME/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWME/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWME/n12 ;
  wire [26:0] \PWME/n13 ;
  wire [31:0] \PWME/n22 ;
  wire [31:0] \PWME/n23 ;
  wire [24:0] \PWME/n26 ;
  wire [23:0] \PWME/n27 ;
  wire [23:0] \PWME/n29 ;
  wire [23:0] \PWME/n31 ;
  wire [31:0] \PWME/pnumr ;  // src/OnePWM.v(47)
  wire [26:0] \PWMF/FreCnt ;  // src/OnePWM.v(13)
  wire [26:0] \PWMF/FreCntr ;  // src/OnePWM.v(13)
  wire [27:0] \PWMF/n12 ;
  wire [26:0] \PWMF/n13 ;
  wire [31:0] \PWMF/n22 ;
  wire [31:0] \PWMF/n23 ;
  wire [24:0] \PWMF/n26 ;
  wire [23:0] \PWMF/n27 ;
  wire [23:0] \PWMF/n29 ;
  wire [23:0] \PWMF/n31 ;
  wire [31:0] \PWMF/pnumr ;  // src/OnePWM.v(47)
  wire [31:0] \U_AHB/h2h_haddr ;  // src/AHB.v(23)
  wire [31:0] \U_AHB/h2h_haddrw ;  // src/AHB.v(16)
  wire [31:0] \U_AHB/h2h_hrdata ;  // src/AHB.v(18)
  wire [31:0] \U_AHB/h2h_hwdata ;  // src/AHB.v(17)
  wire [31:0] \U_AHB/n114 ;
  wire [31:0] \U_AHB/n116 ;
  wire [31:0] \U_AHB/n117 ;
  wire [31:0] \U_AHB/n118 ;
  wire [31:0] \U_AHB/n37 ;
  wire [31:0] \U_AHB/n39 ;
  wire [31:0] \U_AHB/n40 ;
  wire [31:0] \U_AHB/n41 ;
  wire [31:0] \U_AHB/n42 ;
  wire  \U_AHB/sel0_b0/B0 ;
  wire  \U_AHB/sel0_b0/B1 ;
  wire  \U_AHB/sel0_b0/B10 ;
  wire  \U_AHB/sel0_b0/B11 ;
  wire  \U_AHB/sel0_b0/B2 ;
  wire  \U_AHB/sel0_b0/B3 ;
  wire  \U_AHB/sel0_b0/B4 ;
  wire  \U_AHB/sel0_b0/B5 ;
  wire  \U_AHB/sel0_b0/B6 ;
  wire  \U_AHB/sel0_b0/B7 ;
  wire  \U_AHB/sel0_b0/B8 ;
  wire  \U_AHB/sel0_b0/B9 ;
  wire  \U_AHB/sel0_b1/B0 ;
  wire  \U_AHB/sel0_b1/B1 ;
  wire  \U_AHB/sel0_b1/B10 ;
  wire  \U_AHB/sel0_b1/B11 ;
  wire  \U_AHB/sel0_b1/B2 ;
  wire  \U_AHB/sel0_b1/B3 ;
  wire  \U_AHB/sel0_b1/B4 ;
  wire  \U_AHB/sel0_b1/B5 ;
  wire  \U_AHB/sel0_b1/B6 ;
  wire  \U_AHB/sel0_b1/B7 ;
  wire  \U_AHB/sel0_b1/B8 ;
  wire  \U_AHB/sel0_b1/B9 ;
  wire  \U_AHB/sel0_b10/B0 ;
  wire  \U_AHB/sel0_b10/B1 ;
  wire  \U_AHB/sel0_b10/B10 ;
  wire  \U_AHB/sel0_b10/B11 ;
  wire  \U_AHB/sel0_b10/B2 ;
  wire  \U_AHB/sel0_b10/B3 ;
  wire  \U_AHB/sel0_b10/B4 ;
  wire  \U_AHB/sel0_b10/B5 ;
  wire  \U_AHB/sel0_b10/B6 ;
  wire  \U_AHB/sel0_b10/B7 ;
  wire  \U_AHB/sel0_b10/B8 ;
  wire  \U_AHB/sel0_b10/B9 ;
  wire  \U_AHB/sel0_b11/B0 ;
  wire  \U_AHB/sel0_b11/B1 ;
  wire  \U_AHB/sel0_b11/B10 ;
  wire  \U_AHB/sel0_b11/B11 ;
  wire  \U_AHB/sel0_b11/B2 ;
  wire  \U_AHB/sel0_b11/B3 ;
  wire  \U_AHB/sel0_b11/B4 ;
  wire  \U_AHB/sel0_b11/B5 ;
  wire  \U_AHB/sel0_b11/B6 ;
  wire  \U_AHB/sel0_b11/B7 ;
  wire  \U_AHB/sel0_b11/B8 ;
  wire  \U_AHB/sel0_b11/B9 ;
  wire  \U_AHB/sel0_b12/B0 ;
  wire  \U_AHB/sel0_b12/B1 ;
  wire  \U_AHB/sel0_b12/B10 ;
  wire  \U_AHB/sel0_b12/B11 ;
  wire  \U_AHB/sel0_b12/B2 ;
  wire  \U_AHB/sel0_b12/B3 ;
  wire  \U_AHB/sel0_b12/B4 ;
  wire  \U_AHB/sel0_b12/B5 ;
  wire  \U_AHB/sel0_b12/B6 ;
  wire  \U_AHB/sel0_b12/B7 ;
  wire  \U_AHB/sel0_b12/B8 ;
  wire  \U_AHB/sel0_b12/B9 ;
  wire  \U_AHB/sel0_b13/B0 ;
  wire  \U_AHB/sel0_b13/B1 ;
  wire  \U_AHB/sel0_b13/B10 ;
  wire  \U_AHB/sel0_b13/B11 ;
  wire  \U_AHB/sel0_b13/B2 ;
  wire  \U_AHB/sel0_b13/B3 ;
  wire  \U_AHB/sel0_b13/B4 ;
  wire  \U_AHB/sel0_b13/B5 ;
  wire  \U_AHB/sel0_b13/B6 ;
  wire  \U_AHB/sel0_b13/B7 ;
  wire  \U_AHB/sel0_b13/B8 ;
  wire  \U_AHB/sel0_b13/B9 ;
  wire  \U_AHB/sel0_b14/B0 ;
  wire  \U_AHB/sel0_b14/B1 ;
  wire  \U_AHB/sel0_b14/B10 ;
  wire  \U_AHB/sel0_b14/B11 ;
  wire  \U_AHB/sel0_b14/B2 ;
  wire  \U_AHB/sel0_b14/B3 ;
  wire  \U_AHB/sel0_b14/B4 ;
  wire  \U_AHB/sel0_b14/B5 ;
  wire  \U_AHB/sel0_b14/B6 ;
  wire  \U_AHB/sel0_b14/B7 ;
  wire  \U_AHB/sel0_b14/B8 ;
  wire  \U_AHB/sel0_b14/B9 ;
  wire  \U_AHB/sel0_b15/B0 ;
  wire  \U_AHB/sel0_b15/B1 ;
  wire  \U_AHB/sel0_b15/B10 ;
  wire  \U_AHB/sel0_b15/B11 ;
  wire  \U_AHB/sel0_b15/B2 ;
  wire  \U_AHB/sel0_b15/B3 ;
  wire  \U_AHB/sel0_b15/B4 ;
  wire  \U_AHB/sel0_b15/B5 ;
  wire  \U_AHB/sel0_b15/B6 ;
  wire  \U_AHB/sel0_b15/B7 ;
  wire  \U_AHB/sel0_b15/B8 ;
  wire  \U_AHB/sel0_b15/B9 ;
  wire  \U_AHB/sel0_b16/B0 ;
  wire  \U_AHB/sel0_b16/B1 ;
  wire  \U_AHB/sel0_b16/B10 ;
  wire  \U_AHB/sel0_b16/B11 ;
  wire  \U_AHB/sel0_b16/B2 ;
  wire  \U_AHB/sel0_b16/B3 ;
  wire  \U_AHB/sel0_b16/B4 ;
  wire  \U_AHB/sel0_b16/B5 ;
  wire  \U_AHB/sel0_b16/B6 ;
  wire  \U_AHB/sel0_b16/B7 ;
  wire  \U_AHB/sel0_b16/B8 ;
  wire  \U_AHB/sel0_b16/B9 ;
  wire  \U_AHB/sel0_b17/B0 ;
  wire  \U_AHB/sel0_b17/B1 ;
  wire  \U_AHB/sel0_b17/B10 ;
  wire  \U_AHB/sel0_b17/B11 ;
  wire  \U_AHB/sel0_b17/B2 ;
  wire  \U_AHB/sel0_b17/B3 ;
  wire  \U_AHB/sel0_b17/B4 ;
  wire  \U_AHB/sel0_b17/B5 ;
  wire  \U_AHB/sel0_b17/B6 ;
  wire  \U_AHB/sel0_b17/B7 ;
  wire  \U_AHB/sel0_b17/B8 ;
  wire  \U_AHB/sel0_b17/B9 ;
  wire  \U_AHB/sel0_b18/B0 ;
  wire  \U_AHB/sel0_b18/B1 ;
  wire  \U_AHB/sel0_b18/B10 ;
  wire  \U_AHB/sel0_b18/B11 ;
  wire  \U_AHB/sel0_b18/B2 ;
  wire  \U_AHB/sel0_b18/B3 ;
  wire  \U_AHB/sel0_b18/B4 ;
  wire  \U_AHB/sel0_b18/B5 ;
  wire  \U_AHB/sel0_b18/B6 ;
  wire  \U_AHB/sel0_b18/B7 ;
  wire  \U_AHB/sel0_b18/B8 ;
  wire  \U_AHB/sel0_b18/B9 ;
  wire  \U_AHB/sel0_b19/B0 ;
  wire  \U_AHB/sel0_b19/B1 ;
  wire  \U_AHB/sel0_b19/B10 ;
  wire  \U_AHB/sel0_b19/B11 ;
  wire  \U_AHB/sel0_b19/B2 ;
  wire  \U_AHB/sel0_b19/B3 ;
  wire  \U_AHB/sel0_b19/B4 ;
  wire  \U_AHB/sel0_b19/B5 ;
  wire  \U_AHB/sel0_b19/B6 ;
  wire  \U_AHB/sel0_b19/B7 ;
  wire  \U_AHB/sel0_b19/B8 ;
  wire  \U_AHB/sel0_b19/B9 ;
  wire  \U_AHB/sel0_b2/B0 ;
  wire  \U_AHB/sel0_b2/B1 ;
  wire  \U_AHB/sel0_b2/B10 ;
  wire  \U_AHB/sel0_b2/B11 ;
  wire  \U_AHB/sel0_b2/B2 ;
  wire  \U_AHB/sel0_b2/B3 ;
  wire  \U_AHB/sel0_b2/B4 ;
  wire  \U_AHB/sel0_b2/B5 ;
  wire  \U_AHB/sel0_b2/B6 ;
  wire  \U_AHB/sel0_b2/B7 ;
  wire  \U_AHB/sel0_b2/B8 ;
  wire  \U_AHB/sel0_b2/B9 ;
  wire  \U_AHB/sel0_b20/B0 ;
  wire  \U_AHB/sel0_b20/B1 ;
  wire  \U_AHB/sel0_b20/B10 ;
  wire  \U_AHB/sel0_b20/B11 ;
  wire  \U_AHB/sel0_b20/B2 ;
  wire  \U_AHB/sel0_b20/B3 ;
  wire  \U_AHB/sel0_b20/B4 ;
  wire  \U_AHB/sel0_b20/B5 ;
  wire  \U_AHB/sel0_b20/B6 ;
  wire  \U_AHB/sel0_b20/B7 ;
  wire  \U_AHB/sel0_b20/B8 ;
  wire  \U_AHB/sel0_b20/B9 ;
  wire  \U_AHB/sel0_b21/B0 ;
  wire  \U_AHB/sel0_b21/B1 ;
  wire  \U_AHB/sel0_b21/B10 ;
  wire  \U_AHB/sel0_b21/B11 ;
  wire  \U_AHB/sel0_b21/B2 ;
  wire  \U_AHB/sel0_b21/B3 ;
  wire  \U_AHB/sel0_b21/B4 ;
  wire  \U_AHB/sel0_b21/B5 ;
  wire  \U_AHB/sel0_b21/B6 ;
  wire  \U_AHB/sel0_b21/B7 ;
  wire  \U_AHB/sel0_b21/B8 ;
  wire  \U_AHB/sel0_b21/B9 ;
  wire  \U_AHB/sel0_b22/B0 ;
  wire  \U_AHB/sel0_b22/B1 ;
  wire  \U_AHB/sel0_b22/B10 ;
  wire  \U_AHB/sel0_b22/B11 ;
  wire  \U_AHB/sel0_b22/B2 ;
  wire  \U_AHB/sel0_b22/B3 ;
  wire  \U_AHB/sel0_b22/B4 ;
  wire  \U_AHB/sel0_b22/B5 ;
  wire  \U_AHB/sel0_b22/B6 ;
  wire  \U_AHB/sel0_b22/B7 ;
  wire  \U_AHB/sel0_b22/B8 ;
  wire  \U_AHB/sel0_b22/B9 ;
  wire  \U_AHB/sel0_b23/B0 ;
  wire  \U_AHB/sel0_b23/B1 ;
  wire  \U_AHB/sel0_b23/B10 ;
  wire  \U_AHB/sel0_b23/B11 ;
  wire  \U_AHB/sel0_b23/B2 ;
  wire  \U_AHB/sel0_b23/B3 ;
  wire  \U_AHB/sel0_b23/B4 ;
  wire  \U_AHB/sel0_b23/B5 ;
  wire  \U_AHB/sel0_b23/B6 ;
  wire  \U_AHB/sel0_b23/B7 ;
  wire  \U_AHB/sel0_b23/B8 ;
  wire  \U_AHB/sel0_b23/B9 ;
  wire  \U_AHB/sel0_b3/B0 ;
  wire  \U_AHB/sel0_b3/B1 ;
  wire  \U_AHB/sel0_b3/B10 ;
  wire  \U_AHB/sel0_b3/B11 ;
  wire  \U_AHB/sel0_b3/B2 ;
  wire  \U_AHB/sel0_b3/B3 ;
  wire  \U_AHB/sel0_b3/B4 ;
  wire  \U_AHB/sel0_b3/B5 ;
  wire  \U_AHB/sel0_b3/B6 ;
  wire  \U_AHB/sel0_b3/B7 ;
  wire  \U_AHB/sel0_b3/B8 ;
  wire  \U_AHB/sel0_b3/B9 ;
  wire  \U_AHB/sel0_b4/B0 ;
  wire  \U_AHB/sel0_b4/B1 ;
  wire  \U_AHB/sel0_b4/B10 ;
  wire  \U_AHB/sel0_b4/B11 ;
  wire  \U_AHB/sel0_b4/B2 ;
  wire  \U_AHB/sel0_b4/B3 ;
  wire  \U_AHB/sel0_b4/B4 ;
  wire  \U_AHB/sel0_b4/B5 ;
  wire  \U_AHB/sel0_b4/B6 ;
  wire  \U_AHB/sel0_b4/B7 ;
  wire  \U_AHB/sel0_b4/B8 ;
  wire  \U_AHB/sel0_b4/B9 ;
  wire  \U_AHB/sel0_b5/B0 ;
  wire  \U_AHB/sel0_b5/B1 ;
  wire  \U_AHB/sel0_b5/B10 ;
  wire  \U_AHB/sel0_b5/B11 ;
  wire  \U_AHB/sel0_b5/B2 ;
  wire  \U_AHB/sel0_b5/B3 ;
  wire  \U_AHB/sel0_b5/B4 ;
  wire  \U_AHB/sel0_b5/B5 ;
  wire  \U_AHB/sel0_b5/B6 ;
  wire  \U_AHB/sel0_b5/B7 ;
  wire  \U_AHB/sel0_b5/B8 ;
  wire  \U_AHB/sel0_b5/B9 ;
  wire  \U_AHB/sel0_b6/B0 ;
  wire  \U_AHB/sel0_b6/B1 ;
  wire  \U_AHB/sel0_b6/B10 ;
  wire  \U_AHB/sel0_b6/B11 ;
  wire  \U_AHB/sel0_b6/B2 ;
  wire  \U_AHB/sel0_b6/B3 ;
  wire  \U_AHB/sel0_b6/B4 ;
  wire  \U_AHB/sel0_b6/B5 ;
  wire  \U_AHB/sel0_b6/B6 ;
  wire  \U_AHB/sel0_b6/B7 ;
  wire  \U_AHB/sel0_b6/B8 ;
  wire  \U_AHB/sel0_b6/B9 ;
  wire  \U_AHB/sel0_b7/B0 ;
  wire  \U_AHB/sel0_b7/B1 ;
  wire  \U_AHB/sel0_b7/B10 ;
  wire  \U_AHB/sel0_b7/B11 ;
  wire  \U_AHB/sel0_b7/B2 ;
  wire  \U_AHB/sel0_b7/B3 ;
  wire  \U_AHB/sel0_b7/B4 ;
  wire  \U_AHB/sel0_b7/B5 ;
  wire  \U_AHB/sel0_b7/B6 ;
  wire  \U_AHB/sel0_b7/B7 ;
  wire  \U_AHB/sel0_b7/B8 ;
  wire  \U_AHB/sel0_b7/B9 ;
  wire  \U_AHB/sel0_b8/B0 ;
  wire  \U_AHB/sel0_b8/B1 ;
  wire  \U_AHB/sel0_b8/B10 ;
  wire  \U_AHB/sel0_b8/B11 ;
  wire  \U_AHB/sel0_b8/B2 ;
  wire  \U_AHB/sel0_b8/B3 ;
  wire  \U_AHB/sel0_b8/B4 ;
  wire  \U_AHB/sel0_b8/B5 ;
  wire  \U_AHB/sel0_b8/B6 ;
  wire  \U_AHB/sel0_b8/B7 ;
  wire  \U_AHB/sel0_b8/B8 ;
  wire  \U_AHB/sel0_b8/B9 ;
  wire  \U_AHB/sel0_b9/B0 ;
  wire  \U_AHB/sel0_b9/B1 ;
  wire  \U_AHB/sel0_b9/B10 ;
  wire  \U_AHB/sel0_b9/B11 ;
  wire  \U_AHB/sel0_b9/B2 ;
  wire  \U_AHB/sel0_b9/B3 ;
  wire  \U_AHB/sel0_b9/B4 ;
  wire  \U_AHB/sel0_b9/B5 ;
  wire  \U_AHB/sel0_b9/B6 ;
  wire  \U_AHB/sel0_b9/B7 ;
  wire  \U_AHB/sel0_b9/B8 ;
  wire  \U_AHB/sel0_b9/B9 ;
  wire  \U_AHB/sel1_b0/B0 ;
  wire  \U_AHB/sel1_b0/B1 ;
  wire  \U_AHB/sel1_b0/B3 ;
  wire  \U_AHB/sel1_b0/B4 ;
  wire  \U_AHB/sel1_b0/B5 ;
  wire  \U_AHB/sel1_b0/B6 ;
  wire  \U_AHB/sel1_b0/B7 ;
  wire  \U_AHB/sel1_b0/B8 ;
  wire  \U_AHB/sel1_b1/B0 ;
  wire  \U_AHB/sel1_b1/B1 ;
  wire  \U_AHB/sel1_b1/B3 ;
  wire  \U_AHB/sel1_b1/B4 ;
  wire  \U_AHB/sel1_b1/B5 ;
  wire  \U_AHB/sel1_b1/B6 ;
  wire  \U_AHB/sel1_b1/B7 ;
  wire  \U_AHB/sel1_b1/B8 ;
  wire  \U_AHB/sel1_b10/B0 ;
  wire  \U_AHB/sel1_b10/B1 ;
  wire  \U_AHB/sel1_b10/B3 ;
  wire  \U_AHB/sel1_b10/B4 ;
  wire  \U_AHB/sel1_b10/B5 ;
  wire  \U_AHB/sel1_b10/B6 ;
  wire  \U_AHB/sel1_b10/B7 ;
  wire  \U_AHB/sel1_b10/B8 ;
  wire  \U_AHB/sel1_b11/B0 ;
  wire  \U_AHB/sel1_b11/B1 ;
  wire  \U_AHB/sel1_b11/B3 ;
  wire  \U_AHB/sel1_b11/B4 ;
  wire  \U_AHB/sel1_b11/B5 ;
  wire  \U_AHB/sel1_b11/B6 ;
  wire  \U_AHB/sel1_b11/B7 ;
  wire  \U_AHB/sel1_b11/B8 ;
  wire  \U_AHB/sel1_b12/B0 ;
  wire  \U_AHB/sel1_b12/B1 ;
  wire  \U_AHB/sel1_b12/B3 ;
  wire  \U_AHB/sel1_b12/B4 ;
  wire  \U_AHB/sel1_b12/B5 ;
  wire  \U_AHB/sel1_b12/B6 ;
  wire  \U_AHB/sel1_b12/B7 ;
  wire  \U_AHB/sel1_b12/B8 ;
  wire  \U_AHB/sel1_b13/B0 ;
  wire  \U_AHB/sel1_b13/B1 ;
  wire  \U_AHB/sel1_b13/B3 ;
  wire  \U_AHB/sel1_b13/B4 ;
  wire  \U_AHB/sel1_b13/B5 ;
  wire  \U_AHB/sel1_b13/B6 ;
  wire  \U_AHB/sel1_b13/B7 ;
  wire  \U_AHB/sel1_b13/B8 ;
  wire  \U_AHB/sel1_b14/B0 ;
  wire  \U_AHB/sel1_b14/B1 ;
  wire  \U_AHB/sel1_b14/B3 ;
  wire  \U_AHB/sel1_b14/B4 ;
  wire  \U_AHB/sel1_b14/B5 ;
  wire  \U_AHB/sel1_b14/B6 ;
  wire  \U_AHB/sel1_b14/B7 ;
  wire  \U_AHB/sel1_b14/B8 ;
  wire  \U_AHB/sel1_b15/B0 ;
  wire  \U_AHB/sel1_b15/B1 ;
  wire  \U_AHB/sel1_b15/B3 ;
  wire  \U_AHB/sel1_b15/B4 ;
  wire  \U_AHB/sel1_b15/B5 ;
  wire  \U_AHB/sel1_b15/B6 ;
  wire  \U_AHB/sel1_b15/B7 ;
  wire  \U_AHB/sel1_b15/B8 ;
  wire  \U_AHB/sel1_b16/B0 ;
  wire  \U_AHB/sel1_b16/B1 ;
  wire  \U_AHB/sel1_b16/B4 ;
  wire  \U_AHB/sel1_b16/B5 ;
  wire  \U_AHB/sel1_b16/B6 ;
  wire  \U_AHB/sel1_b16/B7 ;
  wire  \U_AHB/sel1_b16/B8 ;
  wire  \U_AHB/sel1_b17/B0 ;
  wire  \U_AHB/sel1_b17/B1 ;
  wire  \U_AHB/sel1_b17/B4 ;
  wire  \U_AHB/sel1_b17/B5 ;
  wire  \U_AHB/sel1_b17/B6 ;
  wire  \U_AHB/sel1_b17/B7 ;
  wire  \U_AHB/sel1_b17/B8 ;
  wire  \U_AHB/sel1_b18/B0 ;
  wire  \U_AHB/sel1_b18/B1 ;
  wire  \U_AHB/sel1_b18/B3 ;
  wire  \U_AHB/sel1_b18/B4 ;
  wire  \U_AHB/sel1_b18/B5 ;
  wire  \U_AHB/sel1_b18/B6 ;
  wire  \U_AHB/sel1_b18/B7 ;
  wire  \U_AHB/sel1_b18/B8 ;
  wire  \U_AHB/sel1_b19/B0 ;
  wire  \U_AHB/sel1_b19/B1 ;
  wire  \U_AHB/sel1_b19/B3 ;
  wire  \U_AHB/sel1_b19/B4 ;
  wire  \U_AHB/sel1_b19/B5 ;
  wire  \U_AHB/sel1_b19/B6 ;
  wire  \U_AHB/sel1_b19/B7 ;
  wire  \U_AHB/sel1_b19/B8 ;
  wire  \U_AHB/sel1_b2/B0 ;
  wire  \U_AHB/sel1_b2/B1 ;
  wire  \U_AHB/sel1_b2/B4 ;
  wire  \U_AHB/sel1_b2/B5 ;
  wire  \U_AHB/sel1_b2/B6 ;
  wire  \U_AHB/sel1_b2/B7 ;
  wire  \U_AHB/sel1_b2/B8 ;
  wire  \U_AHB/sel1_b20/B0 ;
  wire  \U_AHB/sel1_b20/B1 ;
  wire  \U_AHB/sel1_b20/B3 ;
  wire  \U_AHB/sel1_b20/B4 ;
  wire  \U_AHB/sel1_b20/B5 ;
  wire  \U_AHB/sel1_b20/B6 ;
  wire  \U_AHB/sel1_b20/B7 ;
  wire  \U_AHB/sel1_b20/B8 ;
  wire  \U_AHB/sel1_b21/B0 ;
  wire  \U_AHB/sel1_b21/B1 ;
  wire  \U_AHB/sel1_b21/B3 ;
  wire  \U_AHB/sel1_b21/B4 ;
  wire  \U_AHB/sel1_b21/B5 ;
  wire  \U_AHB/sel1_b21/B6 ;
  wire  \U_AHB/sel1_b21/B7 ;
  wire  \U_AHB/sel1_b21/B8 ;
  wire  \U_AHB/sel1_b22/B0 ;
  wire  \U_AHB/sel1_b22/B1 ;
  wire  \U_AHB/sel1_b22/B3 ;
  wire  \U_AHB/sel1_b22/B4 ;
  wire  \U_AHB/sel1_b22/B5 ;
  wire  \U_AHB/sel1_b22/B6 ;
  wire  \U_AHB/sel1_b22/B7 ;
  wire  \U_AHB/sel1_b22/B8 ;
  wire  \U_AHB/sel1_b23/B0 ;
  wire  \U_AHB/sel1_b23/B1 ;
  wire  \U_AHB/sel1_b23/B3 ;
  wire  \U_AHB/sel1_b23/B4 ;
  wire  \U_AHB/sel1_b23/B5 ;
  wire  \U_AHB/sel1_b23/B6 ;
  wire  \U_AHB/sel1_b23/B7 ;
  wire  \U_AHB/sel1_b23/B8 ;
  wire  \U_AHB/sel1_b24/B0 ;
  wire  \U_AHB/sel1_b24/B1 ;
  wire  \U_AHB/sel1_b24/B3 ;
  wire  \U_AHB/sel1_b25/B0 ;
  wire  \U_AHB/sel1_b25/B1 ;
  wire  \U_AHB/sel1_b25/B3 ;
  wire  \U_AHB/sel1_b26/B0 ;
  wire  \U_AHB/sel1_b26/B1 ;
  wire  \U_AHB/sel1_b27/B0 ;
  wire  \U_AHB/sel1_b27/B1 ;
  wire  \U_AHB/sel1_b28/B0 ;
  wire  \U_AHB/sel1_b28/B1 ;
  wire  \U_AHB/sel1_b29/B0 ;
  wire  \U_AHB/sel1_b29/B1 ;
  wire  \U_AHB/sel1_b3/B0 ;
  wire  \U_AHB/sel1_b3/B1 ;
  wire  \U_AHB/sel1_b3/B4 ;
  wire  \U_AHB/sel1_b3/B5 ;
  wire  \U_AHB/sel1_b3/B6 ;
  wire  \U_AHB/sel1_b3/B7 ;
  wire  \U_AHB/sel1_b3/B8 ;
  wire  \U_AHB/sel1_b30/B0 ;
  wire  \U_AHB/sel1_b30/B1 ;
  wire  \U_AHB/sel1_b31/B0 ;
  wire  \U_AHB/sel1_b31/B1 ;
  wire  \U_AHB/sel1_b4/B0 ;
  wire  \U_AHB/sel1_b4/B1 ;
  wire  \U_AHB/sel1_b4/B4 ;
  wire  \U_AHB/sel1_b4/B5 ;
  wire  \U_AHB/sel1_b4/B6 ;
  wire  \U_AHB/sel1_b4/B7 ;
  wire  \U_AHB/sel1_b4/B8 ;
  wire  \U_AHB/sel1_b5/B0 ;
  wire  \U_AHB/sel1_b5/B1 ;
  wire  \U_AHB/sel1_b5/B4 ;
  wire  \U_AHB/sel1_b5/B5 ;
  wire  \U_AHB/sel1_b5/B6 ;
  wire  \U_AHB/sel1_b5/B7 ;
  wire  \U_AHB/sel1_b5/B8 ;
  wire  \U_AHB/sel1_b6/B0 ;
  wire  \U_AHB/sel1_b6/B1 ;
  wire  \U_AHB/sel1_b6/B4 ;
  wire  \U_AHB/sel1_b6/B5 ;
  wire  \U_AHB/sel1_b6/B6 ;
  wire  \U_AHB/sel1_b6/B7 ;
  wire  \U_AHB/sel1_b6/B8 ;
  wire  \U_AHB/sel1_b7/B0 ;
  wire  \U_AHB/sel1_b7/B1 ;
  wire  \U_AHB/sel1_b7/B4 ;
  wire  \U_AHB/sel1_b7/B5 ;
  wire  \U_AHB/sel1_b7/B6 ;
  wire  \U_AHB/sel1_b7/B7 ;
  wire  \U_AHB/sel1_b7/B8 ;
  wire  \U_AHB/sel1_b8/B0 ;
  wire  \U_AHB/sel1_b8/B1 ;
  wire  \U_AHB/sel1_b8/B4 ;
  wire  \U_AHB/sel1_b8/B5 ;
  wire  \U_AHB/sel1_b8/B6 ;
  wire  \U_AHB/sel1_b8/B7 ;
  wire  \U_AHB/sel1_b8/B8 ;
  wire  \U_AHB/sel1_b9/B0 ;
  wire  \U_AHB/sel1_b9/B1 ;
  wire  \U_AHB/sel1_b9/B4 ;
  wire  \U_AHB/sel1_b9/B5 ;
  wire  \U_AHB/sel1_b9/B6 ;
  wire  \U_AHB/sel1_b9/B7 ;
  wire  \U_AHB/sel1_b9/B8 ;
  wire [31:0] freq0;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freq1;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freq2;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freq3;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freq4;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freq5;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freq6;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freq7;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freq8;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freq9;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freqA;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freqB;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freqC;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freqD;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freqE;  // CPLD_SOC_AHB_TOP.v(55)
  wire [31:0] freqF;  // CPLD_SOC_AHB_TOP.v(55)
  wire [3:0] n10;
  wire [31:0] n2;
  wire [31:0] n3;
  wire [3:0] n7;
  wire [3:0] n8;
  wire [3:0] n9;
  wire [32:0] pnum0;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnum1;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnum2;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnum3;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnum4;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnum5;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnum6;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnum7;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnum8;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnum9;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnumA;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnumB;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnumC;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnumD;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnumE;  // CPLD_SOC_AHB_TOP.v(54)
  wire [32:0] pnumF;  // CPLD_SOC_AHB_TOP.v(54)
  wire [23:0] pnumcnt0;  // CPLD_SOC_AHB_TOP.v(61)
  wire [23:0] pnumcnt1;  // CPLD_SOC_AHB_TOP.v(62)
  wire [23:0] pnumcnt2;  // CPLD_SOC_AHB_TOP.v(63)
  wire [23:0] pnumcnt3;  // CPLD_SOC_AHB_TOP.v(64)
  wire [23:0] pnumcnt4;  // CPLD_SOC_AHB_TOP.v(65)
  wire [23:0] pnumcnt5;  // CPLD_SOC_AHB_TOP.v(66)
  wire [23:0] pnumcnt6;  // CPLD_SOC_AHB_TOP.v(67)
  wire [23:0] pnumcnt7;  // CPLD_SOC_AHB_TOP.v(68)
  wire [23:0] pnumcnt8;  // CPLD_SOC_AHB_TOP.v(69)
  wire [23:0] pnumcnt9;  // CPLD_SOC_AHB_TOP.v(70)
  wire [23:0] pnumcntA;  // CPLD_SOC_AHB_TOP.v(71)
  wire [23:0] pnumcntB;  // CPLD_SOC_AHB_TOP.v(72)
  wire [23:0] pnumcntC;  // CPLD_SOC_AHB_TOP.v(73)
  wire [23:0] pnumcntD;  // CPLD_SOC_AHB_TOP.v(74)
  wire [23:0] pnumcntE;  // CPLD_SOC_AHB_TOP.v(75)
  wire [23:0] pnumcntF;  // CPLD_SOC_AHB_TOP.v(76)
  wire [31:0] pwm_start_stop;  // CPLD_SOC_AHB_TOP.v(52)
  wire [15:0] pwm_state_read;  // CPLD_SOC_AHB_TOP.v(78)
  wire [31:0] timer;  // CPLD_SOC_AHB_TOP.v(26)
  wire \PWM0/RemaTxNum[0]_keep ;
  wire \PWM0/RemaTxNum[10]_keep ;
  wire \PWM0/RemaTxNum[11]_keep ;
  wire \PWM0/RemaTxNum[12]_keep ;
  wire \PWM0/RemaTxNum[13]_keep ;
  wire \PWM0/RemaTxNum[14]_keep ;
  wire \PWM0/RemaTxNum[15]_keep ;
  wire \PWM0/RemaTxNum[16]_keep ;
  wire \PWM0/RemaTxNum[17]_keep ;
  wire \PWM0/RemaTxNum[18]_keep ;
  wire \PWM0/RemaTxNum[19]_keep ;
  wire \PWM0/RemaTxNum[1]_keep ;
  wire \PWM0/RemaTxNum[20]_keep ;
  wire \PWM0/RemaTxNum[21]_keep ;
  wire \PWM0/RemaTxNum[22]_keep ;
  wire \PWM0/RemaTxNum[23]_keep ;
  wire \PWM0/RemaTxNum[2]_keep ;
  wire \PWM0/RemaTxNum[3]_keep ;
  wire \PWM0/RemaTxNum[4]_keep ;
  wire \PWM0/RemaTxNum[5]_keep ;
  wire \PWM0/RemaTxNum[6]_keep ;
  wire \PWM0/RemaTxNum[7]_keep ;
  wire \PWM0/RemaTxNum[8]_keep ;
  wire \PWM0/RemaTxNum[9]_keep ;
  wire \PWM0/dir_keep ;
  wire \PWM0/mux3_b0_sel_is_3_o ;
  wire \PWM0/n0 ;
  wire \PWM0/n1 ;
  wire \PWM0/n10 ;
  wire \PWM0/n11 ;
  wire \PWM0/n17 ;
  wire \PWM0/n17_neg ;
  wire \PWM0/n18 ;
  wire \PWM0/n24 ;
  wire \PWM0/n25 ;
  wire \PWM0/n25_neg ;
  wire \PWM0/n32 ;
  wire \PWM0/n4 ;
  wire \PWM0/n4_neg ;
  wire \PWM0/n5 ;
  wire \PWM0/n6 ;
  wire \PWM0/n6_neg ;
  wire \PWM0/n8 ;
  wire \PWM0/n9 ;
  wire \PWM0/pnumr[0]_keep ;
  wire \PWM0/pnumr[10]_keep ;
  wire \PWM0/pnumr[11]_keep ;
  wire \PWM0/pnumr[12]_keep ;
  wire \PWM0/pnumr[13]_keep ;
  wire \PWM0/pnumr[14]_keep ;
  wire \PWM0/pnumr[15]_keep ;
  wire \PWM0/pnumr[16]_keep ;
  wire \PWM0/pnumr[17]_keep ;
  wire \PWM0/pnumr[18]_keep ;
  wire \PWM0/pnumr[19]_keep ;
  wire \PWM0/pnumr[1]_keep ;
  wire \PWM0/pnumr[20]_keep ;
  wire \PWM0/pnumr[21]_keep ;
  wire \PWM0/pnumr[22]_keep ;
  wire \PWM0/pnumr[23]_keep ;
  wire \PWM0/pnumr[24]_keep ;
  wire \PWM0/pnumr[25]_keep ;
  wire \PWM0/pnumr[26]_keep ;
  wire \PWM0/pnumr[27]_keep ;
  wire \PWM0/pnumr[28]_keep ;
  wire \PWM0/pnumr[29]_keep ;
  wire \PWM0/pnumr[2]_keep ;
  wire \PWM0/pnumr[30]_keep ;
  wire \PWM0/pnumr[31]_keep ;
  wire \PWM0/pnumr[3]_keep ;
  wire \PWM0/pnumr[4]_keep ;
  wire \PWM0/pnumr[5]_keep ;
  wire \PWM0/pnumr[6]_keep ;
  wire \PWM0/pnumr[7]_keep ;
  wire \PWM0/pnumr[8]_keep ;
  wire \PWM0/pnumr[9]_keep ;
  wire \PWM0/pwm_keep ;
  wire \PWM0/stopreq ;  // src/OnePWM.v(14)
  wire \PWM0/stopreq_keep ;
  wire \PWM0/u14_sel_is_1_o ;
  wire \PWM0/u17_sel_is_1_o ;
  wire \PWM0/u17_sel_is_1_o_neg ;
  wire \PWM0/u18_sel_is_0_o ;
  wire \PWM0/u8_sel_is_0_o ;
  wire \PWM1/RemaTxNum[0]_keep ;
  wire \PWM1/RemaTxNum[10]_keep ;
  wire \PWM1/RemaTxNum[11]_keep ;
  wire \PWM1/RemaTxNum[12]_keep ;
  wire \PWM1/RemaTxNum[13]_keep ;
  wire \PWM1/RemaTxNum[14]_keep ;
  wire \PWM1/RemaTxNum[15]_keep ;
  wire \PWM1/RemaTxNum[16]_keep ;
  wire \PWM1/RemaTxNum[17]_keep ;
  wire \PWM1/RemaTxNum[18]_keep ;
  wire \PWM1/RemaTxNum[19]_keep ;
  wire \PWM1/RemaTxNum[1]_keep ;
  wire \PWM1/RemaTxNum[20]_keep ;
  wire \PWM1/RemaTxNum[21]_keep ;
  wire \PWM1/RemaTxNum[22]_keep ;
  wire \PWM1/RemaTxNum[23]_keep ;
  wire \PWM1/RemaTxNum[2]_keep ;
  wire \PWM1/RemaTxNum[3]_keep ;
  wire \PWM1/RemaTxNum[4]_keep ;
  wire \PWM1/RemaTxNum[5]_keep ;
  wire \PWM1/RemaTxNum[6]_keep ;
  wire \PWM1/RemaTxNum[7]_keep ;
  wire \PWM1/RemaTxNum[8]_keep ;
  wire \PWM1/RemaTxNum[9]_keep ;
  wire \PWM1/dir_keep ;
  wire \PWM1/mux3_b0_sel_is_3_o ;
  wire \PWM1/n0 ;
  wire \PWM1/n1 ;
  wire \PWM1/n10 ;
  wire \PWM1/n11 ;
  wire \PWM1/n17 ;
  wire \PWM1/n17_neg ;
  wire \PWM1/n18 ;
  wire \PWM1/n24 ;
  wire \PWM1/n25 ;
  wire \PWM1/n25_neg ;
  wire \PWM1/n32 ;
  wire \PWM1/n4 ;
  wire \PWM1/n4_neg ;
  wire \PWM1/n5 ;
  wire \PWM1/n6 ;
  wire \PWM1/n6_neg ;
  wire \PWM1/n8 ;
  wire \PWM1/n9 ;
  wire \PWM1/pnumr[0]_keep ;
  wire \PWM1/pnumr[10]_keep ;
  wire \PWM1/pnumr[11]_keep ;
  wire \PWM1/pnumr[12]_keep ;
  wire \PWM1/pnumr[13]_keep ;
  wire \PWM1/pnumr[14]_keep ;
  wire \PWM1/pnumr[15]_keep ;
  wire \PWM1/pnumr[16]_keep ;
  wire \PWM1/pnumr[17]_keep ;
  wire \PWM1/pnumr[18]_keep ;
  wire \PWM1/pnumr[19]_keep ;
  wire \PWM1/pnumr[1]_keep ;
  wire \PWM1/pnumr[20]_keep ;
  wire \PWM1/pnumr[21]_keep ;
  wire \PWM1/pnumr[22]_keep ;
  wire \PWM1/pnumr[23]_keep ;
  wire \PWM1/pnumr[24]_keep ;
  wire \PWM1/pnumr[25]_keep ;
  wire \PWM1/pnumr[26]_keep ;
  wire \PWM1/pnumr[27]_keep ;
  wire \PWM1/pnumr[28]_keep ;
  wire \PWM1/pnumr[29]_keep ;
  wire \PWM1/pnumr[2]_keep ;
  wire \PWM1/pnumr[30]_keep ;
  wire \PWM1/pnumr[31]_keep ;
  wire \PWM1/pnumr[3]_keep ;
  wire \PWM1/pnumr[4]_keep ;
  wire \PWM1/pnumr[5]_keep ;
  wire \PWM1/pnumr[6]_keep ;
  wire \PWM1/pnumr[7]_keep ;
  wire \PWM1/pnumr[8]_keep ;
  wire \PWM1/pnumr[9]_keep ;
  wire \PWM1/pwm_keep ;
  wire \PWM1/stopreq ;  // src/OnePWM.v(14)
  wire \PWM1/stopreq_keep ;
  wire \PWM1/u14_sel_is_1_o ;
  wire \PWM1/u17_sel_is_1_o ;
  wire \PWM1/u17_sel_is_1_o_neg ;
  wire \PWM1/u18_sel_is_0_o ;
  wire \PWM1/u8_sel_is_0_o ;
  wire \PWM2/RemaTxNum[0]_keep ;
  wire \PWM2/RemaTxNum[10]_keep ;
  wire \PWM2/RemaTxNum[11]_keep ;
  wire \PWM2/RemaTxNum[12]_keep ;
  wire \PWM2/RemaTxNum[13]_keep ;
  wire \PWM2/RemaTxNum[14]_keep ;
  wire \PWM2/RemaTxNum[15]_keep ;
  wire \PWM2/RemaTxNum[16]_keep ;
  wire \PWM2/RemaTxNum[17]_keep ;
  wire \PWM2/RemaTxNum[18]_keep ;
  wire \PWM2/RemaTxNum[19]_keep ;
  wire \PWM2/RemaTxNum[1]_keep ;
  wire \PWM2/RemaTxNum[20]_keep ;
  wire \PWM2/RemaTxNum[21]_keep ;
  wire \PWM2/RemaTxNum[22]_keep ;
  wire \PWM2/RemaTxNum[23]_keep ;
  wire \PWM2/RemaTxNum[2]_keep ;
  wire \PWM2/RemaTxNum[3]_keep ;
  wire \PWM2/RemaTxNum[4]_keep ;
  wire \PWM2/RemaTxNum[5]_keep ;
  wire \PWM2/RemaTxNum[6]_keep ;
  wire \PWM2/RemaTxNum[7]_keep ;
  wire \PWM2/RemaTxNum[8]_keep ;
  wire \PWM2/RemaTxNum[9]_keep ;
  wire \PWM2/dir_keep ;
  wire \PWM2/mux3_b0_sel_is_3_o ;
  wire \PWM2/n0 ;
  wire \PWM2/n1 ;
  wire \PWM2/n10 ;
  wire \PWM2/n11 ;
  wire \PWM2/n17 ;
  wire \PWM2/n17_neg ;
  wire \PWM2/n18 ;
  wire \PWM2/n24 ;
  wire \PWM2/n25 ;
  wire \PWM2/n25_neg ;
  wire \PWM2/n32 ;
  wire \PWM2/n4 ;
  wire \PWM2/n4_neg ;
  wire \PWM2/n5 ;
  wire \PWM2/n6 ;
  wire \PWM2/n6_neg ;
  wire \PWM2/n8 ;
  wire \PWM2/n9 ;
  wire \PWM2/pnumr[0]_keep ;
  wire \PWM2/pnumr[10]_keep ;
  wire \PWM2/pnumr[11]_keep ;
  wire \PWM2/pnumr[12]_keep ;
  wire \PWM2/pnumr[13]_keep ;
  wire \PWM2/pnumr[14]_keep ;
  wire \PWM2/pnumr[15]_keep ;
  wire \PWM2/pnumr[16]_keep ;
  wire \PWM2/pnumr[17]_keep ;
  wire \PWM2/pnumr[18]_keep ;
  wire \PWM2/pnumr[19]_keep ;
  wire \PWM2/pnumr[1]_keep ;
  wire \PWM2/pnumr[20]_keep ;
  wire \PWM2/pnumr[21]_keep ;
  wire \PWM2/pnumr[22]_keep ;
  wire \PWM2/pnumr[23]_keep ;
  wire \PWM2/pnumr[24]_keep ;
  wire \PWM2/pnumr[25]_keep ;
  wire \PWM2/pnumr[26]_keep ;
  wire \PWM2/pnumr[27]_keep ;
  wire \PWM2/pnumr[28]_keep ;
  wire \PWM2/pnumr[29]_keep ;
  wire \PWM2/pnumr[2]_keep ;
  wire \PWM2/pnumr[30]_keep ;
  wire \PWM2/pnumr[31]_keep ;
  wire \PWM2/pnumr[3]_keep ;
  wire \PWM2/pnumr[4]_keep ;
  wire \PWM2/pnumr[5]_keep ;
  wire \PWM2/pnumr[6]_keep ;
  wire \PWM2/pnumr[7]_keep ;
  wire \PWM2/pnumr[8]_keep ;
  wire \PWM2/pnumr[9]_keep ;
  wire \PWM2/pwm_keep ;
  wire \PWM2/stopreq ;  // src/OnePWM.v(14)
  wire \PWM2/stopreq_keep ;
  wire \PWM2/u14_sel_is_1_o ;
  wire \PWM2/u17_sel_is_1_o ;
  wire \PWM2/u17_sel_is_1_o_neg ;
  wire \PWM2/u18_sel_is_0_o ;
  wire \PWM2/u8_sel_is_0_o ;
  wire \PWM3/RemaTxNum[0]_keep ;
  wire \PWM3/RemaTxNum[10]_keep ;
  wire \PWM3/RemaTxNum[11]_keep ;
  wire \PWM3/RemaTxNum[12]_keep ;
  wire \PWM3/RemaTxNum[13]_keep ;
  wire \PWM3/RemaTxNum[14]_keep ;
  wire \PWM3/RemaTxNum[15]_keep ;
  wire \PWM3/RemaTxNum[16]_keep ;
  wire \PWM3/RemaTxNum[17]_keep ;
  wire \PWM3/RemaTxNum[18]_keep ;
  wire \PWM3/RemaTxNum[19]_keep ;
  wire \PWM3/RemaTxNum[1]_keep ;
  wire \PWM3/RemaTxNum[20]_keep ;
  wire \PWM3/RemaTxNum[21]_keep ;
  wire \PWM3/RemaTxNum[22]_keep ;
  wire \PWM3/RemaTxNum[23]_keep ;
  wire \PWM3/RemaTxNum[2]_keep ;
  wire \PWM3/RemaTxNum[3]_keep ;
  wire \PWM3/RemaTxNum[4]_keep ;
  wire \PWM3/RemaTxNum[5]_keep ;
  wire \PWM3/RemaTxNum[6]_keep ;
  wire \PWM3/RemaTxNum[7]_keep ;
  wire \PWM3/RemaTxNum[8]_keep ;
  wire \PWM3/RemaTxNum[9]_keep ;
  wire \PWM3/dir_keep ;
  wire \PWM3/mux3_b0_sel_is_3_o ;
  wire \PWM3/n0 ;
  wire \PWM3/n1 ;
  wire \PWM3/n10 ;
  wire \PWM3/n11 ;
  wire \PWM3/n17 ;
  wire \PWM3/n17_neg ;
  wire \PWM3/n18 ;
  wire \PWM3/n24 ;
  wire \PWM3/n25 ;
  wire \PWM3/n25_neg ;
  wire \PWM3/n32 ;
  wire \PWM3/n4 ;
  wire \PWM3/n4_neg ;
  wire \PWM3/n5 ;
  wire \PWM3/n6 ;
  wire \PWM3/n6_neg ;
  wire \PWM3/n8 ;
  wire \PWM3/n9 ;
  wire \PWM3/pnumr[0]_keep ;
  wire \PWM3/pnumr[10]_keep ;
  wire \PWM3/pnumr[11]_keep ;
  wire \PWM3/pnumr[12]_keep ;
  wire \PWM3/pnumr[13]_keep ;
  wire \PWM3/pnumr[14]_keep ;
  wire \PWM3/pnumr[15]_keep ;
  wire \PWM3/pnumr[16]_keep ;
  wire \PWM3/pnumr[17]_keep ;
  wire \PWM3/pnumr[18]_keep ;
  wire \PWM3/pnumr[19]_keep ;
  wire \PWM3/pnumr[1]_keep ;
  wire \PWM3/pnumr[20]_keep ;
  wire \PWM3/pnumr[21]_keep ;
  wire \PWM3/pnumr[22]_keep ;
  wire \PWM3/pnumr[23]_keep ;
  wire \PWM3/pnumr[24]_keep ;
  wire \PWM3/pnumr[25]_keep ;
  wire \PWM3/pnumr[26]_keep ;
  wire \PWM3/pnumr[27]_keep ;
  wire \PWM3/pnumr[28]_keep ;
  wire \PWM3/pnumr[29]_keep ;
  wire \PWM3/pnumr[2]_keep ;
  wire \PWM3/pnumr[30]_keep ;
  wire \PWM3/pnumr[31]_keep ;
  wire \PWM3/pnumr[3]_keep ;
  wire \PWM3/pnumr[4]_keep ;
  wire \PWM3/pnumr[5]_keep ;
  wire \PWM3/pnumr[6]_keep ;
  wire \PWM3/pnumr[7]_keep ;
  wire \PWM3/pnumr[8]_keep ;
  wire \PWM3/pnumr[9]_keep ;
  wire \PWM3/pwm_keep ;
  wire \PWM3/stopreq ;  // src/OnePWM.v(14)
  wire \PWM3/stopreq_keep ;
  wire \PWM3/u14_sel_is_1_o ;
  wire \PWM3/u17_sel_is_1_o ;
  wire \PWM3/u17_sel_is_1_o_neg ;
  wire \PWM3/u18_sel_is_0_o ;
  wire \PWM3/u8_sel_is_0_o ;
  wire \PWM4/RemaTxNum[0]_keep ;
  wire \PWM4/RemaTxNum[10]_keep ;
  wire \PWM4/RemaTxNum[11]_keep ;
  wire \PWM4/RemaTxNum[12]_keep ;
  wire \PWM4/RemaTxNum[13]_keep ;
  wire \PWM4/RemaTxNum[14]_keep ;
  wire \PWM4/RemaTxNum[15]_keep ;
  wire \PWM4/RemaTxNum[16]_keep ;
  wire \PWM4/RemaTxNum[17]_keep ;
  wire \PWM4/RemaTxNum[18]_keep ;
  wire \PWM4/RemaTxNum[19]_keep ;
  wire \PWM4/RemaTxNum[1]_keep ;
  wire \PWM4/RemaTxNum[20]_keep ;
  wire \PWM4/RemaTxNum[21]_keep ;
  wire \PWM4/RemaTxNum[22]_keep ;
  wire \PWM4/RemaTxNum[23]_keep ;
  wire \PWM4/RemaTxNum[2]_keep ;
  wire \PWM4/RemaTxNum[3]_keep ;
  wire \PWM4/RemaTxNum[4]_keep ;
  wire \PWM4/RemaTxNum[5]_keep ;
  wire \PWM4/RemaTxNum[6]_keep ;
  wire \PWM4/RemaTxNum[7]_keep ;
  wire \PWM4/RemaTxNum[8]_keep ;
  wire \PWM4/RemaTxNum[9]_keep ;
  wire \PWM4/dir_keep ;
  wire \PWM4/mux3_b0_sel_is_3_o ;
  wire \PWM4/n0 ;
  wire \PWM4/n1 ;
  wire \PWM4/n10 ;
  wire \PWM4/n11 ;
  wire \PWM4/n17 ;
  wire \PWM4/n17_neg ;
  wire \PWM4/n18 ;
  wire \PWM4/n24 ;
  wire \PWM4/n25 ;
  wire \PWM4/n25_neg ;
  wire \PWM4/n32 ;
  wire \PWM4/n4 ;
  wire \PWM4/n4_neg ;
  wire \PWM4/n5 ;
  wire \PWM4/n6 ;
  wire \PWM4/n6_neg ;
  wire \PWM4/n8 ;
  wire \PWM4/n9 ;
  wire \PWM4/pnumr[0]_keep ;
  wire \PWM4/pnumr[10]_keep ;
  wire \PWM4/pnumr[11]_keep ;
  wire \PWM4/pnumr[12]_keep ;
  wire \PWM4/pnumr[13]_keep ;
  wire \PWM4/pnumr[14]_keep ;
  wire \PWM4/pnumr[15]_keep ;
  wire \PWM4/pnumr[16]_keep ;
  wire \PWM4/pnumr[17]_keep ;
  wire \PWM4/pnumr[18]_keep ;
  wire \PWM4/pnumr[19]_keep ;
  wire \PWM4/pnumr[1]_keep ;
  wire \PWM4/pnumr[20]_keep ;
  wire \PWM4/pnumr[21]_keep ;
  wire \PWM4/pnumr[22]_keep ;
  wire \PWM4/pnumr[23]_keep ;
  wire \PWM4/pnumr[24]_keep ;
  wire \PWM4/pnumr[25]_keep ;
  wire \PWM4/pnumr[26]_keep ;
  wire \PWM4/pnumr[27]_keep ;
  wire \PWM4/pnumr[28]_keep ;
  wire \PWM4/pnumr[29]_keep ;
  wire \PWM4/pnumr[2]_keep ;
  wire \PWM4/pnumr[30]_keep ;
  wire \PWM4/pnumr[31]_keep ;
  wire \PWM4/pnumr[3]_keep ;
  wire \PWM4/pnumr[4]_keep ;
  wire \PWM4/pnumr[5]_keep ;
  wire \PWM4/pnumr[6]_keep ;
  wire \PWM4/pnumr[7]_keep ;
  wire \PWM4/pnumr[8]_keep ;
  wire \PWM4/pnumr[9]_keep ;
  wire \PWM4/pwm_keep ;
  wire \PWM4/stopreq ;  // src/OnePWM.v(14)
  wire \PWM4/stopreq_keep ;
  wire \PWM4/u14_sel_is_1_o ;
  wire \PWM4/u17_sel_is_1_o ;
  wire \PWM4/u17_sel_is_1_o_neg ;
  wire \PWM4/u18_sel_is_0_o ;
  wire \PWM4/u8_sel_is_0_o ;
  wire \PWM5/RemaTxNum[0]_keep ;
  wire \PWM5/RemaTxNum[10]_keep ;
  wire \PWM5/RemaTxNum[11]_keep ;
  wire \PWM5/RemaTxNum[12]_keep ;
  wire \PWM5/RemaTxNum[13]_keep ;
  wire \PWM5/RemaTxNum[14]_keep ;
  wire \PWM5/RemaTxNum[15]_keep ;
  wire \PWM5/RemaTxNum[16]_keep ;
  wire \PWM5/RemaTxNum[17]_keep ;
  wire \PWM5/RemaTxNum[18]_keep ;
  wire \PWM5/RemaTxNum[19]_keep ;
  wire \PWM5/RemaTxNum[1]_keep ;
  wire \PWM5/RemaTxNum[20]_keep ;
  wire \PWM5/RemaTxNum[21]_keep ;
  wire \PWM5/RemaTxNum[22]_keep ;
  wire \PWM5/RemaTxNum[23]_keep ;
  wire \PWM5/RemaTxNum[2]_keep ;
  wire \PWM5/RemaTxNum[3]_keep ;
  wire \PWM5/RemaTxNum[4]_keep ;
  wire \PWM5/RemaTxNum[5]_keep ;
  wire \PWM5/RemaTxNum[6]_keep ;
  wire \PWM5/RemaTxNum[7]_keep ;
  wire \PWM5/RemaTxNum[8]_keep ;
  wire \PWM5/RemaTxNum[9]_keep ;
  wire \PWM5/dir_keep ;
  wire \PWM5/mux3_b0_sel_is_3_o ;
  wire \PWM5/n0 ;
  wire \PWM5/n1 ;
  wire \PWM5/n10 ;
  wire \PWM5/n11 ;
  wire \PWM5/n17 ;
  wire \PWM5/n17_neg ;
  wire \PWM5/n18 ;
  wire \PWM5/n24 ;
  wire \PWM5/n25 ;
  wire \PWM5/n25_neg ;
  wire \PWM5/n32 ;
  wire \PWM5/n4 ;
  wire \PWM5/n4_neg ;
  wire \PWM5/n5 ;
  wire \PWM5/n6 ;
  wire \PWM5/n6_neg ;
  wire \PWM5/n8 ;
  wire \PWM5/n9 ;
  wire \PWM5/pnumr[0]_keep ;
  wire \PWM5/pnumr[10]_keep ;
  wire \PWM5/pnumr[11]_keep ;
  wire \PWM5/pnumr[12]_keep ;
  wire \PWM5/pnumr[13]_keep ;
  wire \PWM5/pnumr[14]_keep ;
  wire \PWM5/pnumr[15]_keep ;
  wire \PWM5/pnumr[16]_keep ;
  wire \PWM5/pnumr[17]_keep ;
  wire \PWM5/pnumr[18]_keep ;
  wire \PWM5/pnumr[19]_keep ;
  wire \PWM5/pnumr[1]_keep ;
  wire \PWM5/pnumr[20]_keep ;
  wire \PWM5/pnumr[21]_keep ;
  wire \PWM5/pnumr[22]_keep ;
  wire \PWM5/pnumr[23]_keep ;
  wire \PWM5/pnumr[24]_keep ;
  wire \PWM5/pnumr[25]_keep ;
  wire \PWM5/pnumr[26]_keep ;
  wire \PWM5/pnumr[27]_keep ;
  wire \PWM5/pnumr[28]_keep ;
  wire \PWM5/pnumr[29]_keep ;
  wire \PWM5/pnumr[2]_keep ;
  wire \PWM5/pnumr[30]_keep ;
  wire \PWM5/pnumr[31]_keep ;
  wire \PWM5/pnumr[3]_keep ;
  wire \PWM5/pnumr[4]_keep ;
  wire \PWM5/pnumr[5]_keep ;
  wire \PWM5/pnumr[6]_keep ;
  wire \PWM5/pnumr[7]_keep ;
  wire \PWM5/pnumr[8]_keep ;
  wire \PWM5/pnumr[9]_keep ;
  wire \PWM5/pwm_keep ;
  wire \PWM5/stopreq ;  // src/OnePWM.v(14)
  wire \PWM5/stopreq_keep ;
  wire \PWM5/u14_sel_is_1_o ;
  wire \PWM5/u17_sel_is_1_o ;
  wire \PWM5/u17_sel_is_1_o_neg ;
  wire \PWM5/u18_sel_is_0_o ;
  wire \PWM5/u8_sel_is_0_o ;
  wire \PWM6/RemaTxNum[0]_keep ;
  wire \PWM6/RemaTxNum[10]_keep ;
  wire \PWM6/RemaTxNum[11]_keep ;
  wire \PWM6/RemaTxNum[12]_keep ;
  wire \PWM6/RemaTxNum[13]_keep ;
  wire \PWM6/RemaTxNum[14]_keep ;
  wire \PWM6/RemaTxNum[15]_keep ;
  wire \PWM6/RemaTxNum[16]_keep ;
  wire \PWM6/RemaTxNum[17]_keep ;
  wire \PWM6/RemaTxNum[18]_keep ;
  wire \PWM6/RemaTxNum[19]_keep ;
  wire \PWM6/RemaTxNum[1]_keep ;
  wire \PWM6/RemaTxNum[20]_keep ;
  wire \PWM6/RemaTxNum[21]_keep ;
  wire \PWM6/RemaTxNum[22]_keep ;
  wire \PWM6/RemaTxNum[23]_keep ;
  wire \PWM6/RemaTxNum[2]_keep ;
  wire \PWM6/RemaTxNum[3]_keep ;
  wire \PWM6/RemaTxNum[4]_keep ;
  wire \PWM6/RemaTxNum[5]_keep ;
  wire \PWM6/RemaTxNum[6]_keep ;
  wire \PWM6/RemaTxNum[7]_keep ;
  wire \PWM6/RemaTxNum[8]_keep ;
  wire \PWM6/RemaTxNum[9]_keep ;
  wire \PWM6/dir_keep ;
  wire \PWM6/mux3_b0_sel_is_3_o ;
  wire \PWM6/n0 ;
  wire \PWM6/n1 ;
  wire \PWM6/n10 ;
  wire \PWM6/n11 ;
  wire \PWM6/n17 ;
  wire \PWM6/n17_neg ;
  wire \PWM6/n18 ;
  wire \PWM6/n24 ;
  wire \PWM6/n25 ;
  wire \PWM6/n25_neg ;
  wire \PWM6/n32 ;
  wire \PWM6/n4 ;
  wire \PWM6/n4_neg ;
  wire \PWM6/n5 ;
  wire \PWM6/n6 ;
  wire \PWM6/n6_neg ;
  wire \PWM6/n8 ;
  wire \PWM6/n9 ;
  wire \PWM6/pnumr[0]_keep ;
  wire \PWM6/pnumr[10]_keep ;
  wire \PWM6/pnumr[11]_keep ;
  wire \PWM6/pnumr[12]_keep ;
  wire \PWM6/pnumr[13]_keep ;
  wire \PWM6/pnumr[14]_keep ;
  wire \PWM6/pnumr[15]_keep ;
  wire \PWM6/pnumr[16]_keep ;
  wire \PWM6/pnumr[17]_keep ;
  wire \PWM6/pnumr[18]_keep ;
  wire \PWM6/pnumr[19]_keep ;
  wire \PWM6/pnumr[1]_keep ;
  wire \PWM6/pnumr[20]_keep ;
  wire \PWM6/pnumr[21]_keep ;
  wire \PWM6/pnumr[22]_keep ;
  wire \PWM6/pnumr[23]_keep ;
  wire \PWM6/pnumr[24]_keep ;
  wire \PWM6/pnumr[25]_keep ;
  wire \PWM6/pnumr[26]_keep ;
  wire \PWM6/pnumr[27]_keep ;
  wire \PWM6/pnumr[28]_keep ;
  wire \PWM6/pnumr[29]_keep ;
  wire \PWM6/pnumr[2]_keep ;
  wire \PWM6/pnumr[30]_keep ;
  wire \PWM6/pnumr[31]_keep ;
  wire \PWM6/pnumr[3]_keep ;
  wire \PWM6/pnumr[4]_keep ;
  wire \PWM6/pnumr[5]_keep ;
  wire \PWM6/pnumr[6]_keep ;
  wire \PWM6/pnumr[7]_keep ;
  wire \PWM6/pnumr[8]_keep ;
  wire \PWM6/pnumr[9]_keep ;
  wire \PWM6/pwm_keep ;
  wire \PWM6/stopreq ;  // src/OnePWM.v(14)
  wire \PWM6/stopreq_keep ;
  wire \PWM6/u14_sel_is_1_o ;
  wire \PWM6/u17_sel_is_1_o ;
  wire \PWM6/u17_sel_is_1_o_neg ;
  wire \PWM6/u18_sel_is_0_o ;
  wire \PWM6/u8_sel_is_0_o ;
  wire \PWM7/RemaTxNum[0]_keep ;
  wire \PWM7/RemaTxNum[10]_keep ;
  wire \PWM7/RemaTxNum[11]_keep ;
  wire \PWM7/RemaTxNum[12]_keep ;
  wire \PWM7/RemaTxNum[13]_keep ;
  wire \PWM7/RemaTxNum[14]_keep ;
  wire \PWM7/RemaTxNum[15]_keep ;
  wire \PWM7/RemaTxNum[16]_keep ;
  wire \PWM7/RemaTxNum[17]_keep ;
  wire \PWM7/RemaTxNum[18]_keep ;
  wire \PWM7/RemaTxNum[19]_keep ;
  wire \PWM7/RemaTxNum[1]_keep ;
  wire \PWM7/RemaTxNum[20]_keep ;
  wire \PWM7/RemaTxNum[21]_keep ;
  wire \PWM7/RemaTxNum[22]_keep ;
  wire \PWM7/RemaTxNum[23]_keep ;
  wire \PWM7/RemaTxNum[2]_keep ;
  wire \PWM7/RemaTxNum[3]_keep ;
  wire \PWM7/RemaTxNum[4]_keep ;
  wire \PWM7/RemaTxNum[5]_keep ;
  wire \PWM7/RemaTxNum[6]_keep ;
  wire \PWM7/RemaTxNum[7]_keep ;
  wire \PWM7/RemaTxNum[8]_keep ;
  wire \PWM7/RemaTxNum[9]_keep ;
  wire \PWM7/dir_keep ;
  wire \PWM7/mux3_b0_sel_is_3_o ;
  wire \PWM7/n0 ;
  wire \PWM7/n1 ;
  wire \PWM7/n10 ;
  wire \PWM7/n11 ;
  wire \PWM7/n17 ;
  wire \PWM7/n17_neg ;
  wire \PWM7/n18 ;
  wire \PWM7/n24 ;
  wire \PWM7/n25 ;
  wire \PWM7/n25_neg ;
  wire \PWM7/n32 ;
  wire \PWM7/n4 ;
  wire \PWM7/n4_neg ;
  wire \PWM7/n5 ;
  wire \PWM7/n6 ;
  wire \PWM7/n6_neg ;
  wire \PWM7/n8 ;
  wire \PWM7/n9 ;
  wire \PWM7/pnumr[0]_keep ;
  wire \PWM7/pnumr[10]_keep ;
  wire \PWM7/pnumr[11]_keep ;
  wire \PWM7/pnumr[12]_keep ;
  wire \PWM7/pnumr[13]_keep ;
  wire \PWM7/pnumr[14]_keep ;
  wire \PWM7/pnumr[15]_keep ;
  wire \PWM7/pnumr[16]_keep ;
  wire \PWM7/pnumr[17]_keep ;
  wire \PWM7/pnumr[18]_keep ;
  wire \PWM7/pnumr[19]_keep ;
  wire \PWM7/pnumr[1]_keep ;
  wire \PWM7/pnumr[20]_keep ;
  wire \PWM7/pnumr[21]_keep ;
  wire \PWM7/pnumr[22]_keep ;
  wire \PWM7/pnumr[23]_keep ;
  wire \PWM7/pnumr[24]_keep ;
  wire \PWM7/pnumr[25]_keep ;
  wire \PWM7/pnumr[26]_keep ;
  wire \PWM7/pnumr[27]_keep ;
  wire \PWM7/pnumr[28]_keep ;
  wire \PWM7/pnumr[29]_keep ;
  wire \PWM7/pnumr[2]_keep ;
  wire \PWM7/pnumr[30]_keep ;
  wire \PWM7/pnumr[31]_keep ;
  wire \PWM7/pnumr[3]_keep ;
  wire \PWM7/pnumr[4]_keep ;
  wire \PWM7/pnumr[5]_keep ;
  wire \PWM7/pnumr[6]_keep ;
  wire \PWM7/pnumr[7]_keep ;
  wire \PWM7/pnumr[8]_keep ;
  wire \PWM7/pnumr[9]_keep ;
  wire \PWM7/pwm_keep ;
  wire \PWM7/stopreq ;  // src/OnePWM.v(14)
  wire \PWM7/stopreq_keep ;
  wire \PWM7/u14_sel_is_1_o ;
  wire \PWM7/u17_sel_is_1_o ;
  wire \PWM7/u17_sel_is_1_o_neg ;
  wire \PWM7/u18_sel_is_0_o ;
  wire \PWM7/u8_sel_is_0_o ;
  wire \PWM8/RemaTxNum[0]_keep ;
  wire \PWM8/RemaTxNum[10]_keep ;
  wire \PWM8/RemaTxNum[11]_keep ;
  wire \PWM8/RemaTxNum[12]_keep ;
  wire \PWM8/RemaTxNum[13]_keep ;
  wire \PWM8/RemaTxNum[14]_keep ;
  wire \PWM8/RemaTxNum[15]_keep ;
  wire \PWM8/RemaTxNum[16]_keep ;
  wire \PWM8/RemaTxNum[17]_keep ;
  wire \PWM8/RemaTxNum[18]_keep ;
  wire \PWM8/RemaTxNum[19]_keep ;
  wire \PWM8/RemaTxNum[1]_keep ;
  wire \PWM8/RemaTxNum[20]_keep ;
  wire \PWM8/RemaTxNum[21]_keep ;
  wire \PWM8/RemaTxNum[22]_keep ;
  wire \PWM8/RemaTxNum[23]_keep ;
  wire \PWM8/RemaTxNum[2]_keep ;
  wire \PWM8/RemaTxNum[3]_keep ;
  wire \PWM8/RemaTxNum[4]_keep ;
  wire \PWM8/RemaTxNum[5]_keep ;
  wire \PWM8/RemaTxNum[6]_keep ;
  wire \PWM8/RemaTxNum[7]_keep ;
  wire \PWM8/RemaTxNum[8]_keep ;
  wire \PWM8/RemaTxNum[9]_keep ;
  wire \PWM8/dir_keep ;
  wire \PWM8/mux3_b0_sel_is_3_o ;
  wire \PWM8/n0 ;
  wire \PWM8/n1 ;
  wire \PWM8/n10 ;
  wire \PWM8/n11 ;
  wire \PWM8/n17 ;
  wire \PWM8/n17_neg ;
  wire \PWM8/n18 ;
  wire \PWM8/n24 ;
  wire \PWM8/n25 ;
  wire \PWM8/n25_neg ;
  wire \PWM8/n32 ;
  wire \PWM8/n4 ;
  wire \PWM8/n4_neg ;
  wire \PWM8/n5 ;
  wire \PWM8/n6 ;
  wire \PWM8/n6_neg ;
  wire \PWM8/n8 ;
  wire \PWM8/n9 ;
  wire \PWM8/pnumr[0]_keep ;
  wire \PWM8/pnumr[10]_keep ;
  wire \PWM8/pnumr[11]_keep ;
  wire \PWM8/pnumr[12]_keep ;
  wire \PWM8/pnumr[13]_keep ;
  wire \PWM8/pnumr[14]_keep ;
  wire \PWM8/pnumr[15]_keep ;
  wire \PWM8/pnumr[16]_keep ;
  wire \PWM8/pnumr[17]_keep ;
  wire \PWM8/pnumr[18]_keep ;
  wire \PWM8/pnumr[19]_keep ;
  wire \PWM8/pnumr[1]_keep ;
  wire \PWM8/pnumr[20]_keep ;
  wire \PWM8/pnumr[21]_keep ;
  wire \PWM8/pnumr[22]_keep ;
  wire \PWM8/pnumr[23]_keep ;
  wire \PWM8/pnumr[24]_keep ;
  wire \PWM8/pnumr[25]_keep ;
  wire \PWM8/pnumr[26]_keep ;
  wire \PWM8/pnumr[27]_keep ;
  wire \PWM8/pnumr[28]_keep ;
  wire \PWM8/pnumr[29]_keep ;
  wire \PWM8/pnumr[2]_keep ;
  wire \PWM8/pnumr[30]_keep ;
  wire \PWM8/pnumr[31]_keep ;
  wire \PWM8/pnumr[3]_keep ;
  wire \PWM8/pnumr[4]_keep ;
  wire \PWM8/pnumr[5]_keep ;
  wire \PWM8/pnumr[6]_keep ;
  wire \PWM8/pnumr[7]_keep ;
  wire \PWM8/pnumr[8]_keep ;
  wire \PWM8/pnumr[9]_keep ;
  wire \PWM8/pwm_keep ;
  wire \PWM8/stopreq ;  // src/OnePWM.v(14)
  wire \PWM8/stopreq_keep ;
  wire \PWM8/u14_sel_is_1_o ;
  wire \PWM8/u17_sel_is_1_o ;
  wire \PWM8/u17_sel_is_1_o_neg ;
  wire \PWM8/u18_sel_is_0_o ;
  wire \PWM8/u8_sel_is_0_o ;
  wire \PWM9/RemaTxNum[0]_keep ;
  wire \PWM9/RemaTxNum[10]_keep ;
  wire \PWM9/RemaTxNum[11]_keep ;
  wire \PWM9/RemaTxNum[12]_keep ;
  wire \PWM9/RemaTxNum[13]_keep ;
  wire \PWM9/RemaTxNum[14]_keep ;
  wire \PWM9/RemaTxNum[15]_keep ;
  wire \PWM9/RemaTxNum[16]_keep ;
  wire \PWM9/RemaTxNum[17]_keep ;
  wire \PWM9/RemaTxNum[18]_keep ;
  wire \PWM9/RemaTxNum[19]_keep ;
  wire \PWM9/RemaTxNum[1]_keep ;
  wire \PWM9/RemaTxNum[20]_keep ;
  wire \PWM9/RemaTxNum[21]_keep ;
  wire \PWM9/RemaTxNum[22]_keep ;
  wire \PWM9/RemaTxNum[23]_keep ;
  wire \PWM9/RemaTxNum[2]_keep ;
  wire \PWM9/RemaTxNum[3]_keep ;
  wire \PWM9/RemaTxNum[4]_keep ;
  wire \PWM9/RemaTxNum[5]_keep ;
  wire \PWM9/RemaTxNum[6]_keep ;
  wire \PWM9/RemaTxNum[7]_keep ;
  wire \PWM9/RemaTxNum[8]_keep ;
  wire \PWM9/RemaTxNum[9]_keep ;
  wire \PWM9/dir_keep ;
  wire \PWM9/mux3_b0_sel_is_3_o ;
  wire \PWM9/n0 ;
  wire \PWM9/n1 ;
  wire \PWM9/n10 ;
  wire \PWM9/n11 ;
  wire \PWM9/n17 ;
  wire \PWM9/n17_neg ;
  wire \PWM9/n18 ;
  wire \PWM9/n24 ;
  wire \PWM9/n25 ;
  wire \PWM9/n25_neg ;
  wire \PWM9/n32 ;
  wire \PWM9/n4 ;
  wire \PWM9/n4_neg ;
  wire \PWM9/n5 ;
  wire \PWM9/n6 ;
  wire \PWM9/n6_neg ;
  wire \PWM9/n8 ;
  wire \PWM9/n9 ;
  wire \PWM9/pnumr[0]_keep ;
  wire \PWM9/pnumr[10]_keep ;
  wire \PWM9/pnumr[11]_keep ;
  wire \PWM9/pnumr[12]_keep ;
  wire \PWM9/pnumr[13]_keep ;
  wire \PWM9/pnumr[14]_keep ;
  wire \PWM9/pnumr[15]_keep ;
  wire \PWM9/pnumr[16]_keep ;
  wire \PWM9/pnumr[17]_keep ;
  wire \PWM9/pnumr[18]_keep ;
  wire \PWM9/pnumr[19]_keep ;
  wire \PWM9/pnumr[1]_keep ;
  wire \PWM9/pnumr[20]_keep ;
  wire \PWM9/pnumr[21]_keep ;
  wire \PWM9/pnumr[22]_keep ;
  wire \PWM9/pnumr[23]_keep ;
  wire \PWM9/pnumr[24]_keep ;
  wire \PWM9/pnumr[25]_keep ;
  wire \PWM9/pnumr[26]_keep ;
  wire \PWM9/pnumr[27]_keep ;
  wire \PWM9/pnumr[28]_keep ;
  wire \PWM9/pnumr[29]_keep ;
  wire \PWM9/pnumr[2]_keep ;
  wire \PWM9/pnumr[30]_keep ;
  wire \PWM9/pnumr[31]_keep ;
  wire \PWM9/pnumr[3]_keep ;
  wire \PWM9/pnumr[4]_keep ;
  wire \PWM9/pnumr[5]_keep ;
  wire \PWM9/pnumr[6]_keep ;
  wire \PWM9/pnumr[7]_keep ;
  wire \PWM9/pnumr[8]_keep ;
  wire \PWM9/pnumr[9]_keep ;
  wire \PWM9/pwm_keep ;
  wire \PWM9/stopreq ;  // src/OnePWM.v(14)
  wire \PWM9/stopreq_keep ;
  wire \PWM9/u14_sel_is_1_o ;
  wire \PWM9/u17_sel_is_1_o ;
  wire \PWM9/u17_sel_is_1_o_neg ;
  wire \PWM9/u18_sel_is_0_o ;
  wire \PWM9/u8_sel_is_0_o ;
  wire \PWMA/RemaTxNum[0]_keep ;
  wire \PWMA/RemaTxNum[10]_keep ;
  wire \PWMA/RemaTxNum[11]_keep ;
  wire \PWMA/RemaTxNum[12]_keep ;
  wire \PWMA/RemaTxNum[13]_keep ;
  wire \PWMA/RemaTxNum[14]_keep ;
  wire \PWMA/RemaTxNum[15]_keep ;
  wire \PWMA/RemaTxNum[16]_keep ;
  wire \PWMA/RemaTxNum[17]_keep ;
  wire \PWMA/RemaTxNum[18]_keep ;
  wire \PWMA/RemaTxNum[19]_keep ;
  wire \PWMA/RemaTxNum[1]_keep ;
  wire \PWMA/RemaTxNum[20]_keep ;
  wire \PWMA/RemaTxNum[21]_keep ;
  wire \PWMA/RemaTxNum[22]_keep ;
  wire \PWMA/RemaTxNum[23]_keep ;
  wire \PWMA/RemaTxNum[2]_keep ;
  wire \PWMA/RemaTxNum[3]_keep ;
  wire \PWMA/RemaTxNum[4]_keep ;
  wire \PWMA/RemaTxNum[5]_keep ;
  wire \PWMA/RemaTxNum[6]_keep ;
  wire \PWMA/RemaTxNum[7]_keep ;
  wire \PWMA/RemaTxNum[8]_keep ;
  wire \PWMA/RemaTxNum[9]_keep ;
  wire \PWMA/dir_keep ;
  wire \PWMA/mux3_b0_sel_is_3_o ;
  wire \PWMA/n0 ;
  wire \PWMA/n1 ;
  wire \PWMA/n10 ;
  wire \PWMA/n11 ;
  wire \PWMA/n17 ;
  wire \PWMA/n17_neg ;
  wire \PWMA/n18 ;
  wire \PWMA/n24 ;
  wire \PWMA/n25 ;
  wire \PWMA/n25_neg ;
  wire \PWMA/n32 ;
  wire \PWMA/n4 ;
  wire \PWMA/n4_neg ;
  wire \PWMA/n5 ;
  wire \PWMA/n6 ;
  wire \PWMA/n6_neg ;
  wire \PWMA/n8 ;
  wire \PWMA/n9 ;
  wire \PWMA/pnumr[0]_keep ;
  wire \PWMA/pnumr[10]_keep ;
  wire \PWMA/pnumr[11]_keep ;
  wire \PWMA/pnumr[12]_keep ;
  wire \PWMA/pnumr[13]_keep ;
  wire \PWMA/pnumr[14]_keep ;
  wire \PWMA/pnumr[15]_keep ;
  wire \PWMA/pnumr[16]_keep ;
  wire \PWMA/pnumr[17]_keep ;
  wire \PWMA/pnumr[18]_keep ;
  wire \PWMA/pnumr[19]_keep ;
  wire \PWMA/pnumr[1]_keep ;
  wire \PWMA/pnumr[20]_keep ;
  wire \PWMA/pnumr[21]_keep ;
  wire \PWMA/pnumr[22]_keep ;
  wire \PWMA/pnumr[23]_keep ;
  wire \PWMA/pnumr[24]_keep ;
  wire \PWMA/pnumr[25]_keep ;
  wire \PWMA/pnumr[26]_keep ;
  wire \PWMA/pnumr[27]_keep ;
  wire \PWMA/pnumr[28]_keep ;
  wire \PWMA/pnumr[29]_keep ;
  wire \PWMA/pnumr[2]_keep ;
  wire \PWMA/pnumr[30]_keep ;
  wire \PWMA/pnumr[31]_keep ;
  wire \PWMA/pnumr[3]_keep ;
  wire \PWMA/pnumr[4]_keep ;
  wire \PWMA/pnumr[5]_keep ;
  wire \PWMA/pnumr[6]_keep ;
  wire \PWMA/pnumr[7]_keep ;
  wire \PWMA/pnumr[8]_keep ;
  wire \PWMA/pnumr[9]_keep ;
  wire \PWMA/pwm_keep ;
  wire \PWMA/stopreq ;  // src/OnePWM.v(14)
  wire \PWMA/stopreq_keep ;
  wire \PWMA/u14_sel_is_1_o ;
  wire \PWMA/u17_sel_is_1_o ;
  wire \PWMA/u17_sel_is_1_o_neg ;
  wire \PWMA/u18_sel_is_0_o ;
  wire \PWMA/u8_sel_is_0_o ;
  wire \PWMB/RemaTxNum[0]_keep ;
  wire \PWMB/RemaTxNum[10]_keep ;
  wire \PWMB/RemaTxNum[11]_keep ;
  wire \PWMB/RemaTxNum[12]_keep ;
  wire \PWMB/RemaTxNum[13]_keep ;
  wire \PWMB/RemaTxNum[14]_keep ;
  wire \PWMB/RemaTxNum[15]_keep ;
  wire \PWMB/RemaTxNum[16]_keep ;
  wire \PWMB/RemaTxNum[17]_keep ;
  wire \PWMB/RemaTxNum[18]_keep ;
  wire \PWMB/RemaTxNum[19]_keep ;
  wire \PWMB/RemaTxNum[1]_keep ;
  wire \PWMB/RemaTxNum[20]_keep ;
  wire \PWMB/RemaTxNum[21]_keep ;
  wire \PWMB/RemaTxNum[22]_keep ;
  wire \PWMB/RemaTxNum[23]_keep ;
  wire \PWMB/RemaTxNum[2]_keep ;
  wire \PWMB/RemaTxNum[3]_keep ;
  wire \PWMB/RemaTxNum[4]_keep ;
  wire \PWMB/RemaTxNum[5]_keep ;
  wire \PWMB/RemaTxNum[6]_keep ;
  wire \PWMB/RemaTxNum[7]_keep ;
  wire \PWMB/RemaTxNum[8]_keep ;
  wire \PWMB/RemaTxNum[9]_keep ;
  wire \PWMB/dir_keep ;
  wire \PWMB/mux3_b0_sel_is_3_o ;
  wire \PWMB/n0 ;
  wire \PWMB/n1 ;
  wire \PWMB/n10 ;
  wire \PWMB/n11 ;
  wire \PWMB/n17 ;
  wire \PWMB/n17_neg ;
  wire \PWMB/n18 ;
  wire \PWMB/n24 ;
  wire \PWMB/n25 ;
  wire \PWMB/n25_neg ;
  wire \PWMB/n32 ;
  wire \PWMB/n4 ;
  wire \PWMB/n4_neg ;
  wire \PWMB/n5 ;
  wire \PWMB/n6 ;
  wire \PWMB/n6_neg ;
  wire \PWMB/n8 ;
  wire \PWMB/n9 ;
  wire \PWMB/pnumr[0]_keep ;
  wire \PWMB/pnumr[10]_keep ;
  wire \PWMB/pnumr[11]_keep ;
  wire \PWMB/pnumr[12]_keep ;
  wire \PWMB/pnumr[13]_keep ;
  wire \PWMB/pnumr[14]_keep ;
  wire \PWMB/pnumr[15]_keep ;
  wire \PWMB/pnumr[16]_keep ;
  wire \PWMB/pnumr[17]_keep ;
  wire \PWMB/pnumr[18]_keep ;
  wire \PWMB/pnumr[19]_keep ;
  wire \PWMB/pnumr[1]_keep ;
  wire \PWMB/pnumr[20]_keep ;
  wire \PWMB/pnumr[21]_keep ;
  wire \PWMB/pnumr[22]_keep ;
  wire \PWMB/pnumr[23]_keep ;
  wire \PWMB/pnumr[24]_keep ;
  wire \PWMB/pnumr[25]_keep ;
  wire \PWMB/pnumr[26]_keep ;
  wire \PWMB/pnumr[27]_keep ;
  wire \PWMB/pnumr[28]_keep ;
  wire \PWMB/pnumr[29]_keep ;
  wire \PWMB/pnumr[2]_keep ;
  wire \PWMB/pnumr[30]_keep ;
  wire \PWMB/pnumr[31]_keep ;
  wire \PWMB/pnumr[3]_keep ;
  wire \PWMB/pnumr[4]_keep ;
  wire \PWMB/pnumr[5]_keep ;
  wire \PWMB/pnumr[6]_keep ;
  wire \PWMB/pnumr[7]_keep ;
  wire \PWMB/pnumr[8]_keep ;
  wire \PWMB/pnumr[9]_keep ;
  wire \PWMB/pwm_keep ;
  wire \PWMB/stopreq ;  // src/OnePWM.v(14)
  wire \PWMB/stopreq_keep ;
  wire \PWMB/u14_sel_is_1_o ;
  wire \PWMB/u17_sel_is_1_o ;
  wire \PWMB/u17_sel_is_1_o_neg ;
  wire \PWMB/u18_sel_is_0_o ;
  wire \PWMB/u8_sel_is_0_o ;
  wire \PWMC/RemaTxNum[0]_keep ;
  wire \PWMC/RemaTxNum[10]_keep ;
  wire \PWMC/RemaTxNum[11]_keep ;
  wire \PWMC/RemaTxNum[12]_keep ;
  wire \PWMC/RemaTxNum[13]_keep ;
  wire \PWMC/RemaTxNum[14]_keep ;
  wire \PWMC/RemaTxNum[15]_keep ;
  wire \PWMC/RemaTxNum[16]_keep ;
  wire \PWMC/RemaTxNum[17]_keep ;
  wire \PWMC/RemaTxNum[18]_keep ;
  wire \PWMC/RemaTxNum[19]_keep ;
  wire \PWMC/RemaTxNum[1]_keep ;
  wire \PWMC/RemaTxNum[20]_keep ;
  wire \PWMC/RemaTxNum[21]_keep ;
  wire \PWMC/RemaTxNum[22]_keep ;
  wire \PWMC/RemaTxNum[23]_keep ;
  wire \PWMC/RemaTxNum[2]_keep ;
  wire \PWMC/RemaTxNum[3]_keep ;
  wire \PWMC/RemaTxNum[4]_keep ;
  wire \PWMC/RemaTxNum[5]_keep ;
  wire \PWMC/RemaTxNum[6]_keep ;
  wire \PWMC/RemaTxNum[7]_keep ;
  wire \PWMC/RemaTxNum[8]_keep ;
  wire \PWMC/RemaTxNum[9]_keep ;
  wire \PWMC/dir_keep ;
  wire \PWMC/mux3_b0_sel_is_3_o ;
  wire \PWMC/n0 ;
  wire \PWMC/n1 ;
  wire \PWMC/n10 ;
  wire \PWMC/n11 ;
  wire \PWMC/n17 ;
  wire \PWMC/n17_neg ;
  wire \PWMC/n18 ;
  wire \PWMC/n24 ;
  wire \PWMC/n25 ;
  wire \PWMC/n25_neg ;
  wire \PWMC/n32 ;
  wire \PWMC/n4 ;
  wire \PWMC/n4_neg ;
  wire \PWMC/n5 ;
  wire \PWMC/n6 ;
  wire \PWMC/n6_neg ;
  wire \PWMC/n8 ;
  wire \PWMC/n9 ;
  wire \PWMC/pnumr[0]_keep ;
  wire \PWMC/pnumr[10]_keep ;
  wire \PWMC/pnumr[11]_keep ;
  wire \PWMC/pnumr[12]_keep ;
  wire \PWMC/pnumr[13]_keep ;
  wire \PWMC/pnumr[14]_keep ;
  wire \PWMC/pnumr[15]_keep ;
  wire \PWMC/pnumr[16]_keep ;
  wire \PWMC/pnumr[17]_keep ;
  wire \PWMC/pnumr[18]_keep ;
  wire \PWMC/pnumr[19]_keep ;
  wire \PWMC/pnumr[1]_keep ;
  wire \PWMC/pnumr[20]_keep ;
  wire \PWMC/pnumr[21]_keep ;
  wire \PWMC/pnumr[22]_keep ;
  wire \PWMC/pnumr[23]_keep ;
  wire \PWMC/pnumr[24]_keep ;
  wire \PWMC/pnumr[25]_keep ;
  wire \PWMC/pnumr[26]_keep ;
  wire \PWMC/pnumr[27]_keep ;
  wire \PWMC/pnumr[28]_keep ;
  wire \PWMC/pnumr[29]_keep ;
  wire \PWMC/pnumr[2]_keep ;
  wire \PWMC/pnumr[30]_keep ;
  wire \PWMC/pnumr[31]_keep ;
  wire \PWMC/pnumr[3]_keep ;
  wire \PWMC/pnumr[4]_keep ;
  wire \PWMC/pnumr[5]_keep ;
  wire \PWMC/pnumr[6]_keep ;
  wire \PWMC/pnumr[7]_keep ;
  wire \PWMC/pnumr[8]_keep ;
  wire \PWMC/pnumr[9]_keep ;
  wire \PWMC/pwm_keep ;
  wire \PWMC/stopreq ;  // src/OnePWM.v(14)
  wire \PWMC/stopreq_keep ;
  wire \PWMC/u14_sel_is_1_o ;
  wire \PWMC/u17_sel_is_1_o ;
  wire \PWMC/u17_sel_is_1_o_neg ;
  wire \PWMC/u18_sel_is_0_o ;
  wire \PWMC/u8_sel_is_0_o ;
  wire \PWMD/RemaTxNum[0]_keep ;
  wire \PWMD/RemaTxNum[10]_keep ;
  wire \PWMD/RemaTxNum[11]_keep ;
  wire \PWMD/RemaTxNum[12]_keep ;
  wire \PWMD/RemaTxNum[13]_keep ;
  wire \PWMD/RemaTxNum[14]_keep ;
  wire \PWMD/RemaTxNum[15]_keep ;
  wire \PWMD/RemaTxNum[16]_keep ;
  wire \PWMD/RemaTxNum[17]_keep ;
  wire \PWMD/RemaTxNum[18]_keep ;
  wire \PWMD/RemaTxNum[19]_keep ;
  wire \PWMD/RemaTxNum[1]_keep ;
  wire \PWMD/RemaTxNum[20]_keep ;
  wire \PWMD/RemaTxNum[21]_keep ;
  wire \PWMD/RemaTxNum[22]_keep ;
  wire \PWMD/RemaTxNum[23]_keep ;
  wire \PWMD/RemaTxNum[2]_keep ;
  wire \PWMD/RemaTxNum[3]_keep ;
  wire \PWMD/RemaTxNum[4]_keep ;
  wire \PWMD/RemaTxNum[5]_keep ;
  wire \PWMD/RemaTxNum[6]_keep ;
  wire \PWMD/RemaTxNum[7]_keep ;
  wire \PWMD/RemaTxNum[8]_keep ;
  wire \PWMD/RemaTxNum[9]_keep ;
  wire \PWMD/dir_keep ;
  wire \PWMD/mux3_b0_sel_is_3_o ;
  wire \PWMD/n0 ;
  wire \PWMD/n1 ;
  wire \PWMD/n10 ;
  wire \PWMD/n11 ;
  wire \PWMD/n17 ;
  wire \PWMD/n17_neg ;
  wire \PWMD/n18 ;
  wire \PWMD/n24 ;
  wire \PWMD/n25 ;
  wire \PWMD/n25_neg ;
  wire \PWMD/n32 ;
  wire \PWMD/n4 ;
  wire \PWMD/n4_neg ;
  wire \PWMD/n5 ;
  wire \PWMD/n6 ;
  wire \PWMD/n6_neg ;
  wire \PWMD/n8 ;
  wire \PWMD/n9 ;
  wire \PWMD/pnumr[0]_keep ;
  wire \PWMD/pnumr[10]_keep ;
  wire \PWMD/pnumr[11]_keep ;
  wire \PWMD/pnumr[12]_keep ;
  wire \PWMD/pnumr[13]_keep ;
  wire \PWMD/pnumr[14]_keep ;
  wire \PWMD/pnumr[15]_keep ;
  wire \PWMD/pnumr[16]_keep ;
  wire \PWMD/pnumr[17]_keep ;
  wire \PWMD/pnumr[18]_keep ;
  wire \PWMD/pnumr[19]_keep ;
  wire \PWMD/pnumr[1]_keep ;
  wire \PWMD/pnumr[20]_keep ;
  wire \PWMD/pnumr[21]_keep ;
  wire \PWMD/pnumr[22]_keep ;
  wire \PWMD/pnumr[23]_keep ;
  wire \PWMD/pnumr[24]_keep ;
  wire \PWMD/pnumr[25]_keep ;
  wire \PWMD/pnumr[26]_keep ;
  wire \PWMD/pnumr[27]_keep ;
  wire \PWMD/pnumr[28]_keep ;
  wire \PWMD/pnumr[29]_keep ;
  wire \PWMD/pnumr[2]_keep ;
  wire \PWMD/pnumr[30]_keep ;
  wire \PWMD/pnumr[31]_keep ;
  wire \PWMD/pnumr[3]_keep ;
  wire \PWMD/pnumr[4]_keep ;
  wire \PWMD/pnumr[5]_keep ;
  wire \PWMD/pnumr[6]_keep ;
  wire \PWMD/pnumr[7]_keep ;
  wire \PWMD/pnumr[8]_keep ;
  wire \PWMD/pnumr[9]_keep ;
  wire \PWMD/pwm_keep ;
  wire \PWMD/stopreq ;  // src/OnePWM.v(14)
  wire \PWMD/stopreq_keep ;
  wire \PWMD/u14_sel_is_1_o ;
  wire \PWMD/u17_sel_is_1_o ;
  wire \PWMD/u17_sel_is_1_o_neg ;
  wire \PWMD/u18_sel_is_0_o ;
  wire \PWMD/u8_sel_is_0_o ;
  wire \PWME/RemaTxNum[0]_keep ;
  wire \PWME/RemaTxNum[10]_keep ;
  wire \PWME/RemaTxNum[11]_keep ;
  wire \PWME/RemaTxNum[12]_keep ;
  wire \PWME/RemaTxNum[13]_keep ;
  wire \PWME/RemaTxNum[14]_keep ;
  wire \PWME/RemaTxNum[15]_keep ;
  wire \PWME/RemaTxNum[16]_keep ;
  wire \PWME/RemaTxNum[17]_keep ;
  wire \PWME/RemaTxNum[18]_keep ;
  wire \PWME/RemaTxNum[19]_keep ;
  wire \PWME/RemaTxNum[1]_keep ;
  wire \PWME/RemaTxNum[20]_keep ;
  wire \PWME/RemaTxNum[21]_keep ;
  wire \PWME/RemaTxNum[22]_keep ;
  wire \PWME/RemaTxNum[23]_keep ;
  wire \PWME/RemaTxNum[2]_keep ;
  wire \PWME/RemaTxNum[3]_keep ;
  wire \PWME/RemaTxNum[4]_keep ;
  wire \PWME/RemaTxNum[5]_keep ;
  wire \PWME/RemaTxNum[6]_keep ;
  wire \PWME/RemaTxNum[7]_keep ;
  wire \PWME/RemaTxNum[8]_keep ;
  wire \PWME/RemaTxNum[9]_keep ;
  wire \PWME/dir_keep ;
  wire \PWME/mux3_b0_sel_is_3_o ;
  wire \PWME/n0 ;
  wire \PWME/n1 ;
  wire \PWME/n10 ;
  wire \PWME/n11 ;
  wire \PWME/n17 ;
  wire \PWME/n17_neg ;
  wire \PWME/n18 ;
  wire \PWME/n24 ;
  wire \PWME/n25 ;
  wire \PWME/n25_neg ;
  wire \PWME/n32 ;
  wire \PWME/n4 ;
  wire \PWME/n4_neg ;
  wire \PWME/n5 ;
  wire \PWME/n6 ;
  wire \PWME/n6_neg ;
  wire \PWME/n8 ;
  wire \PWME/n9 ;
  wire \PWME/pnumr[0]_keep ;
  wire \PWME/pnumr[10]_keep ;
  wire \PWME/pnumr[11]_keep ;
  wire \PWME/pnumr[12]_keep ;
  wire \PWME/pnumr[13]_keep ;
  wire \PWME/pnumr[14]_keep ;
  wire \PWME/pnumr[15]_keep ;
  wire \PWME/pnumr[16]_keep ;
  wire \PWME/pnumr[17]_keep ;
  wire \PWME/pnumr[18]_keep ;
  wire \PWME/pnumr[19]_keep ;
  wire \PWME/pnumr[1]_keep ;
  wire \PWME/pnumr[20]_keep ;
  wire \PWME/pnumr[21]_keep ;
  wire \PWME/pnumr[22]_keep ;
  wire \PWME/pnumr[23]_keep ;
  wire \PWME/pnumr[24]_keep ;
  wire \PWME/pnumr[25]_keep ;
  wire \PWME/pnumr[26]_keep ;
  wire \PWME/pnumr[27]_keep ;
  wire \PWME/pnumr[28]_keep ;
  wire \PWME/pnumr[29]_keep ;
  wire \PWME/pnumr[2]_keep ;
  wire \PWME/pnumr[30]_keep ;
  wire \PWME/pnumr[31]_keep ;
  wire \PWME/pnumr[3]_keep ;
  wire \PWME/pnumr[4]_keep ;
  wire \PWME/pnumr[5]_keep ;
  wire \PWME/pnumr[6]_keep ;
  wire \PWME/pnumr[7]_keep ;
  wire \PWME/pnumr[8]_keep ;
  wire \PWME/pnumr[9]_keep ;
  wire \PWME/pwm_keep ;
  wire \PWME/stopreq ;  // src/OnePWM.v(14)
  wire \PWME/stopreq_keep ;
  wire \PWME/u14_sel_is_1_o ;
  wire \PWME/u17_sel_is_1_o ;
  wire \PWME/u17_sel_is_1_o_neg ;
  wire \PWME/u18_sel_is_0_o ;
  wire \PWME/u8_sel_is_0_o ;
  wire \PWMF/RemaTxNum[0]_keep ;
  wire \PWMF/RemaTxNum[10]_keep ;
  wire \PWMF/RemaTxNum[11]_keep ;
  wire \PWMF/RemaTxNum[12]_keep ;
  wire \PWMF/RemaTxNum[13]_keep ;
  wire \PWMF/RemaTxNum[14]_keep ;
  wire \PWMF/RemaTxNum[15]_keep ;
  wire \PWMF/RemaTxNum[16]_keep ;
  wire \PWMF/RemaTxNum[17]_keep ;
  wire \PWMF/RemaTxNum[18]_keep ;
  wire \PWMF/RemaTxNum[19]_keep ;
  wire \PWMF/RemaTxNum[1]_keep ;
  wire \PWMF/RemaTxNum[20]_keep ;
  wire \PWMF/RemaTxNum[21]_keep ;
  wire \PWMF/RemaTxNum[22]_keep ;
  wire \PWMF/RemaTxNum[23]_keep ;
  wire \PWMF/RemaTxNum[2]_keep ;
  wire \PWMF/RemaTxNum[3]_keep ;
  wire \PWMF/RemaTxNum[4]_keep ;
  wire \PWMF/RemaTxNum[5]_keep ;
  wire \PWMF/RemaTxNum[6]_keep ;
  wire \PWMF/RemaTxNum[7]_keep ;
  wire \PWMF/RemaTxNum[8]_keep ;
  wire \PWMF/RemaTxNum[9]_keep ;
  wire \PWMF/dir_keep ;
  wire \PWMF/mux3_b0_sel_is_3_o ;
  wire \PWMF/n0 ;
  wire \PWMF/n1 ;
  wire \PWMF/n10 ;
  wire \PWMF/n11 ;
  wire \PWMF/n17 ;
  wire \PWMF/n17_neg ;
  wire \PWMF/n18 ;
  wire \PWMF/n24 ;
  wire \PWMF/n25 ;
  wire \PWMF/n25_neg ;
  wire \PWMF/n32 ;
  wire \PWMF/n4 ;
  wire \PWMF/n4_neg ;
  wire \PWMF/n5 ;
  wire \PWMF/n6 ;
  wire \PWMF/n6_neg ;
  wire \PWMF/n8 ;
  wire \PWMF/n9 ;
  wire \PWMF/pnumr[0]_keep ;
  wire \PWMF/pnumr[10]_keep ;
  wire \PWMF/pnumr[11]_keep ;
  wire \PWMF/pnumr[12]_keep ;
  wire \PWMF/pnumr[13]_keep ;
  wire \PWMF/pnumr[14]_keep ;
  wire \PWMF/pnumr[15]_keep ;
  wire \PWMF/pnumr[16]_keep ;
  wire \PWMF/pnumr[17]_keep ;
  wire \PWMF/pnumr[18]_keep ;
  wire \PWMF/pnumr[19]_keep ;
  wire \PWMF/pnumr[1]_keep ;
  wire \PWMF/pnumr[20]_keep ;
  wire \PWMF/pnumr[21]_keep ;
  wire \PWMF/pnumr[22]_keep ;
  wire \PWMF/pnumr[23]_keep ;
  wire \PWMF/pnumr[24]_keep ;
  wire \PWMF/pnumr[25]_keep ;
  wire \PWMF/pnumr[26]_keep ;
  wire \PWMF/pnumr[27]_keep ;
  wire \PWMF/pnumr[28]_keep ;
  wire \PWMF/pnumr[29]_keep ;
  wire \PWMF/pnumr[2]_keep ;
  wire \PWMF/pnumr[30]_keep ;
  wire \PWMF/pnumr[31]_keep ;
  wire \PWMF/pnumr[3]_keep ;
  wire \PWMF/pnumr[4]_keep ;
  wire \PWMF/pnumr[5]_keep ;
  wire \PWMF/pnumr[6]_keep ;
  wire \PWMF/pnumr[7]_keep ;
  wire \PWMF/pnumr[8]_keep ;
  wire \PWMF/pnumr[9]_keep ;
  wire \PWMF/pwm_keep ;
  wire \PWMF/stopreq ;  // src/OnePWM.v(14)
  wire \PWMF/stopreq_keep ;
  wire \PWMF/u14_sel_is_1_o ;
  wire \PWMF/u17_sel_is_1_o ;
  wire \PWMF/u17_sel_is_1_o_neg ;
  wire \PWMF/u18_sel_is_0_o ;
  wire \PWMF/u8_sel_is_0_o ;
  wire \U_AHB/h2h_hwrite ;  // src/AHB.v(22)
  wire \U_AHB/h2h_hwritew ;  // src/AHB.v(19)
  wire \U_AHB/n0 ;
  wire \U_AHB/n1 ;
  wire \U_AHB/n10 ;
  wire \U_AHB/n100 ;
  wire \U_AHB/n101 ;
  wire \U_AHB/n102 ;
  wire \U_AHB/n103 ;
  wire \U_AHB/n104 ;
  wire \U_AHB/n105 ;
  wire \U_AHB/n106 ;
  wire \U_AHB/n107 ;
  wire \U_AHB/n108 ;
  wire \U_AHB/n109 ;
  wire \U_AHB/n110 ;
  wire \U_AHB/n111 ;
  wire \U_AHB/n112 ;
  wire \U_AHB/n113 ;
  wire \U_AHB/n115 ;
  wire \U_AHB/n12 ;
  wire \U_AHB/n14 ;
  wire \U_AHB/n16 ;
  wire \U_AHB/n18 ;
  wire \U_AHB/n2 ;
  wire \U_AHB/n20 ;
  wire \U_AHB/n22 ;
  wire \U_AHB/n24 ;
  wire \U_AHB/n26 ;
  wire \U_AHB/n28 ;
  wire \U_AHB/n30 ;
  wire \U_AHB/n32 ;
  wire \U_AHB/n34 ;
  wire \U_AHB/n36 ;
  wire \U_AHB/n38 ;
  wire \U_AHB/n4 ;
  wire \U_AHB/n43 ;
  wire \U_AHB/n44 ;
  wire \U_AHB/n45 ;
  wire \U_AHB/n47 ;
  wire \U_AHB/n49 ;
  wire \U_AHB/n50 ;
  wire \U_AHB/n51 ;
  wire \U_AHB/n53 ;
  wire \U_AHB/n55 ;
  wire \U_AHB/n57 ;
  wire \U_AHB/n59 ;
  wire \U_AHB/n6 ;
  wire \U_AHB/n61 ;
  wire \U_AHB/n63 ;
  wire \U_AHB/n65 ;
  wire \U_AHB/n67 ;
  wire \U_AHB/n69 ;
  wire \U_AHB/n7 ;
  wire \U_AHB/n71 ;
  wire \U_AHB/n73 ;
  wire \U_AHB/n75 ;
  wire \U_AHB/n77 ;
  wire \U_AHB/n79 ;
  wire \U_AHB/n8 ;
  wire \U_AHB/n81 ;
  wire \U_AHB/n82 ;
  wire \U_AHB/n83 ;
  wire \U_AHB/n84 ;
  wire \U_AHB/n85 ;
  wire \U_AHB/n86 ;
  wire \U_AHB/n87 ;
  wire \U_AHB/n88 ;
  wire \U_AHB/n89 ;
  wire \U_AHB/n90 ;
  wire \U_AHB/n91 ;
  wire \U_AHB/n92 ;
  wire \U_AHB/n93 ;
  wire \U_AHB/n94 ;
  wire \U_AHB/n95 ;
  wire \U_AHB/n96 ;
  wire \U_AHB/n97 ;
  wire \U_AHB/n98 ;
  wire \U_AHB/n99 ;
  wire \U_AHB/sel0_b0/or_B0_or_B1_B2_o_o ;
  wire \U_AHB/sel0_b0/or_B10_B11_o ;
  wire \U_AHB/sel0_b0/or_B1_B2_o ;
  wire \U_AHB/sel0_b0/or_B3_or_B4_B5_o_o ;
  wire \U_AHB/sel0_b0/or_B4_B5_o ;
  wire \U_AHB/sel0_b0/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel0_b0/or_B7_B8_o ;
  wire \U_AHB/sel0_b0/or_B9_or_B10_B11_o_o ;
  wire \U_AHB/sel0_b0/or_or_B0_or_B1_B2_o__o ;
  wire \U_AHB/sel0_b0/or_or_B6_or_B7_B8_o__o ;
  wire \U_AHB/sel0_b1/or_B0_or_B1_B2_o_o ;
  wire \U_AHB/sel0_b1/or_B10_B11_o ;
  wire \U_AHB/sel0_b1/or_B1_B2_o ;
  wire \U_AHB/sel0_b1/or_B3_or_B4_B5_o_o ;
  wire \U_AHB/sel0_b1/or_B4_B5_o ;
  wire \U_AHB/sel0_b1/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel0_b1/or_B7_B8_o ;
  wire \U_AHB/sel0_b1/or_B9_or_B10_B11_o_o ;
  wire \U_AHB/sel0_b1/or_or_B0_or_B1_B2_o__o ;
  wire \U_AHB/sel0_b1/or_or_B6_or_B7_B8_o__o ;
  wire \U_AHB/sel0_b10/or_B0_or_B1_B2_o_o ;
  wire \U_AHB/sel0_b10/or_B10_B11_o ;
  wire \U_AHB/sel0_b10/or_B1_B2_o ;
  wire \U_AHB/sel0_b10/or_B3_or_B4_B5_o_o ;
  wire \U_AHB/sel0_b10/or_B4_B5_o ;
  wire \U_AHB/sel0_b10/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel0_b10/or_B7_B8_o ;
  wire \U_AHB/sel0_b10/or_B9_or_B10_B11_o_o ;
  wire \U_AHB/sel0_b10/or_or_B0_or_B1_B2_o__o ;
  wire \U_AHB/sel0_b10/or_or_B6_or_B7_B8_o__o ;
  wire \U_AHB/sel0_b11/or_B0_or_B1_B2_o_o ;
  wire \U_AHB/sel0_b11/or_B10_B11_o ;
  wire \U_AHB/sel0_b11/or_B1_B2_o ;
  wire \U_AHB/sel0_b11/or_B3_or_B4_B5_o_o ;
  wire \U_AHB/sel0_b11/or_B4_B5_o ;
  wire \U_AHB/sel0_b11/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel0_b11/or_B7_B8_o ;
  wire \U_AHB/sel0_b11/or_B9_or_B10_B11_o_o ;
  wire \U_AHB/sel0_b11/or_or_B0_or_B1_B2_o__o ;
  wire \U_AHB/sel0_b11/or_or_B6_or_B7_B8_o__o ;
  wire \U_AHB/sel0_b12/or_B0_or_B1_B2_o_o ;
  wire \U_AHB/sel0_b12/or_B10_B11_o ;
  wire \U_AHB/sel0_b12/or_B1_B2_o ;
  wire \U_AHB/sel0_b12/or_B3_or_B4_B5_o_o ;
  wire \U_AHB/sel0_b12/or_B4_B5_o ;
  wire \U_AHB/sel0_b12/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel0_b12/or_B7_B8_o ;
  wire \U_AHB/sel0_b12/or_B9_or_B10_B11_o_o ;
  wire \U_AHB/sel0_b12/or_or_B0_or_B1_B2_o__o ;
  wire \U_AHB/sel0_b12/or_or_B6_or_B7_B8_o__o ;
  wire \U_AHB/sel0_b13/or_B0_or_B1_B2_o_o ;
  wire \U_AHB/sel0_b13/or_B10_B11_o ;
  wire \U_AHB/sel0_b13/or_B1_B2_o ;
  wire \U_AHB/sel0_b13/or_B3_or_B4_B5_o_o ;
  wire \U_AHB/sel0_b13/or_B4_B5_o ;
  wire \U_AHB/sel0_b13/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel0_b13/or_B7_B8_o ;
  wire \U_AHB/sel0_b13/or_B9_or_B10_B11_o_o ;
  wire \U_AHB/sel0_b13/or_or_B0_or_B1_B2_o__o ;
  wire \U_AHB/sel0_b13/or_or_B6_or_B7_B8_o__o ;
  wire \U_AHB/sel0_b14/or_B0_or_B1_B2_o_o ;
  wire \U_AHB/sel0_b14/or_B10_B11_o ;
  wire \U_AHB/sel0_b14/or_B1_B2_o ;
  wire \U_AHB/sel0_b14/or_B3_or_B4_B5_o_o ;
  wire \U_AHB/sel0_b14/or_B4_B5_o ;
  wire \U_AHB/sel0_b14/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel0_b14/or_B7_B8_o ;
  wire \U_AHB/sel0_b14/or_B9_or_B10_B11_o_o ;
  wire \U_AHB/sel0_b14/or_or_B0_or_B1_B2_o__o ;
  wire \U_AHB/sel0_b14/or_or_B6_or_B7_B8_o__o ;
  wire \U_AHB/sel0_b15/or_B0_or_B1_B2_o_o ;
  wire \U_AHB/sel0_b15/or_B10_B11_o ;
  wire \U_AHB/sel0_b15/or_B1_B2_o ;
  wire \U_AHB/sel0_b15/or_B3_or_B4_B5_o_o ;
  wire \U_AHB/sel0_b15/or_B4_B5_o ;
  wire \U_AHB/sel0_b15/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel0_b15/or_B7_B8_o ;
  wire \U_AHB/sel0_b15/or_B9_or_B10_B11_o_o ;
  wire \U_AHB/sel0_b15/or_or_B0_or_B1_B2_o__o ;
  wire \U_AHB/sel0_b15/or_or_B6_or_B7_B8_o__o ;
  wire \U_AHB/sel0_b16/or_B0_or_B1_B2_o_o ;
  wire \U_AHB/sel0_b16/or_B10_B11_o ;
  wire \U_AHB/sel0_b16/or_B1_B2_o ;
  wire \U_AHB/sel0_b16/or_B3_or_B4_B5_o_o ;
  wire \U_AHB/sel0_b16/or_B4_B5_o ;
  wire \U_AHB/sel0_b16/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel0_b16/or_B7_B8_o ;
  wire \U_AHB/sel0_b16/or_B9_or_B10_B11_o_o ;
  wire \U_AHB/sel0_b16/or_or_B0_or_B1_B2_o__o ;
  wire \U_AHB/sel0_b16/or_or_B6_or_B7_B8_o__o ;
  wire \U_AHB/sel0_b17/or_B0_or_B1_B2_o_o ;
  wire \U_AHB/sel0_b17/or_B10_B11_o ;
  wire \U_AHB/sel0_b17/or_B1_B2_o ;
  wire \U_AHB/sel0_b17/or_B3_or_B4_B5_o_o ;
  wire \U_AHB/sel0_b17/or_B4_B5_o ;
  wire \U_AHB/sel0_b17/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel0_b17/or_B7_B8_o ;
  wire \U_AHB/sel0_b17/or_B9_or_B10_B11_o_o ;
  wire \U_AHB/sel0_b17/or_or_B0_or_B1_B2_o__o ;
  wire \U_AHB/sel0_b17/or_or_B6_or_B7_B8_o__o ;
  wire \U_AHB/sel0_b18/or_B0_or_B1_B2_o_o ;
  wire \U_AHB/sel0_b18/or_B10_B11_o ;
  wire \U_AHB/sel0_b18/or_B1_B2_o ;
  wire \U_AHB/sel0_b18/or_B3_or_B4_B5_o_o ;
  wire \U_AHB/sel0_b18/or_B4_B5_o ;
  wire \U_AHB/sel0_b18/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel0_b18/or_B7_B8_o ;
  wire \U_AHB/sel0_b18/or_B9_or_B10_B11_o_o ;
  wire \U_AHB/sel0_b18/or_or_B0_or_B1_B2_o__o ;
  wire \U_AHB/sel0_b18/or_or_B6_or_B7_B8_o__o ;
  wire \U_AHB/sel0_b19/or_B0_or_B1_B2_o_o ;
  wire \U_AHB/sel0_b19/or_B10_B11_o ;
  wire \U_AHB/sel0_b19/or_B1_B2_o ;
  wire \U_AHB/sel0_b19/or_B3_or_B4_B5_o_o ;
  wire \U_AHB/sel0_b19/or_B4_B5_o ;
  wire \U_AHB/sel0_b19/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel0_b19/or_B7_B8_o ;
  wire \U_AHB/sel0_b19/or_B9_or_B10_B11_o_o ;
  wire \U_AHB/sel0_b19/or_or_B0_or_B1_B2_o__o ;
  wire \U_AHB/sel0_b19/or_or_B6_or_B7_B8_o__o ;
  wire \U_AHB/sel0_b2/or_B0_or_B1_B2_o_o ;
  wire \U_AHB/sel0_b2/or_B10_B11_o ;
  wire \U_AHB/sel0_b2/or_B1_B2_o ;
  wire \U_AHB/sel0_b2/or_B3_or_B4_B5_o_o ;
  wire \U_AHB/sel0_b2/or_B4_B5_o ;
  wire \U_AHB/sel0_b2/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel0_b2/or_B7_B8_o ;
  wire \U_AHB/sel0_b2/or_B9_or_B10_B11_o_o ;
  wire \U_AHB/sel0_b2/or_or_B0_or_B1_B2_o__o ;
  wire \U_AHB/sel0_b2/or_or_B6_or_B7_B8_o__o ;
  wire \U_AHB/sel0_b20/or_B0_or_B1_B2_o_o ;
  wire \U_AHB/sel0_b20/or_B10_B11_o ;
  wire \U_AHB/sel0_b20/or_B1_B2_o ;
  wire \U_AHB/sel0_b20/or_B3_or_B4_B5_o_o ;
  wire \U_AHB/sel0_b20/or_B4_B5_o ;
  wire \U_AHB/sel0_b20/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel0_b20/or_B7_B8_o ;
  wire \U_AHB/sel0_b20/or_B9_or_B10_B11_o_o ;
  wire \U_AHB/sel0_b20/or_or_B0_or_B1_B2_o__o ;
  wire \U_AHB/sel0_b20/or_or_B6_or_B7_B8_o__o ;
  wire \U_AHB/sel0_b21/or_B0_or_B1_B2_o_o ;
  wire \U_AHB/sel0_b21/or_B10_B11_o ;
  wire \U_AHB/sel0_b21/or_B1_B2_o ;
  wire \U_AHB/sel0_b21/or_B3_or_B4_B5_o_o ;
  wire \U_AHB/sel0_b21/or_B4_B5_o ;
  wire \U_AHB/sel0_b21/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel0_b21/or_B7_B8_o ;
  wire \U_AHB/sel0_b21/or_B9_or_B10_B11_o_o ;
  wire \U_AHB/sel0_b21/or_or_B0_or_B1_B2_o__o ;
  wire \U_AHB/sel0_b21/or_or_B6_or_B7_B8_o__o ;
  wire \U_AHB/sel0_b22/or_B0_or_B1_B2_o_o ;
  wire \U_AHB/sel0_b22/or_B10_B11_o ;
  wire \U_AHB/sel0_b22/or_B1_B2_o ;
  wire \U_AHB/sel0_b22/or_B3_or_B4_B5_o_o ;
  wire \U_AHB/sel0_b22/or_B4_B5_o ;
  wire \U_AHB/sel0_b22/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel0_b22/or_B7_B8_o ;
  wire \U_AHB/sel0_b22/or_B9_or_B10_B11_o_o ;
  wire \U_AHB/sel0_b22/or_or_B0_or_B1_B2_o__o ;
  wire \U_AHB/sel0_b22/or_or_B6_or_B7_B8_o__o ;
  wire \U_AHB/sel0_b23/or_B0_or_B1_B2_o_o ;
  wire \U_AHB/sel0_b23/or_B10_B11_o ;
  wire \U_AHB/sel0_b23/or_B1_B2_o ;
  wire \U_AHB/sel0_b23/or_B3_or_B4_B5_o_o ;
  wire \U_AHB/sel0_b23/or_B4_B5_o ;
  wire \U_AHB/sel0_b23/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel0_b23/or_B7_B8_o ;
  wire \U_AHB/sel0_b23/or_B9_or_B10_B11_o_o ;
  wire \U_AHB/sel0_b23/or_or_B0_or_B1_B2_o__o ;
  wire \U_AHB/sel0_b23/or_or_B6_or_B7_B8_o__o ;
  wire \U_AHB/sel0_b3/or_B0_or_B1_B2_o_o ;
  wire \U_AHB/sel0_b3/or_B10_B11_o ;
  wire \U_AHB/sel0_b3/or_B1_B2_o ;
  wire \U_AHB/sel0_b3/or_B3_or_B4_B5_o_o ;
  wire \U_AHB/sel0_b3/or_B4_B5_o ;
  wire \U_AHB/sel0_b3/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel0_b3/or_B7_B8_o ;
  wire \U_AHB/sel0_b3/or_B9_or_B10_B11_o_o ;
  wire \U_AHB/sel0_b3/or_or_B0_or_B1_B2_o__o ;
  wire \U_AHB/sel0_b3/or_or_B6_or_B7_B8_o__o ;
  wire \U_AHB/sel0_b4/or_B0_or_B1_B2_o_o ;
  wire \U_AHB/sel0_b4/or_B10_B11_o ;
  wire \U_AHB/sel0_b4/or_B1_B2_o ;
  wire \U_AHB/sel0_b4/or_B3_or_B4_B5_o_o ;
  wire \U_AHB/sel0_b4/or_B4_B5_o ;
  wire \U_AHB/sel0_b4/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel0_b4/or_B7_B8_o ;
  wire \U_AHB/sel0_b4/or_B9_or_B10_B11_o_o ;
  wire \U_AHB/sel0_b4/or_or_B0_or_B1_B2_o__o ;
  wire \U_AHB/sel0_b4/or_or_B6_or_B7_B8_o__o ;
  wire \U_AHB/sel0_b5/or_B0_or_B1_B2_o_o ;
  wire \U_AHB/sel0_b5/or_B10_B11_o ;
  wire \U_AHB/sel0_b5/or_B1_B2_o ;
  wire \U_AHB/sel0_b5/or_B3_or_B4_B5_o_o ;
  wire \U_AHB/sel0_b5/or_B4_B5_o ;
  wire \U_AHB/sel0_b5/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel0_b5/or_B7_B8_o ;
  wire \U_AHB/sel0_b5/or_B9_or_B10_B11_o_o ;
  wire \U_AHB/sel0_b5/or_or_B0_or_B1_B2_o__o ;
  wire \U_AHB/sel0_b5/or_or_B6_or_B7_B8_o__o ;
  wire \U_AHB/sel0_b6/or_B0_or_B1_B2_o_o ;
  wire \U_AHB/sel0_b6/or_B10_B11_o ;
  wire \U_AHB/sel0_b6/or_B1_B2_o ;
  wire \U_AHB/sel0_b6/or_B3_or_B4_B5_o_o ;
  wire \U_AHB/sel0_b6/or_B4_B5_o ;
  wire \U_AHB/sel0_b6/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel0_b6/or_B7_B8_o ;
  wire \U_AHB/sel0_b6/or_B9_or_B10_B11_o_o ;
  wire \U_AHB/sel0_b6/or_or_B0_or_B1_B2_o__o ;
  wire \U_AHB/sel0_b6/or_or_B6_or_B7_B8_o__o ;
  wire \U_AHB/sel0_b7/or_B0_or_B1_B2_o_o ;
  wire \U_AHB/sel0_b7/or_B10_B11_o ;
  wire \U_AHB/sel0_b7/or_B1_B2_o ;
  wire \U_AHB/sel0_b7/or_B3_or_B4_B5_o_o ;
  wire \U_AHB/sel0_b7/or_B4_B5_o ;
  wire \U_AHB/sel0_b7/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel0_b7/or_B7_B8_o ;
  wire \U_AHB/sel0_b7/or_B9_or_B10_B11_o_o ;
  wire \U_AHB/sel0_b7/or_or_B0_or_B1_B2_o__o ;
  wire \U_AHB/sel0_b7/or_or_B6_or_B7_B8_o__o ;
  wire \U_AHB/sel0_b8/or_B0_or_B1_B2_o_o ;
  wire \U_AHB/sel0_b8/or_B10_B11_o ;
  wire \U_AHB/sel0_b8/or_B1_B2_o ;
  wire \U_AHB/sel0_b8/or_B3_or_B4_B5_o_o ;
  wire \U_AHB/sel0_b8/or_B4_B5_o ;
  wire \U_AHB/sel0_b8/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel0_b8/or_B7_B8_o ;
  wire \U_AHB/sel0_b8/or_B9_or_B10_B11_o_o ;
  wire \U_AHB/sel0_b8/or_or_B0_or_B1_B2_o__o ;
  wire \U_AHB/sel0_b8/or_or_B6_or_B7_B8_o__o ;
  wire \U_AHB/sel0_b9/or_B0_or_B1_B2_o_o ;
  wire \U_AHB/sel0_b9/or_B10_B11_o ;
  wire \U_AHB/sel0_b9/or_B1_B2_o ;
  wire \U_AHB/sel0_b9/or_B3_or_B4_B5_o_o ;
  wire \U_AHB/sel0_b9/or_B4_B5_o ;
  wire \U_AHB/sel0_b9/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel0_b9/or_B7_B8_o ;
  wire \U_AHB/sel0_b9/or_B9_or_B10_B11_o_o ;
  wire \U_AHB/sel0_b9/or_or_B0_or_B1_B2_o__o ;
  wire \U_AHB/sel0_b9/or_or_B6_or_B7_B8_o__o ;
  wire \U_AHB/sel1_b0/or_B0_B1_o ;
  wire \U_AHB/sel1_b0/or_B4_B5_o ;
  wire \U_AHB/sel1_b0/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel1_b0/or_B7_B8_o ;
  wire \U_AHB/sel1_b0/or_or_B0_B1_o_or_B2__o ;
  wire \U_AHB/sel1_b0/or_or_B4_B5_o_or_B6__o ;
  wire \U_AHB/sel1_b1/or_B0_B1_o ;
  wire \U_AHB/sel1_b1/or_B4_B5_o ;
  wire \U_AHB/sel1_b1/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel1_b1/or_B7_B8_o ;
  wire \U_AHB/sel1_b1/or_or_B0_B1_o_or_B2__o ;
  wire \U_AHB/sel1_b1/or_or_B4_B5_o_or_B6__o ;
  wire \U_AHB/sel1_b10/or_B0_B1_o ;
  wire \U_AHB/sel1_b10/or_B4_B5_o ;
  wire \U_AHB/sel1_b10/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel1_b10/or_B7_B8_o ;
  wire \U_AHB/sel1_b10/or_or_B0_B1_o_or_B2__o ;
  wire \U_AHB/sel1_b10/or_or_B4_B5_o_or_B6__o ;
  wire \U_AHB/sel1_b11/or_B0_B1_o ;
  wire \U_AHB/sel1_b11/or_B4_B5_o ;
  wire \U_AHB/sel1_b11/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel1_b11/or_B7_B8_o ;
  wire \U_AHB/sel1_b11/or_or_B0_B1_o_or_B2__o ;
  wire \U_AHB/sel1_b11/or_or_B4_B5_o_or_B6__o ;
  wire \U_AHB/sel1_b12/or_B0_B1_o ;
  wire \U_AHB/sel1_b12/or_B4_B5_o ;
  wire \U_AHB/sel1_b12/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel1_b12/or_B7_B8_o ;
  wire \U_AHB/sel1_b12/or_or_B0_B1_o_or_B2__o ;
  wire \U_AHB/sel1_b12/or_or_B4_B5_o_or_B6__o ;
  wire \U_AHB/sel1_b13/or_B0_B1_o ;
  wire \U_AHB/sel1_b13/or_B4_B5_o ;
  wire \U_AHB/sel1_b13/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel1_b13/or_B7_B8_o ;
  wire \U_AHB/sel1_b13/or_or_B0_B1_o_or_B2__o ;
  wire \U_AHB/sel1_b13/or_or_B4_B5_o_or_B6__o ;
  wire \U_AHB/sel1_b14/or_B0_B1_o ;
  wire \U_AHB/sel1_b14/or_B4_B5_o ;
  wire \U_AHB/sel1_b14/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel1_b14/or_B7_B8_o ;
  wire \U_AHB/sel1_b14/or_or_B0_B1_o_or_B2__o ;
  wire \U_AHB/sel1_b14/or_or_B4_B5_o_or_B6__o ;
  wire \U_AHB/sel1_b15/or_B0_B1_o ;
  wire \U_AHB/sel1_b15/or_B4_B5_o ;
  wire \U_AHB/sel1_b15/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel1_b15/or_B7_B8_o ;
  wire \U_AHB/sel1_b15/or_or_B0_B1_o_or_B2__o ;
  wire \U_AHB/sel1_b15/or_or_B4_B5_o_or_B6__o ;
  wire \U_AHB/sel1_b16/or_B0_B1_o ;
  wire \U_AHB/sel1_b16/or_B4_B5_o ;
  wire \U_AHB/sel1_b16/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel1_b16/or_B7_B8_o ;
  wire \U_AHB/sel1_b16/or_or_B0_B1_o_or_B2__o ;
  wire \U_AHB/sel1_b16/or_or_B4_B5_o_or_B6__o ;
  wire \U_AHB/sel1_b17/or_B0_B1_o ;
  wire \U_AHB/sel1_b17/or_B4_B5_o ;
  wire \U_AHB/sel1_b17/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel1_b17/or_B7_B8_o ;
  wire \U_AHB/sel1_b17/or_or_B0_B1_o_or_B2__o ;
  wire \U_AHB/sel1_b17/or_or_B4_B5_o_or_B6__o ;
  wire \U_AHB/sel1_b18/or_B0_B1_o ;
  wire \U_AHB/sel1_b18/or_B4_B5_o ;
  wire \U_AHB/sel1_b18/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel1_b18/or_B7_B8_o ;
  wire \U_AHB/sel1_b18/or_or_B0_B1_o_or_B2__o ;
  wire \U_AHB/sel1_b18/or_or_B4_B5_o_or_B6__o ;
  wire \U_AHB/sel1_b19/or_B0_B1_o ;
  wire \U_AHB/sel1_b19/or_B4_B5_o ;
  wire \U_AHB/sel1_b19/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel1_b19/or_B7_B8_o ;
  wire \U_AHB/sel1_b19/or_or_B0_B1_o_or_B2__o ;
  wire \U_AHB/sel1_b19/or_or_B4_B5_o_or_B6__o ;
  wire \U_AHB/sel1_b2/or_B0_B1_o ;
  wire \U_AHB/sel1_b2/or_B4_B5_o ;
  wire \U_AHB/sel1_b2/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel1_b2/or_B7_B8_o ;
  wire \U_AHB/sel1_b2/or_or_B0_B1_o_or_B2__o ;
  wire \U_AHB/sel1_b2/or_or_B4_B5_o_or_B6__o ;
  wire \U_AHB/sel1_b20/or_B0_B1_o ;
  wire \U_AHB/sel1_b20/or_B4_B5_o ;
  wire \U_AHB/sel1_b20/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel1_b20/or_B7_B8_o ;
  wire \U_AHB/sel1_b20/or_or_B0_B1_o_or_B2__o ;
  wire \U_AHB/sel1_b20/or_or_B4_B5_o_or_B6__o ;
  wire \U_AHB/sel1_b21/or_B0_B1_o ;
  wire \U_AHB/sel1_b21/or_B4_B5_o ;
  wire \U_AHB/sel1_b21/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel1_b21/or_B7_B8_o ;
  wire \U_AHB/sel1_b21/or_or_B0_B1_o_or_B2__o ;
  wire \U_AHB/sel1_b21/or_or_B4_B5_o_or_B6__o ;
  wire \U_AHB/sel1_b22/or_B0_B1_o ;
  wire \U_AHB/sel1_b22/or_B4_B5_o ;
  wire \U_AHB/sel1_b22/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel1_b22/or_B7_B8_o ;
  wire \U_AHB/sel1_b22/or_or_B0_B1_o_or_B2__o ;
  wire \U_AHB/sel1_b22/or_or_B4_B5_o_or_B6__o ;
  wire \U_AHB/sel1_b23/or_B0_B1_o ;
  wire \U_AHB/sel1_b23/or_B4_B5_o ;
  wire \U_AHB/sel1_b23/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel1_b23/or_B7_B8_o ;
  wire \U_AHB/sel1_b23/or_or_B0_B1_o_or_B2__o ;
  wire \U_AHB/sel1_b23/or_or_B4_B5_o_or_B6__o ;
  wire \U_AHB/sel1_b24/or_B0_B1_o ;
  wire \U_AHB/sel1_b24/or_or_B0_B1_o_or_B2__o ;
  wire \U_AHB/sel1_b25/or_B0_B1_o ;
  wire \U_AHB/sel1_b25/or_or_B0_B1_o_or_B2__o ;
  wire \U_AHB/sel1_b26/or_B0_B1_o ;
  wire \U_AHB/sel1_b26/or_or_B0_B1_o_or_B2__o ;
  wire \U_AHB/sel1_b27/or_B0_B1_o ;
  wire \U_AHB/sel1_b27/or_or_B0_B1_o_or_B2__o ;
  wire \U_AHB/sel1_b28/or_B0_B1_o ;
  wire \U_AHB/sel1_b28/or_or_B0_B1_o_or_B2__o ;
  wire \U_AHB/sel1_b29/or_B0_B1_o ;
  wire \U_AHB/sel1_b29/or_or_B0_B1_o_or_B2__o ;
  wire \U_AHB/sel1_b3/or_B0_B1_o ;
  wire \U_AHB/sel1_b3/or_B4_B5_o ;
  wire \U_AHB/sel1_b3/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel1_b3/or_B7_B8_o ;
  wire \U_AHB/sel1_b3/or_or_B0_B1_o_or_B2__o ;
  wire \U_AHB/sel1_b3/or_or_B4_B5_o_or_B6__o ;
  wire \U_AHB/sel1_b30/or_B0_B1_o ;
  wire \U_AHB/sel1_b30/or_or_B0_B1_o_or_B2__o ;
  wire \U_AHB/sel1_b31/or_B0_B1_o ;
  wire \U_AHB/sel1_b31/or_or_B0_B1_o_or_B2__o ;
  wire \U_AHB/sel1_b4/or_B0_B1_o ;
  wire \U_AHB/sel1_b4/or_B4_B5_o ;
  wire \U_AHB/sel1_b4/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel1_b4/or_B7_B8_o ;
  wire \U_AHB/sel1_b4/or_or_B0_B1_o_or_B2__o ;
  wire \U_AHB/sel1_b4/or_or_B4_B5_o_or_B6__o ;
  wire \U_AHB/sel1_b5/or_B0_B1_o ;
  wire \U_AHB/sel1_b5/or_B4_B5_o ;
  wire \U_AHB/sel1_b5/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel1_b5/or_B7_B8_o ;
  wire \U_AHB/sel1_b5/or_or_B0_B1_o_or_B2__o ;
  wire \U_AHB/sel1_b5/or_or_B4_B5_o_or_B6__o ;
  wire \U_AHB/sel1_b6/or_B0_B1_o ;
  wire \U_AHB/sel1_b6/or_B4_B5_o ;
  wire \U_AHB/sel1_b6/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel1_b6/or_B7_B8_o ;
  wire \U_AHB/sel1_b6/or_or_B0_B1_o_or_B2__o ;
  wire \U_AHB/sel1_b6/or_or_B4_B5_o_or_B6__o ;
  wire \U_AHB/sel1_b7/or_B0_B1_o ;
  wire \U_AHB/sel1_b7/or_B4_B5_o ;
  wire \U_AHB/sel1_b7/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel1_b7/or_B7_B8_o ;
  wire \U_AHB/sel1_b7/or_or_B0_B1_o_or_B2__o ;
  wire \U_AHB/sel1_b7/or_or_B4_B5_o_or_B6__o ;
  wire \U_AHB/sel1_b8/or_B0_B1_o ;
  wire \U_AHB/sel1_b8/or_B4_B5_o ;
  wire \U_AHB/sel1_b8/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel1_b8/or_B7_B8_o ;
  wire \U_AHB/sel1_b8/or_or_B0_B1_o_or_B2__o ;
  wire \U_AHB/sel1_b8/or_or_B4_B5_o_or_B6__o ;
  wire \U_AHB/sel1_b9/or_B0_B1_o ;
  wire \U_AHB/sel1_b9/or_B4_B5_o ;
  wire \U_AHB/sel1_b9/or_B6_or_B7_B8_o_o ;
  wire \U_AHB/sel1_b9/or_B7_B8_o ;
  wire \U_AHB/sel1_b9/or_or_B0_B1_o_or_B2__o ;
  wire \U_AHB/sel1_b9/or_or_B4_B5_o_or_B6__o ;
  wire clk100m;  // CPLD_SOC_AHB_TOP.v(13)
  wire clk25m;  // CPLD_SOC_AHB_TOP.v(13)
  wire mux2_b0_sel_is_0_o;
  wire mux3_b0_sel_is_2_o;
  wire mux3_b3_sel_is_0_o;
  wire mux4_b2_sel_is_0_o;
  wire mux4_b3_sel_is_2_o;
  wire n1;
  wire n11;
  wire n12;
  wire n13;
  wire n14;
  wire n15;
  wire n16;
  wire n17;
  wire n18;
  wire n19;
  wire n1_neg;
  wire n20;
  wire n21;
  wire n22;
  wire n23;
  wire n24;
  wire n25;
  wire n26;
  wire n4;
  wire n4_neg;
  wire n5;
  wire n5_neg;
  wire n6;
  wire n6_neg;
  wire \pwm_start_stop[16]_neg ;
  wire \pwm_start_stop[17]_neg ;
  wire \pwm_start_stop[18]_neg ;
  wire \pwm_start_stop[19]_neg ;
  wire \pwm_start_stop[20]_neg ;
  wire \pwm_start_stop[21]_neg ;
  wire \pwm_start_stop[22]_neg ;
  wire \pwm_start_stop[23]_neg ;
  wire \pwm_start_stop[24]_neg ;
  wire \pwm_start_stop[25]_neg ;
  wire \pwm_start_stop[26]_neg ;
  wire \pwm_start_stop[27]_neg ;
  wire \pwm_start_stop[28]_neg ;
  wire \pwm_start_stop[29]_neg ;
  wire \pwm_start_stop[30]_neg ;
  wire \pwm_start_stop[31]_neg ;
  wire rstn;  // CPLD_SOC_AHB_TOP.v(13)

  reg_ar_as_w1 \PWM0/State_reg  (
    .clk(clk100m),
    .d(\PWM0/n10 ),
    .en(1'b1),
    .reset(~rstn),
    .set(1'b0),
    .q(pwm_state_read[0]));  // src/OnePWM.v(26)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[0]  (
    .i(\PWM0/RemaTxNum[0]_keep ),
    .o(pnumcnt0[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[10]  (
    .i(\PWM0/RemaTxNum[10]_keep ),
    .o(pnumcnt0[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[11]  (
    .i(\PWM0/RemaTxNum[11]_keep ),
    .o(pnumcnt0[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[12]  (
    .i(\PWM0/RemaTxNum[12]_keep ),
    .o(pnumcnt0[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[13]  (
    .i(\PWM0/RemaTxNum[13]_keep ),
    .o(pnumcnt0[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[14]  (
    .i(\PWM0/RemaTxNum[14]_keep ),
    .o(pnumcnt0[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[15]  (
    .i(\PWM0/RemaTxNum[15]_keep ),
    .o(pnumcnt0[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[16]  (
    .i(\PWM0/RemaTxNum[16]_keep ),
    .o(pnumcnt0[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[17]  (
    .i(\PWM0/RemaTxNum[17]_keep ),
    .o(pnumcnt0[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[18]  (
    .i(\PWM0/RemaTxNum[18]_keep ),
    .o(pnumcnt0[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[19]  (
    .i(\PWM0/RemaTxNum[19]_keep ),
    .o(pnumcnt0[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[1]  (
    .i(\PWM0/RemaTxNum[1]_keep ),
    .o(pnumcnt0[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[20]  (
    .i(\PWM0/RemaTxNum[20]_keep ),
    .o(pnumcnt0[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[21]  (
    .i(\PWM0/RemaTxNum[21]_keep ),
    .o(pnumcnt0[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[22]  (
    .i(\PWM0/RemaTxNum[22]_keep ),
    .o(pnumcnt0[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[23]  (
    .i(\PWM0/RemaTxNum[23]_keep ),
    .o(pnumcnt0[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[2]  (
    .i(\PWM0/RemaTxNum[2]_keep ),
    .o(pnumcnt0[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[3]  (
    .i(\PWM0/RemaTxNum[3]_keep ),
    .o(pnumcnt0[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[4]  (
    .i(\PWM0/RemaTxNum[4]_keep ),
    .o(pnumcnt0[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[5]  (
    .i(\PWM0/RemaTxNum[5]_keep ),
    .o(pnumcnt0[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[6]  (
    .i(\PWM0/RemaTxNum[6]_keep ),
    .o(pnumcnt0[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[7]  (
    .i(\PWM0/RemaTxNum[7]_keep ),
    .o(pnumcnt0[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[8]  (
    .i(\PWM0/RemaTxNum[8]_keep ),
    .o(pnumcnt0[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_RemaTxNum[9]  (
    .i(\PWM0/RemaTxNum[9]_keep ),
    .o(pnumcnt0[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_dir  (
    .i(\PWM0/dir_keep ),
    .o(dir[0]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[0]  (
    .i(\PWM0/pnumr[0]_keep ),
    .o(\PWM0/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[10]  (
    .i(\PWM0/pnumr[10]_keep ),
    .o(\PWM0/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[11]  (
    .i(\PWM0/pnumr[11]_keep ),
    .o(\PWM0/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[12]  (
    .i(\PWM0/pnumr[12]_keep ),
    .o(\PWM0/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[13]  (
    .i(\PWM0/pnumr[13]_keep ),
    .o(\PWM0/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[14]  (
    .i(\PWM0/pnumr[14]_keep ),
    .o(\PWM0/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[15]  (
    .i(\PWM0/pnumr[15]_keep ),
    .o(\PWM0/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[16]  (
    .i(\PWM0/pnumr[16]_keep ),
    .o(\PWM0/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[17]  (
    .i(\PWM0/pnumr[17]_keep ),
    .o(\PWM0/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[18]  (
    .i(\PWM0/pnumr[18]_keep ),
    .o(\PWM0/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[19]  (
    .i(\PWM0/pnumr[19]_keep ),
    .o(\PWM0/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[1]  (
    .i(\PWM0/pnumr[1]_keep ),
    .o(\PWM0/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[20]  (
    .i(\PWM0/pnumr[20]_keep ),
    .o(\PWM0/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[21]  (
    .i(\PWM0/pnumr[21]_keep ),
    .o(\PWM0/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[22]  (
    .i(\PWM0/pnumr[22]_keep ),
    .o(\PWM0/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[23]  (
    .i(\PWM0/pnumr[23]_keep ),
    .o(\PWM0/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[24]  (
    .i(\PWM0/pnumr[24]_keep ),
    .o(\PWM0/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[25]  (
    .i(\PWM0/pnumr[25]_keep ),
    .o(\PWM0/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[26]  (
    .i(\PWM0/pnumr[26]_keep ),
    .o(\PWM0/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[27]  (
    .i(\PWM0/pnumr[27]_keep ),
    .o(\PWM0/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[28]  (
    .i(\PWM0/pnumr[28]_keep ),
    .o(\PWM0/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[29]  (
    .i(\PWM0/pnumr[29]_keep ),
    .o(\PWM0/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[2]  (
    .i(\PWM0/pnumr[2]_keep ),
    .o(\PWM0/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[30]  (
    .i(\PWM0/pnumr[30]_keep ),
    .o(\PWM0/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[31]  (
    .i(\PWM0/pnumr[31]_keep ),
    .o(\PWM0/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[3]  (
    .i(\PWM0/pnumr[3]_keep ),
    .o(\PWM0/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[4]  (
    .i(\PWM0/pnumr[4]_keep ),
    .o(\PWM0/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[5]  (
    .i(\PWM0/pnumr[5]_keep ),
    .o(\PWM0/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[6]  (
    .i(\PWM0/pnumr[6]_keep ),
    .o(\PWM0/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[7]  (
    .i(\PWM0/pnumr[7]_keep ),
    .o(\PWM0/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[8]  (
    .i(\PWM0/pnumr[8]_keep ),
    .o(\PWM0/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pnumr[9]  (
    .i(\PWM0/pnumr[9]_keep ),
    .o(\PWM0/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_pwm  (
    .i(\PWM0/pwm_keep ),
    .o(pwm[0]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM0/_bufkeep_stopreq  (
    .i(\PWM0/stopreq_keep ),
    .o(\PWM0/stopreq ));  // src/OnePWM.v(14)
  reg_ar_as_w1 \PWM0/dir_reg  (
    .clk(clk100m),
    .d(\PWM0/n32 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/dir_keep ));  // src/OnePWM.v(58)
  eq_w27 \PWM0/eq0  (
    .i0(\PWM0/FreCnt ),
    .i1(27'b000000000000000000000000000),
    .o(\PWM0/n0 ));  // src/OnePWM.v(15)
  eq_w24 \PWM0/eq1  (
    .i0(pnumcnt0),
    .i1(24'b000000000000000000000001),
    .o(\PWM0/n5 ));  // src/OnePWM.v(25)
  eq_w27 \PWM0/eq2  (
    .i0(\PWM0/FreCnt ),
    .i1({1'b0,\PWM0/FreCntr [26:1]}),
    .o(\PWM0/n17 ));  // src/OnePWM.v(41)
  eq_w27 \PWM0/eq3  (
    .i0(\PWM0/FreCnt ),
    .i1(\PWM0/FreCntr ),
    .o(\PWM0/n18 ));  // src/OnePWM.v(43)
  binary_mux_s1_w1 \PWM0/mux0_b0  (
    .i0(\PWM0/n12 [0]),
    .i1(freq0[0]),
    .sel(\PWM0/n0 ),
    .o(\PWM0/n13 [0]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM0/mux0_b1  (
    .i0(\PWM0/n12 [1]),
    .i1(freq0[1]),
    .sel(\PWM0/n0 ),
    .o(\PWM0/n13 [1]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM0/mux0_b10  (
    .i0(\PWM0/n12 [10]),
    .i1(freq0[10]),
    .sel(\PWM0/n0 ),
    .o(\PWM0/n13 [10]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM0/mux0_b11  (
    .i0(\PWM0/n12 [11]),
    .i1(freq0[11]),
    .sel(\PWM0/n0 ),
    .o(\PWM0/n13 [11]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM0/mux0_b12  (
    .i0(\PWM0/n12 [12]),
    .i1(freq0[12]),
    .sel(\PWM0/n0 ),
    .o(\PWM0/n13 [12]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM0/mux0_b13  (
    .i0(\PWM0/n12 [13]),
    .i1(freq0[13]),
    .sel(\PWM0/n0 ),
    .o(\PWM0/n13 [13]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM0/mux0_b14  (
    .i0(\PWM0/n12 [14]),
    .i1(freq0[14]),
    .sel(\PWM0/n0 ),
    .o(\PWM0/n13 [14]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM0/mux0_b15  (
    .i0(\PWM0/n12 [15]),
    .i1(freq0[15]),
    .sel(\PWM0/n0 ),
    .o(\PWM0/n13 [15]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM0/mux0_b16  (
    .i0(\PWM0/n12 [16]),
    .i1(freq0[16]),
    .sel(\PWM0/n0 ),
    .o(\PWM0/n13 [16]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM0/mux0_b17  (
    .i0(\PWM0/n12 [17]),
    .i1(freq0[17]),
    .sel(\PWM0/n0 ),
    .o(\PWM0/n13 [17]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM0/mux0_b18  (
    .i0(\PWM0/n12 [18]),
    .i1(freq0[18]),
    .sel(\PWM0/n0 ),
    .o(\PWM0/n13 [18]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM0/mux0_b19  (
    .i0(\PWM0/n12 [19]),
    .i1(freq0[19]),
    .sel(\PWM0/n0 ),
    .o(\PWM0/n13 [19]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM0/mux0_b2  (
    .i0(\PWM0/n12 [2]),
    .i1(freq0[2]),
    .sel(\PWM0/n0 ),
    .o(\PWM0/n13 [2]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM0/mux0_b20  (
    .i0(\PWM0/n12 [20]),
    .i1(freq0[20]),
    .sel(\PWM0/n0 ),
    .o(\PWM0/n13 [20]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM0/mux0_b21  (
    .i0(\PWM0/n12 [21]),
    .i1(freq0[21]),
    .sel(\PWM0/n0 ),
    .o(\PWM0/n13 [21]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM0/mux0_b22  (
    .i0(\PWM0/n12 [22]),
    .i1(freq0[22]),
    .sel(\PWM0/n0 ),
    .o(\PWM0/n13 [22]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM0/mux0_b23  (
    .i0(\PWM0/n12 [23]),
    .i1(freq0[23]),
    .sel(\PWM0/n0 ),
    .o(\PWM0/n13 [23]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM0/mux0_b24  (
    .i0(\PWM0/n12 [24]),
    .i1(freq0[24]),
    .sel(\PWM0/n0 ),
    .o(\PWM0/n13 [24]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM0/mux0_b25  (
    .i0(\PWM0/n12 [25]),
    .i1(freq0[25]),
    .sel(\PWM0/n0 ),
    .o(\PWM0/n13 [25]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM0/mux0_b26  (
    .i0(\PWM0/n12 [26]),
    .i1(freq0[26]),
    .sel(\PWM0/n0 ),
    .o(\PWM0/n13 [26]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM0/mux0_b3  (
    .i0(\PWM0/n12 [3]),
    .i1(freq0[3]),
    .sel(\PWM0/n0 ),
    .o(\PWM0/n13 [3]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM0/mux0_b4  (
    .i0(\PWM0/n12 [4]),
    .i1(freq0[4]),
    .sel(\PWM0/n0 ),
    .o(\PWM0/n13 [4]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM0/mux0_b5  (
    .i0(\PWM0/n12 [5]),
    .i1(freq0[5]),
    .sel(\PWM0/n0 ),
    .o(\PWM0/n13 [5]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM0/mux0_b6  (
    .i0(\PWM0/n12 [6]),
    .i1(freq0[6]),
    .sel(\PWM0/n0 ),
    .o(\PWM0/n13 [6]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM0/mux0_b7  (
    .i0(\PWM0/n12 [7]),
    .i1(freq0[7]),
    .sel(\PWM0/n0 ),
    .o(\PWM0/n13 [7]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM0/mux0_b8  (
    .i0(\PWM0/n12 [8]),
    .i1(freq0[8]),
    .sel(\PWM0/n0 ),
    .o(\PWM0/n13 [8]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM0/mux0_b9  (
    .i0(\PWM0/n12 [9]),
    .i1(freq0[9]),
    .sel(\PWM0/n0 ),
    .o(\PWM0/n13 [9]));  // src/OnePWM.v(32)
  and \PWM0/mux3_b0_sel_is_3  (\PWM0/mux3_b0_sel_is_3_o , \PWM0/n11 , \PWM0/n0 );
  binary_mux_s1_w1 \PWM0/mux4_b0  (
    .i0(\PWM0/pnumr [0]),
    .i1(1'b0),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n22 [0]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux4_b1  (
    .i0(\PWM0/pnumr [1]),
    .i1(1'b0),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n22 [1]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux4_b10  (
    .i0(\PWM0/pnumr [10]),
    .i1(1'b0),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n22 [10]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux4_b11  (
    .i0(\PWM0/pnumr [11]),
    .i1(1'b0),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n22 [11]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux4_b12  (
    .i0(\PWM0/pnumr [12]),
    .i1(1'b0),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n22 [12]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux4_b13  (
    .i0(\PWM0/pnumr [13]),
    .i1(1'b0),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n22 [13]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux4_b14  (
    .i0(\PWM0/pnumr [14]),
    .i1(1'b0),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n22 [14]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux4_b15  (
    .i0(\PWM0/pnumr [15]),
    .i1(1'b0),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n22 [15]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux4_b16  (
    .i0(\PWM0/pnumr [16]),
    .i1(1'b0),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n22 [16]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux4_b17  (
    .i0(\PWM0/pnumr [17]),
    .i1(1'b0),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n22 [17]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux4_b18  (
    .i0(\PWM0/pnumr [18]),
    .i1(1'b0),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n22 [18]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux4_b19  (
    .i0(\PWM0/pnumr [19]),
    .i1(1'b0),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n22 [19]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux4_b2  (
    .i0(\PWM0/pnumr [2]),
    .i1(1'b0),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n22 [2]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux4_b20  (
    .i0(\PWM0/pnumr [20]),
    .i1(1'b0),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n22 [20]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux4_b21  (
    .i0(\PWM0/pnumr [21]),
    .i1(1'b0),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n22 [21]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux4_b22  (
    .i0(\PWM0/pnumr [22]),
    .i1(1'b0),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n22 [22]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux4_b23  (
    .i0(\PWM0/pnumr [23]),
    .i1(1'b0),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n22 [23]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux4_b24  (
    .i0(\PWM0/pnumr [24]),
    .i1(1'b0),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n22 [24]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux4_b25  (
    .i0(\PWM0/pnumr [25]),
    .i1(1'b0),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n22 [25]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux4_b26  (
    .i0(\PWM0/pnumr [26]),
    .i1(1'b0),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n22 [26]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux4_b27  (
    .i0(\PWM0/pnumr [27]),
    .i1(1'b0),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n22 [27]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux4_b28  (
    .i0(\PWM0/pnumr [28]),
    .i1(1'b0),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n22 [28]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux4_b29  (
    .i0(\PWM0/pnumr [29]),
    .i1(1'b0),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n22 [29]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux4_b3  (
    .i0(\PWM0/pnumr [3]),
    .i1(1'b0),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n22 [3]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux4_b30  (
    .i0(\PWM0/pnumr [30]),
    .i1(1'b0),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n22 [30]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux4_b31  (
    .i0(\PWM0/pnumr [31]),
    .i1(1'b0),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n22 [31]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux4_b4  (
    .i0(\PWM0/pnumr [4]),
    .i1(1'b0),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n22 [4]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux4_b5  (
    .i0(\PWM0/pnumr [5]),
    .i1(1'b0),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n22 [5]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux4_b6  (
    .i0(\PWM0/pnumr [6]),
    .i1(1'b0),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n22 [6]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux4_b7  (
    .i0(\PWM0/pnumr [7]),
    .i1(1'b0),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n22 [7]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux4_b8  (
    .i0(\PWM0/pnumr [8]),
    .i1(1'b0),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n22 [8]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux4_b9  (
    .i0(\PWM0/pnumr [9]),
    .i1(1'b0),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n22 [9]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux5_b0  (
    .i0(\PWM0/n22 [0]),
    .i1(pnum0[0]),
    .sel(pnum0[32]),
    .o(\PWM0/n23 [0]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux5_b1  (
    .i0(\PWM0/n22 [1]),
    .i1(pnum0[1]),
    .sel(pnum0[32]),
    .o(\PWM0/n23 [1]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux5_b10  (
    .i0(\PWM0/n22 [10]),
    .i1(pnum0[10]),
    .sel(pnum0[32]),
    .o(\PWM0/n23 [10]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux5_b11  (
    .i0(\PWM0/n22 [11]),
    .i1(pnum0[11]),
    .sel(pnum0[32]),
    .o(\PWM0/n23 [11]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux5_b12  (
    .i0(\PWM0/n22 [12]),
    .i1(pnum0[12]),
    .sel(pnum0[32]),
    .o(\PWM0/n23 [12]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux5_b13  (
    .i0(\PWM0/n22 [13]),
    .i1(pnum0[13]),
    .sel(pnum0[32]),
    .o(\PWM0/n23 [13]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux5_b14  (
    .i0(\PWM0/n22 [14]),
    .i1(pnum0[14]),
    .sel(pnum0[32]),
    .o(\PWM0/n23 [14]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux5_b15  (
    .i0(\PWM0/n22 [15]),
    .i1(pnum0[15]),
    .sel(pnum0[32]),
    .o(\PWM0/n23 [15]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux5_b16  (
    .i0(\PWM0/n22 [16]),
    .i1(pnum0[16]),
    .sel(pnum0[32]),
    .o(\PWM0/n23 [16]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux5_b17  (
    .i0(\PWM0/n22 [17]),
    .i1(pnum0[17]),
    .sel(pnum0[32]),
    .o(\PWM0/n23 [17]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux5_b18  (
    .i0(\PWM0/n22 [18]),
    .i1(pnum0[18]),
    .sel(pnum0[32]),
    .o(\PWM0/n23 [18]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux5_b19  (
    .i0(\PWM0/n22 [19]),
    .i1(pnum0[19]),
    .sel(pnum0[32]),
    .o(\PWM0/n23 [19]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux5_b2  (
    .i0(\PWM0/n22 [2]),
    .i1(pnum0[2]),
    .sel(pnum0[32]),
    .o(\PWM0/n23 [2]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux5_b20  (
    .i0(\PWM0/n22 [20]),
    .i1(pnum0[20]),
    .sel(pnum0[32]),
    .o(\PWM0/n23 [20]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux5_b21  (
    .i0(\PWM0/n22 [21]),
    .i1(pnum0[21]),
    .sel(pnum0[32]),
    .o(\PWM0/n23 [21]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux5_b22  (
    .i0(\PWM0/n22 [22]),
    .i1(pnum0[22]),
    .sel(pnum0[32]),
    .o(\PWM0/n23 [22]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux5_b23  (
    .i0(\PWM0/n22 [23]),
    .i1(pnum0[23]),
    .sel(pnum0[32]),
    .o(\PWM0/n23 [23]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux5_b24  (
    .i0(\PWM0/n22 [24]),
    .i1(pnum0[24]),
    .sel(pnum0[32]),
    .o(\PWM0/n23 [24]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux5_b25  (
    .i0(\PWM0/n22 [25]),
    .i1(pnum0[25]),
    .sel(pnum0[32]),
    .o(\PWM0/n23 [25]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux5_b26  (
    .i0(\PWM0/n22 [26]),
    .i1(pnum0[26]),
    .sel(pnum0[32]),
    .o(\PWM0/n23 [26]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux5_b27  (
    .i0(\PWM0/n22 [27]),
    .i1(pnum0[27]),
    .sel(pnum0[32]),
    .o(\PWM0/n23 [27]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux5_b28  (
    .i0(\PWM0/n22 [28]),
    .i1(pnum0[28]),
    .sel(pnum0[32]),
    .o(\PWM0/n23 [28]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux5_b29  (
    .i0(\PWM0/n22 [29]),
    .i1(pnum0[29]),
    .sel(pnum0[32]),
    .o(\PWM0/n23 [29]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux5_b3  (
    .i0(\PWM0/n22 [3]),
    .i1(pnum0[3]),
    .sel(pnum0[32]),
    .o(\PWM0/n23 [3]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux5_b30  (
    .i0(\PWM0/n22 [30]),
    .i1(pnum0[30]),
    .sel(pnum0[32]),
    .o(\PWM0/n23 [30]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux5_b31  (
    .i0(\PWM0/n22 [31]),
    .i1(pnum0[31]),
    .sel(pnum0[32]),
    .o(\PWM0/n23 [31]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux5_b4  (
    .i0(\PWM0/n22 [4]),
    .i1(pnum0[4]),
    .sel(pnum0[32]),
    .o(\PWM0/n23 [4]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux5_b5  (
    .i0(\PWM0/n22 [5]),
    .i1(pnum0[5]),
    .sel(pnum0[32]),
    .o(\PWM0/n23 [5]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux5_b6  (
    .i0(\PWM0/n22 [6]),
    .i1(pnum0[6]),
    .sel(pnum0[32]),
    .o(\PWM0/n23 [6]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux5_b7  (
    .i0(\PWM0/n22 [7]),
    .i1(pnum0[7]),
    .sel(pnum0[32]),
    .o(\PWM0/n23 [7]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux5_b8  (
    .i0(\PWM0/n22 [8]),
    .i1(pnum0[8]),
    .sel(pnum0[32]),
    .o(\PWM0/n23 [8]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux5_b9  (
    .i0(\PWM0/n22 [9]),
    .i1(pnum0[9]),
    .sel(pnum0[32]),
    .o(\PWM0/n23 [9]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM0/mux6_b0  (
    .i0(\PWM0/pnumr [0]),
    .i1(\PWM0/n26 [0]),
    .sel(\PWM0/n25 ),
    .o(\PWM0/n27 [0]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM0/mux6_b1  (
    .i0(\PWM0/pnumr [1]),
    .i1(\PWM0/n26 [1]),
    .sel(\PWM0/n25 ),
    .o(\PWM0/n27 [1]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM0/mux6_b10  (
    .i0(\PWM0/pnumr [10]),
    .i1(\PWM0/n26 [10]),
    .sel(\PWM0/n25 ),
    .o(\PWM0/n27 [10]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM0/mux6_b11  (
    .i0(\PWM0/pnumr [11]),
    .i1(\PWM0/n26 [11]),
    .sel(\PWM0/n25 ),
    .o(\PWM0/n27 [11]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM0/mux6_b12  (
    .i0(\PWM0/pnumr [12]),
    .i1(\PWM0/n26 [12]),
    .sel(\PWM0/n25 ),
    .o(\PWM0/n27 [12]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM0/mux6_b13  (
    .i0(\PWM0/pnumr [13]),
    .i1(\PWM0/n26 [13]),
    .sel(\PWM0/n25 ),
    .o(\PWM0/n27 [13]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM0/mux6_b14  (
    .i0(\PWM0/pnumr [14]),
    .i1(\PWM0/n26 [14]),
    .sel(\PWM0/n25 ),
    .o(\PWM0/n27 [14]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM0/mux6_b15  (
    .i0(\PWM0/pnumr [15]),
    .i1(\PWM0/n26 [15]),
    .sel(\PWM0/n25 ),
    .o(\PWM0/n27 [15]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM0/mux6_b16  (
    .i0(\PWM0/pnumr [16]),
    .i1(\PWM0/n26 [16]),
    .sel(\PWM0/n25 ),
    .o(\PWM0/n27 [16]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM0/mux6_b17  (
    .i0(\PWM0/pnumr [17]),
    .i1(\PWM0/n26 [17]),
    .sel(\PWM0/n25 ),
    .o(\PWM0/n27 [17]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM0/mux6_b18  (
    .i0(\PWM0/pnumr [18]),
    .i1(\PWM0/n26 [18]),
    .sel(\PWM0/n25 ),
    .o(\PWM0/n27 [18]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM0/mux6_b19  (
    .i0(\PWM0/pnumr [19]),
    .i1(\PWM0/n26 [19]),
    .sel(\PWM0/n25 ),
    .o(\PWM0/n27 [19]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM0/mux6_b2  (
    .i0(\PWM0/pnumr [2]),
    .i1(\PWM0/n26 [2]),
    .sel(\PWM0/n25 ),
    .o(\PWM0/n27 [2]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM0/mux6_b20  (
    .i0(\PWM0/pnumr [20]),
    .i1(\PWM0/n26 [20]),
    .sel(\PWM0/n25 ),
    .o(\PWM0/n27 [20]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM0/mux6_b21  (
    .i0(\PWM0/pnumr [21]),
    .i1(\PWM0/n26 [21]),
    .sel(\PWM0/n25 ),
    .o(\PWM0/n27 [21]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM0/mux6_b22  (
    .i0(\PWM0/pnumr [22]),
    .i1(\PWM0/n26 [22]),
    .sel(\PWM0/n25 ),
    .o(\PWM0/n27 [22]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM0/mux6_b23  (
    .i0(\PWM0/pnumr [23]),
    .i1(\PWM0/n26 [23]),
    .sel(\PWM0/n25 ),
    .o(\PWM0/n27 [23]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM0/mux6_b3  (
    .i0(\PWM0/pnumr [3]),
    .i1(\PWM0/n26 [3]),
    .sel(\PWM0/n25 ),
    .o(\PWM0/n27 [3]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM0/mux6_b4  (
    .i0(\PWM0/pnumr [4]),
    .i1(\PWM0/n26 [4]),
    .sel(\PWM0/n25 ),
    .o(\PWM0/n27 [4]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM0/mux6_b5  (
    .i0(\PWM0/pnumr [5]),
    .i1(\PWM0/n26 [5]),
    .sel(\PWM0/n25 ),
    .o(\PWM0/n27 [5]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM0/mux6_b6  (
    .i0(\PWM0/pnumr [6]),
    .i1(\PWM0/n26 [6]),
    .sel(\PWM0/n25 ),
    .o(\PWM0/n27 [6]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM0/mux6_b7  (
    .i0(\PWM0/pnumr [7]),
    .i1(\PWM0/n26 [7]),
    .sel(\PWM0/n25 ),
    .o(\PWM0/n27 [7]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM0/mux6_b8  (
    .i0(\PWM0/pnumr [8]),
    .i1(\PWM0/n26 [8]),
    .sel(\PWM0/n25 ),
    .o(\PWM0/n27 [8]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM0/mux6_b9  (
    .i0(\PWM0/pnumr [9]),
    .i1(\PWM0/n26 [9]),
    .sel(\PWM0/n25 ),
    .o(\PWM0/n27 [9]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM0/mux7_b0  (
    .i0(pnumcnt0[0]),
    .i1(\PWM0/n27 [0]),
    .sel(\PWM0/n24 ),
    .o(\PWM0/n29 [0]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux7_b1  (
    .i0(pnumcnt0[1]),
    .i1(\PWM0/n27 [1]),
    .sel(\PWM0/n24 ),
    .o(\PWM0/n29 [1]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux7_b10  (
    .i0(pnumcnt0[10]),
    .i1(\PWM0/n27 [10]),
    .sel(\PWM0/n24 ),
    .o(\PWM0/n29 [10]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux7_b11  (
    .i0(pnumcnt0[11]),
    .i1(\PWM0/n27 [11]),
    .sel(\PWM0/n24 ),
    .o(\PWM0/n29 [11]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux7_b12  (
    .i0(pnumcnt0[12]),
    .i1(\PWM0/n27 [12]),
    .sel(\PWM0/n24 ),
    .o(\PWM0/n29 [12]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux7_b13  (
    .i0(pnumcnt0[13]),
    .i1(\PWM0/n27 [13]),
    .sel(\PWM0/n24 ),
    .o(\PWM0/n29 [13]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux7_b14  (
    .i0(pnumcnt0[14]),
    .i1(\PWM0/n27 [14]),
    .sel(\PWM0/n24 ),
    .o(\PWM0/n29 [14]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux7_b15  (
    .i0(pnumcnt0[15]),
    .i1(\PWM0/n27 [15]),
    .sel(\PWM0/n24 ),
    .o(\PWM0/n29 [15]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux7_b16  (
    .i0(pnumcnt0[16]),
    .i1(\PWM0/n27 [16]),
    .sel(\PWM0/n24 ),
    .o(\PWM0/n29 [16]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux7_b17  (
    .i0(pnumcnt0[17]),
    .i1(\PWM0/n27 [17]),
    .sel(\PWM0/n24 ),
    .o(\PWM0/n29 [17]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux7_b18  (
    .i0(pnumcnt0[18]),
    .i1(\PWM0/n27 [18]),
    .sel(\PWM0/n24 ),
    .o(\PWM0/n29 [18]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux7_b19  (
    .i0(pnumcnt0[19]),
    .i1(\PWM0/n27 [19]),
    .sel(\PWM0/n24 ),
    .o(\PWM0/n29 [19]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux7_b2  (
    .i0(pnumcnt0[2]),
    .i1(\PWM0/n27 [2]),
    .sel(\PWM0/n24 ),
    .o(\PWM0/n29 [2]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux7_b20  (
    .i0(pnumcnt0[20]),
    .i1(\PWM0/n27 [20]),
    .sel(\PWM0/n24 ),
    .o(\PWM0/n29 [20]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux7_b21  (
    .i0(pnumcnt0[21]),
    .i1(\PWM0/n27 [21]),
    .sel(\PWM0/n24 ),
    .o(\PWM0/n29 [21]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux7_b22  (
    .i0(pnumcnt0[22]),
    .i1(\PWM0/n27 [22]),
    .sel(\PWM0/n24 ),
    .o(\PWM0/n29 [22]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux7_b23  (
    .i0(pnumcnt0[23]),
    .i1(\PWM0/n27 [23]),
    .sel(\PWM0/n24 ),
    .o(\PWM0/n29 [23]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux7_b3  (
    .i0(pnumcnt0[3]),
    .i1(\PWM0/n27 [3]),
    .sel(\PWM0/n24 ),
    .o(\PWM0/n29 [3]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux7_b4  (
    .i0(pnumcnt0[4]),
    .i1(\PWM0/n27 [4]),
    .sel(\PWM0/n24 ),
    .o(\PWM0/n29 [4]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux7_b5  (
    .i0(pnumcnt0[5]),
    .i1(\PWM0/n27 [5]),
    .sel(\PWM0/n24 ),
    .o(\PWM0/n29 [5]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux7_b6  (
    .i0(pnumcnt0[6]),
    .i1(\PWM0/n27 [6]),
    .sel(\PWM0/n24 ),
    .o(\PWM0/n29 [6]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux7_b7  (
    .i0(pnumcnt0[7]),
    .i1(\PWM0/n27 [7]),
    .sel(\PWM0/n24 ),
    .o(\PWM0/n29 [7]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux7_b8  (
    .i0(pnumcnt0[8]),
    .i1(\PWM0/n27 [8]),
    .sel(\PWM0/n24 ),
    .o(\PWM0/n29 [8]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux7_b9  (
    .i0(pnumcnt0[9]),
    .i1(\PWM0/n27 [9]),
    .sel(\PWM0/n24 ),
    .o(\PWM0/n29 [9]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux8_b0  (
    .i0(\PWM0/n29 [0]),
    .i1(\PWM0/pnumr [0]),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n31 [0]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux8_b1  (
    .i0(\PWM0/n29 [1]),
    .i1(\PWM0/pnumr [1]),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n31 [1]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux8_b10  (
    .i0(\PWM0/n29 [10]),
    .i1(\PWM0/pnumr [10]),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n31 [10]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux8_b11  (
    .i0(\PWM0/n29 [11]),
    .i1(\PWM0/pnumr [11]),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n31 [11]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux8_b12  (
    .i0(\PWM0/n29 [12]),
    .i1(\PWM0/pnumr [12]),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n31 [12]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux8_b13  (
    .i0(\PWM0/n29 [13]),
    .i1(\PWM0/pnumr [13]),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n31 [13]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux8_b14  (
    .i0(\PWM0/n29 [14]),
    .i1(\PWM0/pnumr [14]),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n31 [14]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux8_b15  (
    .i0(\PWM0/n29 [15]),
    .i1(\PWM0/pnumr [15]),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n31 [15]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux8_b16  (
    .i0(\PWM0/n29 [16]),
    .i1(\PWM0/pnumr [16]),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n31 [16]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux8_b17  (
    .i0(\PWM0/n29 [17]),
    .i1(\PWM0/pnumr [17]),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n31 [17]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux8_b18  (
    .i0(\PWM0/n29 [18]),
    .i1(\PWM0/pnumr [18]),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n31 [18]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux8_b19  (
    .i0(\PWM0/n29 [19]),
    .i1(\PWM0/pnumr [19]),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n31 [19]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux8_b2  (
    .i0(\PWM0/n29 [2]),
    .i1(\PWM0/pnumr [2]),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n31 [2]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux8_b20  (
    .i0(\PWM0/n29 [20]),
    .i1(\PWM0/pnumr [20]),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n31 [20]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux8_b21  (
    .i0(\PWM0/n29 [21]),
    .i1(\PWM0/pnumr [21]),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n31 [21]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux8_b22  (
    .i0(\PWM0/n29 [22]),
    .i1(\PWM0/pnumr [22]),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n31 [22]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux8_b23  (
    .i0(\PWM0/n29 [23]),
    .i1(\PWM0/pnumr [23]),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n31 [23]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux8_b3  (
    .i0(\PWM0/n29 [3]),
    .i1(\PWM0/pnumr [3]),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n31 [3]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux8_b4  (
    .i0(\PWM0/n29 [4]),
    .i1(\PWM0/pnumr [4]),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n31 [4]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux8_b5  (
    .i0(\PWM0/n29 [5]),
    .i1(\PWM0/pnumr [5]),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n31 [5]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux8_b6  (
    .i0(\PWM0/n29 [6]),
    .i1(\PWM0/pnumr [6]),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n31 [6]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux8_b7  (
    .i0(\PWM0/n29 [7]),
    .i1(\PWM0/pnumr [7]),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n31 [7]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux8_b8  (
    .i0(\PWM0/n29 [8]),
    .i1(\PWM0/pnumr [8]),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n31 [8]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM0/mux8_b9  (
    .i0(\PWM0/n29 [9]),
    .i1(\PWM0/pnumr [9]),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n31 [9]));  // src/OnePWM.v(57)
  not \PWM0/n17_inv  (\PWM0/n17_neg , \PWM0/n17 );
  not \PWM0/n25_inv  (\PWM0/n25_neg , \PWM0/n25 );
  not \PWM0/n4_inv  (\PWM0/n4_neg , \PWM0/n4 );
  not \PWM0/n6_inv  (\PWM0/n6_neg , \PWM0/n6 );
  ne_w24 \PWM0/neq0  (
    .i0(pnumcnt0),
    .i1(24'b000000000000000000000000),
    .o(\PWM0/n25 ));  // src/OnePWM.v(55)
  reg_sr_ss_w1 \PWM0/pwm_reg  (
    .clk(clk100m),
    .d(pwm[0]),
    .en(1'b1),
    .reset(~\PWM0/u14_sel_is_1_o ),
    .set(\PWM0/n18 ),
    .q(\PWM0/pwm_keep ));  // src/OnePWM.v(45)
  reg_sr_as_w1 \PWM0/reg0_b0  (
    .clk(clk100m),
    .d(\PWM0/n13 [0]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [0]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b1  (
    .clk(clk100m),
    .d(\PWM0/n13 [1]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [1]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b10  (
    .clk(clk100m),
    .d(\PWM0/n13 [10]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [10]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b11  (
    .clk(clk100m),
    .d(\PWM0/n13 [11]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [11]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b12  (
    .clk(clk100m),
    .d(\PWM0/n13 [12]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [12]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b13  (
    .clk(clk100m),
    .d(\PWM0/n13 [13]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [13]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b14  (
    .clk(clk100m),
    .d(\PWM0/n13 [14]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [14]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b15  (
    .clk(clk100m),
    .d(\PWM0/n13 [15]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [15]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b16  (
    .clk(clk100m),
    .d(\PWM0/n13 [16]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [16]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b17  (
    .clk(clk100m),
    .d(\PWM0/n13 [17]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [17]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b18  (
    .clk(clk100m),
    .d(\PWM0/n13 [18]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [18]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b19  (
    .clk(clk100m),
    .d(\PWM0/n13 [19]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [19]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b2  (
    .clk(clk100m),
    .d(\PWM0/n13 [2]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [2]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b20  (
    .clk(clk100m),
    .d(\PWM0/n13 [20]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [20]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b21  (
    .clk(clk100m),
    .d(\PWM0/n13 [21]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [21]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b22  (
    .clk(clk100m),
    .d(\PWM0/n13 [22]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [22]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b23  (
    .clk(clk100m),
    .d(\PWM0/n13 [23]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [23]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b24  (
    .clk(clk100m),
    .d(\PWM0/n13 [24]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [24]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b25  (
    .clk(clk100m),
    .d(\PWM0/n13 [25]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [25]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b26  (
    .clk(clk100m),
    .d(\PWM0/n13 [26]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [26]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b3  (
    .clk(clk100m),
    .d(\PWM0/n13 [3]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [3]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b4  (
    .clk(clk100m),
    .d(\PWM0/n13 [4]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [4]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b5  (
    .clk(clk100m),
    .d(\PWM0/n13 [5]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [5]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b6  (
    .clk(clk100m),
    .d(\PWM0/n13 [6]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [6]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b7  (
    .clk(clk100m),
    .d(\PWM0/n13 [7]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [7]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b8  (
    .clk(clk100m),
    .d(\PWM0/n13 [8]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [8]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM0/reg0_b9  (
    .clk(clk100m),
    .d(\PWM0/n13 [9]),
    .en(1'b1),
    .reset(~\PWM0/n11 ),
    .set(1'b0),
    .q(\PWM0/FreCnt [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b0  (
    .clk(clk100m),
    .d(freq0[0]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [0]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b1  (
    .clk(clk100m),
    .d(freq0[1]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [1]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b10  (
    .clk(clk100m),
    .d(freq0[10]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [10]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b11  (
    .clk(clk100m),
    .d(freq0[11]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [11]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b12  (
    .clk(clk100m),
    .d(freq0[12]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [12]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b13  (
    .clk(clk100m),
    .d(freq0[13]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [13]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b14  (
    .clk(clk100m),
    .d(freq0[14]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [14]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b15  (
    .clk(clk100m),
    .d(freq0[15]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [15]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b16  (
    .clk(clk100m),
    .d(freq0[16]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [16]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b17  (
    .clk(clk100m),
    .d(freq0[17]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [17]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b18  (
    .clk(clk100m),
    .d(freq0[18]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [18]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b19  (
    .clk(clk100m),
    .d(freq0[19]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [19]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b2  (
    .clk(clk100m),
    .d(freq0[2]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [2]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b20  (
    .clk(clk100m),
    .d(freq0[20]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [20]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b21  (
    .clk(clk100m),
    .d(freq0[21]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [21]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b22  (
    .clk(clk100m),
    .d(freq0[22]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [22]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b23  (
    .clk(clk100m),
    .d(freq0[23]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [23]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b24  (
    .clk(clk100m),
    .d(freq0[24]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [24]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b25  (
    .clk(clk100m),
    .d(freq0[25]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [25]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b26  (
    .clk(clk100m),
    .d(freq0[26]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [26]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b3  (
    .clk(clk100m),
    .d(freq0[3]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [3]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b4  (
    .clk(clk100m),
    .d(freq0[4]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [4]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b5  (
    .clk(clk100m),
    .d(freq0[5]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [5]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b6  (
    .clk(clk100m),
    .d(freq0[6]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [6]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b7  (
    .clk(clk100m),
    .d(freq0[7]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [7]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b8  (
    .clk(clk100m),
    .d(freq0[8]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [8]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg1_b9  (
    .clk(clk100m),
    .d(freq0[9]),
    .en(\PWM0/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/FreCntr [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM0/reg2_b0  (
    .clk(clk100m),
    .d(\PWM0/n23 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[0]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b1  (
    .clk(clk100m),
    .d(\PWM0/n23 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[1]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b10  (
    .clk(clk100m),
    .d(\PWM0/n23 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[10]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b11  (
    .clk(clk100m),
    .d(\PWM0/n23 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[11]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b12  (
    .clk(clk100m),
    .d(\PWM0/n23 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[12]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b13  (
    .clk(clk100m),
    .d(\PWM0/n23 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[13]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b14  (
    .clk(clk100m),
    .d(\PWM0/n23 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[14]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b15  (
    .clk(clk100m),
    .d(\PWM0/n23 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[15]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b16  (
    .clk(clk100m),
    .d(\PWM0/n23 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[16]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b17  (
    .clk(clk100m),
    .d(\PWM0/n23 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[17]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b18  (
    .clk(clk100m),
    .d(\PWM0/n23 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[18]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b19  (
    .clk(clk100m),
    .d(\PWM0/n23 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[19]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b2  (
    .clk(clk100m),
    .d(\PWM0/n23 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[2]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b20  (
    .clk(clk100m),
    .d(\PWM0/n23 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[20]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b21  (
    .clk(clk100m),
    .d(\PWM0/n23 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[21]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b22  (
    .clk(clk100m),
    .d(\PWM0/n23 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[22]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b23  (
    .clk(clk100m),
    .d(\PWM0/n23 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[23]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b24  (
    .clk(clk100m),
    .d(\PWM0/n23 [24]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[24]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b25  (
    .clk(clk100m),
    .d(\PWM0/n23 [25]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[25]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b26  (
    .clk(clk100m),
    .d(\PWM0/n23 [26]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[26]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b27  (
    .clk(clk100m),
    .d(\PWM0/n23 [27]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[27]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b28  (
    .clk(clk100m),
    .d(\PWM0/n23 [28]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[28]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b29  (
    .clk(clk100m),
    .d(\PWM0/n23 [29]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[29]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b3  (
    .clk(clk100m),
    .d(\PWM0/n23 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[3]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b30  (
    .clk(clk100m),
    .d(\PWM0/n23 [30]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[30]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b31  (
    .clk(clk100m),
    .d(\PWM0/n23 [31]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[31]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b4  (
    .clk(clk100m),
    .d(\PWM0/n23 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[4]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b5  (
    .clk(clk100m),
    .d(\PWM0/n23 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[5]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b6  (
    .clk(clk100m),
    .d(\PWM0/n23 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[6]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b7  (
    .clk(clk100m),
    .d(\PWM0/n23 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[7]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b8  (
    .clk(clk100m),
    .d(\PWM0/n23 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[8]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg2_b9  (
    .clk(clk100m),
    .d(\PWM0/n23 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/pnumr[9]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM0/reg3_b0  (
    .clk(clk100m),
    .d(\PWM0/n31 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[0]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b1  (
    .clk(clk100m),
    .d(\PWM0/n31 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[1]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b10  (
    .clk(clk100m),
    .d(\PWM0/n31 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[10]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b11  (
    .clk(clk100m),
    .d(\PWM0/n31 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[11]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b12  (
    .clk(clk100m),
    .d(\PWM0/n31 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[12]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b13  (
    .clk(clk100m),
    .d(\PWM0/n31 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[13]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b14  (
    .clk(clk100m),
    .d(\PWM0/n31 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[14]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b15  (
    .clk(clk100m),
    .d(\PWM0/n31 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[15]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b16  (
    .clk(clk100m),
    .d(\PWM0/n31 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[16]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b17  (
    .clk(clk100m),
    .d(\PWM0/n31 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[17]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b18  (
    .clk(clk100m),
    .d(\PWM0/n31 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[18]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b19  (
    .clk(clk100m),
    .d(\PWM0/n31 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[19]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b2  (
    .clk(clk100m),
    .d(\PWM0/n31 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[2]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b20  (
    .clk(clk100m),
    .d(\PWM0/n31 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[20]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b21  (
    .clk(clk100m),
    .d(\PWM0/n31 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[21]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b22  (
    .clk(clk100m),
    .d(\PWM0/n31 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[22]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b23  (
    .clk(clk100m),
    .d(\PWM0/n31 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[23]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b3  (
    .clk(clk100m),
    .d(\PWM0/n31 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[3]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b4  (
    .clk(clk100m),
    .d(\PWM0/n31 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[4]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b5  (
    .clk(clk100m),
    .d(\PWM0/n31 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[5]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b6  (
    .clk(clk100m),
    .d(\PWM0/n31 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[6]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b7  (
    .clk(clk100m),
    .d(\PWM0/n31 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[7]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b8  (
    .clk(clk100m),
    .d(\PWM0/n31 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[8]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM0/reg3_b9  (
    .clk(clk100m),
    .d(\PWM0/n31 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM0/RemaTxNum[9]_keep ));  // src/OnePWM.v(58)
  reg_ar_ss_w1 \PWM0/stopreq_reg  (
    .clk(clk100m),
    .d(\PWM0/n1 ),
    .en(1'b1),
    .reset(1'b0),
    .set(pwm_start_stop[0]),
    .q(\PWM0/stopreq_keep ));  // src/OnePWM.v(15)
  add_pu27_mu27_o27 \PWM0/sub0  (
    .i0(\PWM0/FreCnt ),
    .i1(27'b000000000000000000000000001),
    .o(\PWM0/n12 [26:0]));  // src/OnePWM.v(32)
  add_pu24_mu24_o24 \PWM0/sub1  (
    .i0(pnumcnt0),
    .i1(24'b000000000000000000000001),
    .o(\PWM0/n26 [23:0]));  // src/OnePWM.v(55)
  AL_MUX \PWM0/u10  (
    .i0(1'b0),
    .i1(\PWM0/n9 ),
    .sel(n11),
    .o(\PWM0/n10 ));  // src/OnePWM.v(26)
  or \PWM0/u11  (\PWM0/n11 , pwm_state_read[0], pwm_start_stop[16]);  // src/OnePWM.v(30)
  and \PWM0/u14_sel_is_1  (\PWM0/u14_sel_is_1_o , pwm_state_read[0], \PWM0/n17_neg );
  and \PWM0/u15  (\PWM0/n24 , \PWM0/n0 , pwm_state_read[0]);  // src/OnePWM.v(54)
  and \PWM0/u17_sel_is_1  (\PWM0/u17_sel_is_1_o , \PWM0/n24 , \PWM0/n25_neg );
  not \PWM0/u17_sel_is_1_o_inv  (\PWM0/u17_sel_is_1_o_neg , \PWM0/u17_sel_is_1_o );
  AL_MUX \PWM0/u18  (
    .i0(\PWM0/pnumr [31]),
    .i1(dir[0]),
    .sel(\PWM0/u18_sel_is_0_o ),
    .o(\PWM0/n32 ));
  and \PWM0/u18_sel_is_0  (\PWM0/u18_sel_is_0_o , \pwm_start_stop[16]_neg , \PWM0/u17_sel_is_1_o_neg );
  AL_MUX \PWM0/u2  (
    .i0(\PWM0/stopreq ),
    .i1(1'b0),
    .sel(\PWM0/n0 ),
    .o(\PWM0/n1 ));  // src/OnePWM.v(15)
  and \PWM0/u5  (\PWM0/n4 , \PWM0/stopreq , \PWM0/n0 );  // src/OnePWM.v(23)
  and \PWM0/u6  (\PWM0/n6 , \PWM0/n5 , \PWM0/n0 );  // src/OnePWM.v(25)
  AL_MUX \PWM0/u8  (
    .i0(1'b0),
    .i1(pwm_state_read[0]),
    .sel(\PWM0/u8_sel_is_0_o ),
    .o(\PWM0/n8 ));
  and \PWM0/u8_sel_is_0  (\PWM0/u8_sel_is_0_o , \PWM0/n4_neg , \PWM0/n6_neg );
  AL_MUX \PWM0/u9  (
    .i0(\PWM0/n8 ),
    .i1(1'b1),
    .sel(pwm_start_stop[16]),
    .o(\PWM0/n9 ));  // src/OnePWM.v(26)
  reg_ar_as_w1 \PWM1/State_reg  (
    .clk(clk100m),
    .d(\PWM1/n10 ),
    .en(1'b1),
    .reset(~rstn),
    .set(1'b0),
    .q(pwm_state_read[1]));  // src/OnePWM.v(26)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[0]  (
    .i(\PWM1/RemaTxNum[0]_keep ),
    .o(pnumcnt1[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[10]  (
    .i(\PWM1/RemaTxNum[10]_keep ),
    .o(pnumcnt1[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[11]  (
    .i(\PWM1/RemaTxNum[11]_keep ),
    .o(pnumcnt1[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[12]  (
    .i(\PWM1/RemaTxNum[12]_keep ),
    .o(pnumcnt1[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[13]  (
    .i(\PWM1/RemaTxNum[13]_keep ),
    .o(pnumcnt1[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[14]  (
    .i(\PWM1/RemaTxNum[14]_keep ),
    .o(pnumcnt1[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[15]  (
    .i(\PWM1/RemaTxNum[15]_keep ),
    .o(pnumcnt1[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[16]  (
    .i(\PWM1/RemaTxNum[16]_keep ),
    .o(pnumcnt1[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[17]  (
    .i(\PWM1/RemaTxNum[17]_keep ),
    .o(pnumcnt1[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[18]  (
    .i(\PWM1/RemaTxNum[18]_keep ),
    .o(pnumcnt1[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[19]  (
    .i(\PWM1/RemaTxNum[19]_keep ),
    .o(pnumcnt1[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[1]  (
    .i(\PWM1/RemaTxNum[1]_keep ),
    .o(pnumcnt1[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[20]  (
    .i(\PWM1/RemaTxNum[20]_keep ),
    .o(pnumcnt1[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[21]  (
    .i(\PWM1/RemaTxNum[21]_keep ),
    .o(pnumcnt1[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[22]  (
    .i(\PWM1/RemaTxNum[22]_keep ),
    .o(pnumcnt1[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[23]  (
    .i(\PWM1/RemaTxNum[23]_keep ),
    .o(pnumcnt1[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[2]  (
    .i(\PWM1/RemaTxNum[2]_keep ),
    .o(pnumcnt1[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[3]  (
    .i(\PWM1/RemaTxNum[3]_keep ),
    .o(pnumcnt1[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[4]  (
    .i(\PWM1/RemaTxNum[4]_keep ),
    .o(pnumcnt1[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[5]  (
    .i(\PWM1/RemaTxNum[5]_keep ),
    .o(pnumcnt1[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[6]  (
    .i(\PWM1/RemaTxNum[6]_keep ),
    .o(pnumcnt1[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[7]  (
    .i(\PWM1/RemaTxNum[7]_keep ),
    .o(pnumcnt1[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[8]  (
    .i(\PWM1/RemaTxNum[8]_keep ),
    .o(pnumcnt1[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_RemaTxNum[9]  (
    .i(\PWM1/RemaTxNum[9]_keep ),
    .o(pnumcnt1[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_dir  (
    .i(\PWM1/dir_keep ),
    .o(dir[1]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[0]  (
    .i(\PWM1/pnumr[0]_keep ),
    .o(\PWM1/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[10]  (
    .i(\PWM1/pnumr[10]_keep ),
    .o(\PWM1/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[11]  (
    .i(\PWM1/pnumr[11]_keep ),
    .o(\PWM1/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[12]  (
    .i(\PWM1/pnumr[12]_keep ),
    .o(\PWM1/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[13]  (
    .i(\PWM1/pnumr[13]_keep ),
    .o(\PWM1/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[14]  (
    .i(\PWM1/pnumr[14]_keep ),
    .o(\PWM1/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[15]  (
    .i(\PWM1/pnumr[15]_keep ),
    .o(\PWM1/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[16]  (
    .i(\PWM1/pnumr[16]_keep ),
    .o(\PWM1/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[17]  (
    .i(\PWM1/pnumr[17]_keep ),
    .o(\PWM1/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[18]  (
    .i(\PWM1/pnumr[18]_keep ),
    .o(\PWM1/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[19]  (
    .i(\PWM1/pnumr[19]_keep ),
    .o(\PWM1/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[1]  (
    .i(\PWM1/pnumr[1]_keep ),
    .o(\PWM1/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[20]  (
    .i(\PWM1/pnumr[20]_keep ),
    .o(\PWM1/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[21]  (
    .i(\PWM1/pnumr[21]_keep ),
    .o(\PWM1/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[22]  (
    .i(\PWM1/pnumr[22]_keep ),
    .o(\PWM1/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[23]  (
    .i(\PWM1/pnumr[23]_keep ),
    .o(\PWM1/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[24]  (
    .i(\PWM1/pnumr[24]_keep ),
    .o(\PWM1/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[25]  (
    .i(\PWM1/pnumr[25]_keep ),
    .o(\PWM1/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[26]  (
    .i(\PWM1/pnumr[26]_keep ),
    .o(\PWM1/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[27]  (
    .i(\PWM1/pnumr[27]_keep ),
    .o(\PWM1/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[28]  (
    .i(\PWM1/pnumr[28]_keep ),
    .o(\PWM1/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[29]  (
    .i(\PWM1/pnumr[29]_keep ),
    .o(\PWM1/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[2]  (
    .i(\PWM1/pnumr[2]_keep ),
    .o(\PWM1/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[30]  (
    .i(\PWM1/pnumr[30]_keep ),
    .o(\PWM1/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[31]  (
    .i(\PWM1/pnumr[31]_keep ),
    .o(\PWM1/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[3]  (
    .i(\PWM1/pnumr[3]_keep ),
    .o(\PWM1/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[4]  (
    .i(\PWM1/pnumr[4]_keep ),
    .o(\PWM1/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[5]  (
    .i(\PWM1/pnumr[5]_keep ),
    .o(\PWM1/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[6]  (
    .i(\PWM1/pnumr[6]_keep ),
    .o(\PWM1/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[7]  (
    .i(\PWM1/pnumr[7]_keep ),
    .o(\PWM1/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[8]  (
    .i(\PWM1/pnumr[8]_keep ),
    .o(\PWM1/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pnumr[9]  (
    .i(\PWM1/pnumr[9]_keep ),
    .o(\PWM1/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_pwm  (
    .i(\PWM1/pwm_keep ),
    .o(pwm[1]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM1/_bufkeep_stopreq  (
    .i(\PWM1/stopreq_keep ),
    .o(\PWM1/stopreq ));  // src/OnePWM.v(14)
  reg_ar_as_w1 \PWM1/dir_reg  (
    .clk(clk100m),
    .d(\PWM1/n32 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/dir_keep ));  // src/OnePWM.v(58)
  eq_w27 \PWM1/eq0  (
    .i0(\PWM1/FreCnt ),
    .i1(27'b000000000000000000000000000),
    .o(\PWM1/n0 ));  // src/OnePWM.v(15)
  eq_w24 \PWM1/eq1  (
    .i0(pnumcnt1),
    .i1(24'b000000000000000000000001),
    .o(\PWM1/n5 ));  // src/OnePWM.v(25)
  eq_w27 \PWM1/eq2  (
    .i0(\PWM1/FreCnt ),
    .i1({1'b0,\PWM1/FreCntr [26:1]}),
    .o(\PWM1/n17 ));  // src/OnePWM.v(41)
  eq_w27 \PWM1/eq3  (
    .i0(\PWM1/FreCnt ),
    .i1(\PWM1/FreCntr ),
    .o(\PWM1/n18 ));  // src/OnePWM.v(43)
  binary_mux_s1_w1 \PWM1/mux0_b0  (
    .i0(\PWM1/n12 [0]),
    .i1(freq1[0]),
    .sel(\PWM1/n0 ),
    .o(\PWM1/n13 [0]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM1/mux0_b1  (
    .i0(\PWM1/n12 [1]),
    .i1(freq1[1]),
    .sel(\PWM1/n0 ),
    .o(\PWM1/n13 [1]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM1/mux0_b10  (
    .i0(\PWM1/n12 [10]),
    .i1(freq1[10]),
    .sel(\PWM1/n0 ),
    .o(\PWM1/n13 [10]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM1/mux0_b11  (
    .i0(\PWM1/n12 [11]),
    .i1(freq1[11]),
    .sel(\PWM1/n0 ),
    .o(\PWM1/n13 [11]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM1/mux0_b12  (
    .i0(\PWM1/n12 [12]),
    .i1(freq1[12]),
    .sel(\PWM1/n0 ),
    .o(\PWM1/n13 [12]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM1/mux0_b13  (
    .i0(\PWM1/n12 [13]),
    .i1(freq1[13]),
    .sel(\PWM1/n0 ),
    .o(\PWM1/n13 [13]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM1/mux0_b14  (
    .i0(\PWM1/n12 [14]),
    .i1(freq1[14]),
    .sel(\PWM1/n0 ),
    .o(\PWM1/n13 [14]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM1/mux0_b15  (
    .i0(\PWM1/n12 [15]),
    .i1(freq1[15]),
    .sel(\PWM1/n0 ),
    .o(\PWM1/n13 [15]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM1/mux0_b16  (
    .i0(\PWM1/n12 [16]),
    .i1(freq1[16]),
    .sel(\PWM1/n0 ),
    .o(\PWM1/n13 [16]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM1/mux0_b17  (
    .i0(\PWM1/n12 [17]),
    .i1(freq1[17]),
    .sel(\PWM1/n0 ),
    .o(\PWM1/n13 [17]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM1/mux0_b18  (
    .i0(\PWM1/n12 [18]),
    .i1(freq1[18]),
    .sel(\PWM1/n0 ),
    .o(\PWM1/n13 [18]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM1/mux0_b19  (
    .i0(\PWM1/n12 [19]),
    .i1(freq1[19]),
    .sel(\PWM1/n0 ),
    .o(\PWM1/n13 [19]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM1/mux0_b2  (
    .i0(\PWM1/n12 [2]),
    .i1(freq1[2]),
    .sel(\PWM1/n0 ),
    .o(\PWM1/n13 [2]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM1/mux0_b20  (
    .i0(\PWM1/n12 [20]),
    .i1(freq1[20]),
    .sel(\PWM1/n0 ),
    .o(\PWM1/n13 [20]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM1/mux0_b21  (
    .i0(\PWM1/n12 [21]),
    .i1(freq1[21]),
    .sel(\PWM1/n0 ),
    .o(\PWM1/n13 [21]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM1/mux0_b22  (
    .i0(\PWM1/n12 [22]),
    .i1(freq1[22]),
    .sel(\PWM1/n0 ),
    .o(\PWM1/n13 [22]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM1/mux0_b23  (
    .i0(\PWM1/n12 [23]),
    .i1(freq1[23]),
    .sel(\PWM1/n0 ),
    .o(\PWM1/n13 [23]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM1/mux0_b24  (
    .i0(\PWM1/n12 [24]),
    .i1(freq1[24]),
    .sel(\PWM1/n0 ),
    .o(\PWM1/n13 [24]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM1/mux0_b25  (
    .i0(\PWM1/n12 [25]),
    .i1(freq1[25]),
    .sel(\PWM1/n0 ),
    .o(\PWM1/n13 [25]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM1/mux0_b26  (
    .i0(\PWM1/n12 [26]),
    .i1(freq1[26]),
    .sel(\PWM1/n0 ),
    .o(\PWM1/n13 [26]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM1/mux0_b3  (
    .i0(\PWM1/n12 [3]),
    .i1(freq1[3]),
    .sel(\PWM1/n0 ),
    .o(\PWM1/n13 [3]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM1/mux0_b4  (
    .i0(\PWM1/n12 [4]),
    .i1(freq1[4]),
    .sel(\PWM1/n0 ),
    .o(\PWM1/n13 [4]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM1/mux0_b5  (
    .i0(\PWM1/n12 [5]),
    .i1(freq1[5]),
    .sel(\PWM1/n0 ),
    .o(\PWM1/n13 [5]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM1/mux0_b6  (
    .i0(\PWM1/n12 [6]),
    .i1(freq1[6]),
    .sel(\PWM1/n0 ),
    .o(\PWM1/n13 [6]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM1/mux0_b7  (
    .i0(\PWM1/n12 [7]),
    .i1(freq1[7]),
    .sel(\PWM1/n0 ),
    .o(\PWM1/n13 [7]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM1/mux0_b8  (
    .i0(\PWM1/n12 [8]),
    .i1(freq1[8]),
    .sel(\PWM1/n0 ),
    .o(\PWM1/n13 [8]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM1/mux0_b9  (
    .i0(\PWM1/n12 [9]),
    .i1(freq1[9]),
    .sel(\PWM1/n0 ),
    .o(\PWM1/n13 [9]));  // src/OnePWM.v(32)
  and \PWM1/mux3_b0_sel_is_3  (\PWM1/mux3_b0_sel_is_3_o , \PWM1/n11 , \PWM1/n0 );
  binary_mux_s1_w1 \PWM1/mux4_b0  (
    .i0(\PWM1/pnumr [0]),
    .i1(1'b0),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n22 [0]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux4_b1  (
    .i0(\PWM1/pnumr [1]),
    .i1(1'b0),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n22 [1]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux4_b10  (
    .i0(\PWM1/pnumr [10]),
    .i1(1'b0),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n22 [10]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux4_b11  (
    .i0(\PWM1/pnumr [11]),
    .i1(1'b0),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n22 [11]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux4_b12  (
    .i0(\PWM1/pnumr [12]),
    .i1(1'b0),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n22 [12]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux4_b13  (
    .i0(\PWM1/pnumr [13]),
    .i1(1'b0),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n22 [13]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux4_b14  (
    .i0(\PWM1/pnumr [14]),
    .i1(1'b0),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n22 [14]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux4_b15  (
    .i0(\PWM1/pnumr [15]),
    .i1(1'b0),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n22 [15]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux4_b16  (
    .i0(\PWM1/pnumr [16]),
    .i1(1'b0),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n22 [16]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux4_b17  (
    .i0(\PWM1/pnumr [17]),
    .i1(1'b0),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n22 [17]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux4_b18  (
    .i0(\PWM1/pnumr [18]),
    .i1(1'b0),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n22 [18]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux4_b19  (
    .i0(\PWM1/pnumr [19]),
    .i1(1'b0),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n22 [19]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux4_b2  (
    .i0(\PWM1/pnumr [2]),
    .i1(1'b0),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n22 [2]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux4_b20  (
    .i0(\PWM1/pnumr [20]),
    .i1(1'b0),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n22 [20]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux4_b21  (
    .i0(\PWM1/pnumr [21]),
    .i1(1'b0),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n22 [21]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux4_b22  (
    .i0(\PWM1/pnumr [22]),
    .i1(1'b0),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n22 [22]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux4_b23  (
    .i0(\PWM1/pnumr [23]),
    .i1(1'b0),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n22 [23]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux4_b24  (
    .i0(\PWM1/pnumr [24]),
    .i1(1'b0),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n22 [24]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux4_b25  (
    .i0(\PWM1/pnumr [25]),
    .i1(1'b0),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n22 [25]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux4_b26  (
    .i0(\PWM1/pnumr [26]),
    .i1(1'b0),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n22 [26]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux4_b27  (
    .i0(\PWM1/pnumr [27]),
    .i1(1'b0),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n22 [27]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux4_b28  (
    .i0(\PWM1/pnumr [28]),
    .i1(1'b0),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n22 [28]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux4_b29  (
    .i0(\PWM1/pnumr [29]),
    .i1(1'b0),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n22 [29]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux4_b3  (
    .i0(\PWM1/pnumr [3]),
    .i1(1'b0),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n22 [3]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux4_b30  (
    .i0(\PWM1/pnumr [30]),
    .i1(1'b0),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n22 [30]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux4_b31  (
    .i0(\PWM1/pnumr [31]),
    .i1(1'b0),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n22 [31]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux4_b4  (
    .i0(\PWM1/pnumr [4]),
    .i1(1'b0),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n22 [4]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux4_b5  (
    .i0(\PWM1/pnumr [5]),
    .i1(1'b0),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n22 [5]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux4_b6  (
    .i0(\PWM1/pnumr [6]),
    .i1(1'b0),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n22 [6]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux4_b7  (
    .i0(\PWM1/pnumr [7]),
    .i1(1'b0),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n22 [7]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux4_b8  (
    .i0(\PWM1/pnumr [8]),
    .i1(1'b0),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n22 [8]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux4_b9  (
    .i0(\PWM1/pnumr [9]),
    .i1(1'b0),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n22 [9]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux5_b0  (
    .i0(\PWM1/n22 [0]),
    .i1(pnum1[0]),
    .sel(pnum1[32]),
    .o(\PWM1/n23 [0]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux5_b1  (
    .i0(\PWM1/n22 [1]),
    .i1(pnum1[1]),
    .sel(pnum1[32]),
    .o(\PWM1/n23 [1]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux5_b10  (
    .i0(\PWM1/n22 [10]),
    .i1(pnum1[10]),
    .sel(pnum1[32]),
    .o(\PWM1/n23 [10]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux5_b11  (
    .i0(\PWM1/n22 [11]),
    .i1(pnum1[11]),
    .sel(pnum1[32]),
    .o(\PWM1/n23 [11]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux5_b12  (
    .i0(\PWM1/n22 [12]),
    .i1(pnum1[12]),
    .sel(pnum1[32]),
    .o(\PWM1/n23 [12]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux5_b13  (
    .i0(\PWM1/n22 [13]),
    .i1(pnum1[13]),
    .sel(pnum1[32]),
    .o(\PWM1/n23 [13]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux5_b14  (
    .i0(\PWM1/n22 [14]),
    .i1(pnum1[14]),
    .sel(pnum1[32]),
    .o(\PWM1/n23 [14]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux5_b15  (
    .i0(\PWM1/n22 [15]),
    .i1(pnum1[15]),
    .sel(pnum1[32]),
    .o(\PWM1/n23 [15]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux5_b16  (
    .i0(\PWM1/n22 [16]),
    .i1(pnum1[16]),
    .sel(pnum1[32]),
    .o(\PWM1/n23 [16]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux5_b17  (
    .i0(\PWM1/n22 [17]),
    .i1(pnum1[17]),
    .sel(pnum1[32]),
    .o(\PWM1/n23 [17]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux5_b18  (
    .i0(\PWM1/n22 [18]),
    .i1(pnum1[18]),
    .sel(pnum1[32]),
    .o(\PWM1/n23 [18]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux5_b19  (
    .i0(\PWM1/n22 [19]),
    .i1(pnum1[19]),
    .sel(pnum1[32]),
    .o(\PWM1/n23 [19]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux5_b2  (
    .i0(\PWM1/n22 [2]),
    .i1(pnum1[2]),
    .sel(pnum1[32]),
    .o(\PWM1/n23 [2]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux5_b20  (
    .i0(\PWM1/n22 [20]),
    .i1(pnum1[20]),
    .sel(pnum1[32]),
    .o(\PWM1/n23 [20]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux5_b21  (
    .i0(\PWM1/n22 [21]),
    .i1(pnum1[21]),
    .sel(pnum1[32]),
    .o(\PWM1/n23 [21]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux5_b22  (
    .i0(\PWM1/n22 [22]),
    .i1(pnum1[22]),
    .sel(pnum1[32]),
    .o(\PWM1/n23 [22]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux5_b23  (
    .i0(\PWM1/n22 [23]),
    .i1(pnum1[23]),
    .sel(pnum1[32]),
    .o(\PWM1/n23 [23]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux5_b24  (
    .i0(\PWM1/n22 [24]),
    .i1(pnum1[24]),
    .sel(pnum1[32]),
    .o(\PWM1/n23 [24]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux5_b25  (
    .i0(\PWM1/n22 [25]),
    .i1(pnum1[25]),
    .sel(pnum1[32]),
    .o(\PWM1/n23 [25]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux5_b26  (
    .i0(\PWM1/n22 [26]),
    .i1(pnum1[26]),
    .sel(pnum1[32]),
    .o(\PWM1/n23 [26]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux5_b27  (
    .i0(\PWM1/n22 [27]),
    .i1(pnum1[27]),
    .sel(pnum1[32]),
    .o(\PWM1/n23 [27]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux5_b28  (
    .i0(\PWM1/n22 [28]),
    .i1(pnum1[28]),
    .sel(pnum1[32]),
    .o(\PWM1/n23 [28]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux5_b29  (
    .i0(\PWM1/n22 [29]),
    .i1(pnum1[29]),
    .sel(pnum1[32]),
    .o(\PWM1/n23 [29]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux5_b3  (
    .i0(\PWM1/n22 [3]),
    .i1(pnum1[3]),
    .sel(pnum1[32]),
    .o(\PWM1/n23 [3]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux5_b30  (
    .i0(\PWM1/n22 [30]),
    .i1(pnum1[30]),
    .sel(pnum1[32]),
    .o(\PWM1/n23 [30]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux5_b31  (
    .i0(\PWM1/n22 [31]),
    .i1(pnum1[31]),
    .sel(pnum1[32]),
    .o(\PWM1/n23 [31]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux5_b4  (
    .i0(\PWM1/n22 [4]),
    .i1(pnum1[4]),
    .sel(pnum1[32]),
    .o(\PWM1/n23 [4]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux5_b5  (
    .i0(\PWM1/n22 [5]),
    .i1(pnum1[5]),
    .sel(pnum1[32]),
    .o(\PWM1/n23 [5]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux5_b6  (
    .i0(\PWM1/n22 [6]),
    .i1(pnum1[6]),
    .sel(pnum1[32]),
    .o(\PWM1/n23 [6]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux5_b7  (
    .i0(\PWM1/n22 [7]),
    .i1(pnum1[7]),
    .sel(pnum1[32]),
    .o(\PWM1/n23 [7]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux5_b8  (
    .i0(\PWM1/n22 [8]),
    .i1(pnum1[8]),
    .sel(pnum1[32]),
    .o(\PWM1/n23 [8]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux5_b9  (
    .i0(\PWM1/n22 [9]),
    .i1(pnum1[9]),
    .sel(pnum1[32]),
    .o(\PWM1/n23 [9]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM1/mux6_b0  (
    .i0(\PWM1/pnumr [0]),
    .i1(\PWM1/n26 [0]),
    .sel(\PWM1/n25 ),
    .o(\PWM1/n27 [0]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM1/mux6_b1  (
    .i0(\PWM1/pnumr [1]),
    .i1(\PWM1/n26 [1]),
    .sel(\PWM1/n25 ),
    .o(\PWM1/n27 [1]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM1/mux6_b10  (
    .i0(\PWM1/pnumr [10]),
    .i1(\PWM1/n26 [10]),
    .sel(\PWM1/n25 ),
    .o(\PWM1/n27 [10]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM1/mux6_b11  (
    .i0(\PWM1/pnumr [11]),
    .i1(\PWM1/n26 [11]),
    .sel(\PWM1/n25 ),
    .o(\PWM1/n27 [11]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM1/mux6_b12  (
    .i0(\PWM1/pnumr [12]),
    .i1(\PWM1/n26 [12]),
    .sel(\PWM1/n25 ),
    .o(\PWM1/n27 [12]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM1/mux6_b13  (
    .i0(\PWM1/pnumr [13]),
    .i1(\PWM1/n26 [13]),
    .sel(\PWM1/n25 ),
    .o(\PWM1/n27 [13]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM1/mux6_b14  (
    .i0(\PWM1/pnumr [14]),
    .i1(\PWM1/n26 [14]),
    .sel(\PWM1/n25 ),
    .o(\PWM1/n27 [14]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM1/mux6_b15  (
    .i0(\PWM1/pnumr [15]),
    .i1(\PWM1/n26 [15]),
    .sel(\PWM1/n25 ),
    .o(\PWM1/n27 [15]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM1/mux6_b16  (
    .i0(\PWM1/pnumr [16]),
    .i1(\PWM1/n26 [16]),
    .sel(\PWM1/n25 ),
    .o(\PWM1/n27 [16]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM1/mux6_b17  (
    .i0(\PWM1/pnumr [17]),
    .i1(\PWM1/n26 [17]),
    .sel(\PWM1/n25 ),
    .o(\PWM1/n27 [17]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM1/mux6_b18  (
    .i0(\PWM1/pnumr [18]),
    .i1(\PWM1/n26 [18]),
    .sel(\PWM1/n25 ),
    .o(\PWM1/n27 [18]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM1/mux6_b19  (
    .i0(\PWM1/pnumr [19]),
    .i1(\PWM1/n26 [19]),
    .sel(\PWM1/n25 ),
    .o(\PWM1/n27 [19]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM1/mux6_b2  (
    .i0(\PWM1/pnumr [2]),
    .i1(\PWM1/n26 [2]),
    .sel(\PWM1/n25 ),
    .o(\PWM1/n27 [2]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM1/mux6_b20  (
    .i0(\PWM1/pnumr [20]),
    .i1(\PWM1/n26 [20]),
    .sel(\PWM1/n25 ),
    .o(\PWM1/n27 [20]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM1/mux6_b21  (
    .i0(\PWM1/pnumr [21]),
    .i1(\PWM1/n26 [21]),
    .sel(\PWM1/n25 ),
    .o(\PWM1/n27 [21]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM1/mux6_b22  (
    .i0(\PWM1/pnumr [22]),
    .i1(\PWM1/n26 [22]),
    .sel(\PWM1/n25 ),
    .o(\PWM1/n27 [22]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM1/mux6_b23  (
    .i0(\PWM1/pnumr [23]),
    .i1(\PWM1/n26 [23]),
    .sel(\PWM1/n25 ),
    .o(\PWM1/n27 [23]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM1/mux6_b3  (
    .i0(\PWM1/pnumr [3]),
    .i1(\PWM1/n26 [3]),
    .sel(\PWM1/n25 ),
    .o(\PWM1/n27 [3]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM1/mux6_b4  (
    .i0(\PWM1/pnumr [4]),
    .i1(\PWM1/n26 [4]),
    .sel(\PWM1/n25 ),
    .o(\PWM1/n27 [4]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM1/mux6_b5  (
    .i0(\PWM1/pnumr [5]),
    .i1(\PWM1/n26 [5]),
    .sel(\PWM1/n25 ),
    .o(\PWM1/n27 [5]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM1/mux6_b6  (
    .i0(\PWM1/pnumr [6]),
    .i1(\PWM1/n26 [6]),
    .sel(\PWM1/n25 ),
    .o(\PWM1/n27 [6]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM1/mux6_b7  (
    .i0(\PWM1/pnumr [7]),
    .i1(\PWM1/n26 [7]),
    .sel(\PWM1/n25 ),
    .o(\PWM1/n27 [7]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM1/mux6_b8  (
    .i0(\PWM1/pnumr [8]),
    .i1(\PWM1/n26 [8]),
    .sel(\PWM1/n25 ),
    .o(\PWM1/n27 [8]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM1/mux6_b9  (
    .i0(\PWM1/pnumr [9]),
    .i1(\PWM1/n26 [9]),
    .sel(\PWM1/n25 ),
    .o(\PWM1/n27 [9]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM1/mux7_b0  (
    .i0(pnumcnt1[0]),
    .i1(\PWM1/n27 [0]),
    .sel(\PWM1/n24 ),
    .o(\PWM1/n29 [0]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux7_b1  (
    .i0(pnumcnt1[1]),
    .i1(\PWM1/n27 [1]),
    .sel(\PWM1/n24 ),
    .o(\PWM1/n29 [1]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux7_b10  (
    .i0(pnumcnt1[10]),
    .i1(\PWM1/n27 [10]),
    .sel(\PWM1/n24 ),
    .o(\PWM1/n29 [10]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux7_b11  (
    .i0(pnumcnt1[11]),
    .i1(\PWM1/n27 [11]),
    .sel(\PWM1/n24 ),
    .o(\PWM1/n29 [11]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux7_b12  (
    .i0(pnumcnt1[12]),
    .i1(\PWM1/n27 [12]),
    .sel(\PWM1/n24 ),
    .o(\PWM1/n29 [12]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux7_b13  (
    .i0(pnumcnt1[13]),
    .i1(\PWM1/n27 [13]),
    .sel(\PWM1/n24 ),
    .o(\PWM1/n29 [13]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux7_b14  (
    .i0(pnumcnt1[14]),
    .i1(\PWM1/n27 [14]),
    .sel(\PWM1/n24 ),
    .o(\PWM1/n29 [14]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux7_b15  (
    .i0(pnumcnt1[15]),
    .i1(\PWM1/n27 [15]),
    .sel(\PWM1/n24 ),
    .o(\PWM1/n29 [15]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux7_b16  (
    .i0(pnumcnt1[16]),
    .i1(\PWM1/n27 [16]),
    .sel(\PWM1/n24 ),
    .o(\PWM1/n29 [16]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux7_b17  (
    .i0(pnumcnt1[17]),
    .i1(\PWM1/n27 [17]),
    .sel(\PWM1/n24 ),
    .o(\PWM1/n29 [17]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux7_b18  (
    .i0(pnumcnt1[18]),
    .i1(\PWM1/n27 [18]),
    .sel(\PWM1/n24 ),
    .o(\PWM1/n29 [18]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux7_b19  (
    .i0(pnumcnt1[19]),
    .i1(\PWM1/n27 [19]),
    .sel(\PWM1/n24 ),
    .o(\PWM1/n29 [19]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux7_b2  (
    .i0(pnumcnt1[2]),
    .i1(\PWM1/n27 [2]),
    .sel(\PWM1/n24 ),
    .o(\PWM1/n29 [2]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux7_b20  (
    .i0(pnumcnt1[20]),
    .i1(\PWM1/n27 [20]),
    .sel(\PWM1/n24 ),
    .o(\PWM1/n29 [20]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux7_b21  (
    .i0(pnumcnt1[21]),
    .i1(\PWM1/n27 [21]),
    .sel(\PWM1/n24 ),
    .o(\PWM1/n29 [21]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux7_b22  (
    .i0(pnumcnt1[22]),
    .i1(\PWM1/n27 [22]),
    .sel(\PWM1/n24 ),
    .o(\PWM1/n29 [22]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux7_b23  (
    .i0(pnumcnt1[23]),
    .i1(\PWM1/n27 [23]),
    .sel(\PWM1/n24 ),
    .o(\PWM1/n29 [23]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux7_b3  (
    .i0(pnumcnt1[3]),
    .i1(\PWM1/n27 [3]),
    .sel(\PWM1/n24 ),
    .o(\PWM1/n29 [3]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux7_b4  (
    .i0(pnumcnt1[4]),
    .i1(\PWM1/n27 [4]),
    .sel(\PWM1/n24 ),
    .o(\PWM1/n29 [4]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux7_b5  (
    .i0(pnumcnt1[5]),
    .i1(\PWM1/n27 [5]),
    .sel(\PWM1/n24 ),
    .o(\PWM1/n29 [5]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux7_b6  (
    .i0(pnumcnt1[6]),
    .i1(\PWM1/n27 [6]),
    .sel(\PWM1/n24 ),
    .o(\PWM1/n29 [6]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux7_b7  (
    .i0(pnumcnt1[7]),
    .i1(\PWM1/n27 [7]),
    .sel(\PWM1/n24 ),
    .o(\PWM1/n29 [7]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux7_b8  (
    .i0(pnumcnt1[8]),
    .i1(\PWM1/n27 [8]),
    .sel(\PWM1/n24 ),
    .o(\PWM1/n29 [8]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux7_b9  (
    .i0(pnumcnt1[9]),
    .i1(\PWM1/n27 [9]),
    .sel(\PWM1/n24 ),
    .o(\PWM1/n29 [9]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux8_b0  (
    .i0(\PWM1/n29 [0]),
    .i1(\PWM1/pnumr [0]),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n31 [0]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux8_b1  (
    .i0(\PWM1/n29 [1]),
    .i1(\PWM1/pnumr [1]),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n31 [1]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux8_b10  (
    .i0(\PWM1/n29 [10]),
    .i1(\PWM1/pnumr [10]),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n31 [10]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux8_b11  (
    .i0(\PWM1/n29 [11]),
    .i1(\PWM1/pnumr [11]),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n31 [11]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux8_b12  (
    .i0(\PWM1/n29 [12]),
    .i1(\PWM1/pnumr [12]),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n31 [12]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux8_b13  (
    .i0(\PWM1/n29 [13]),
    .i1(\PWM1/pnumr [13]),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n31 [13]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux8_b14  (
    .i0(\PWM1/n29 [14]),
    .i1(\PWM1/pnumr [14]),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n31 [14]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux8_b15  (
    .i0(\PWM1/n29 [15]),
    .i1(\PWM1/pnumr [15]),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n31 [15]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux8_b16  (
    .i0(\PWM1/n29 [16]),
    .i1(\PWM1/pnumr [16]),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n31 [16]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux8_b17  (
    .i0(\PWM1/n29 [17]),
    .i1(\PWM1/pnumr [17]),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n31 [17]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux8_b18  (
    .i0(\PWM1/n29 [18]),
    .i1(\PWM1/pnumr [18]),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n31 [18]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux8_b19  (
    .i0(\PWM1/n29 [19]),
    .i1(\PWM1/pnumr [19]),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n31 [19]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux8_b2  (
    .i0(\PWM1/n29 [2]),
    .i1(\PWM1/pnumr [2]),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n31 [2]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux8_b20  (
    .i0(\PWM1/n29 [20]),
    .i1(\PWM1/pnumr [20]),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n31 [20]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux8_b21  (
    .i0(\PWM1/n29 [21]),
    .i1(\PWM1/pnumr [21]),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n31 [21]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux8_b22  (
    .i0(\PWM1/n29 [22]),
    .i1(\PWM1/pnumr [22]),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n31 [22]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux8_b23  (
    .i0(\PWM1/n29 [23]),
    .i1(\PWM1/pnumr [23]),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n31 [23]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux8_b3  (
    .i0(\PWM1/n29 [3]),
    .i1(\PWM1/pnumr [3]),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n31 [3]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux8_b4  (
    .i0(\PWM1/n29 [4]),
    .i1(\PWM1/pnumr [4]),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n31 [4]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux8_b5  (
    .i0(\PWM1/n29 [5]),
    .i1(\PWM1/pnumr [5]),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n31 [5]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux8_b6  (
    .i0(\PWM1/n29 [6]),
    .i1(\PWM1/pnumr [6]),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n31 [6]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux8_b7  (
    .i0(\PWM1/n29 [7]),
    .i1(\PWM1/pnumr [7]),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n31 [7]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux8_b8  (
    .i0(\PWM1/n29 [8]),
    .i1(\PWM1/pnumr [8]),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n31 [8]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM1/mux8_b9  (
    .i0(\PWM1/n29 [9]),
    .i1(\PWM1/pnumr [9]),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n31 [9]));  // src/OnePWM.v(57)
  not \PWM1/n17_inv  (\PWM1/n17_neg , \PWM1/n17 );
  not \PWM1/n25_inv  (\PWM1/n25_neg , \PWM1/n25 );
  not \PWM1/n4_inv  (\PWM1/n4_neg , \PWM1/n4 );
  not \PWM1/n6_inv  (\PWM1/n6_neg , \PWM1/n6 );
  ne_w24 \PWM1/neq0  (
    .i0(pnumcnt1),
    .i1(24'b000000000000000000000000),
    .o(\PWM1/n25 ));  // src/OnePWM.v(55)
  reg_sr_ss_w1 \PWM1/pwm_reg  (
    .clk(clk100m),
    .d(pwm[1]),
    .en(1'b1),
    .reset(~\PWM1/u14_sel_is_1_o ),
    .set(\PWM1/n18 ),
    .q(\PWM1/pwm_keep ));  // src/OnePWM.v(45)
  reg_sr_as_w1 \PWM1/reg0_b0  (
    .clk(clk100m),
    .d(\PWM1/n13 [0]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [0]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b1  (
    .clk(clk100m),
    .d(\PWM1/n13 [1]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [1]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b10  (
    .clk(clk100m),
    .d(\PWM1/n13 [10]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [10]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b11  (
    .clk(clk100m),
    .d(\PWM1/n13 [11]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [11]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b12  (
    .clk(clk100m),
    .d(\PWM1/n13 [12]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [12]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b13  (
    .clk(clk100m),
    .d(\PWM1/n13 [13]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [13]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b14  (
    .clk(clk100m),
    .d(\PWM1/n13 [14]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [14]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b15  (
    .clk(clk100m),
    .d(\PWM1/n13 [15]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [15]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b16  (
    .clk(clk100m),
    .d(\PWM1/n13 [16]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [16]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b17  (
    .clk(clk100m),
    .d(\PWM1/n13 [17]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [17]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b18  (
    .clk(clk100m),
    .d(\PWM1/n13 [18]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [18]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b19  (
    .clk(clk100m),
    .d(\PWM1/n13 [19]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [19]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b2  (
    .clk(clk100m),
    .d(\PWM1/n13 [2]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [2]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b20  (
    .clk(clk100m),
    .d(\PWM1/n13 [20]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [20]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b21  (
    .clk(clk100m),
    .d(\PWM1/n13 [21]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [21]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b22  (
    .clk(clk100m),
    .d(\PWM1/n13 [22]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [22]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b23  (
    .clk(clk100m),
    .d(\PWM1/n13 [23]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [23]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b24  (
    .clk(clk100m),
    .d(\PWM1/n13 [24]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [24]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b25  (
    .clk(clk100m),
    .d(\PWM1/n13 [25]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [25]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b26  (
    .clk(clk100m),
    .d(\PWM1/n13 [26]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [26]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b3  (
    .clk(clk100m),
    .d(\PWM1/n13 [3]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [3]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b4  (
    .clk(clk100m),
    .d(\PWM1/n13 [4]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [4]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b5  (
    .clk(clk100m),
    .d(\PWM1/n13 [5]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [5]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b6  (
    .clk(clk100m),
    .d(\PWM1/n13 [6]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [6]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b7  (
    .clk(clk100m),
    .d(\PWM1/n13 [7]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [7]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b8  (
    .clk(clk100m),
    .d(\PWM1/n13 [8]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [8]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM1/reg0_b9  (
    .clk(clk100m),
    .d(\PWM1/n13 [9]),
    .en(1'b1),
    .reset(~\PWM1/n11 ),
    .set(1'b0),
    .q(\PWM1/FreCnt [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b0  (
    .clk(clk100m),
    .d(freq1[0]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [0]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b1  (
    .clk(clk100m),
    .d(freq1[1]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [1]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b10  (
    .clk(clk100m),
    .d(freq1[10]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [10]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b11  (
    .clk(clk100m),
    .d(freq1[11]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [11]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b12  (
    .clk(clk100m),
    .d(freq1[12]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [12]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b13  (
    .clk(clk100m),
    .d(freq1[13]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [13]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b14  (
    .clk(clk100m),
    .d(freq1[14]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [14]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b15  (
    .clk(clk100m),
    .d(freq1[15]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [15]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b16  (
    .clk(clk100m),
    .d(freq1[16]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [16]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b17  (
    .clk(clk100m),
    .d(freq1[17]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [17]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b18  (
    .clk(clk100m),
    .d(freq1[18]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [18]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b19  (
    .clk(clk100m),
    .d(freq1[19]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [19]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b2  (
    .clk(clk100m),
    .d(freq1[2]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [2]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b20  (
    .clk(clk100m),
    .d(freq1[20]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [20]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b21  (
    .clk(clk100m),
    .d(freq1[21]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [21]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b22  (
    .clk(clk100m),
    .d(freq1[22]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [22]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b23  (
    .clk(clk100m),
    .d(freq1[23]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [23]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b24  (
    .clk(clk100m),
    .d(freq1[24]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [24]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b25  (
    .clk(clk100m),
    .d(freq1[25]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [25]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b26  (
    .clk(clk100m),
    .d(freq1[26]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [26]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b3  (
    .clk(clk100m),
    .d(freq1[3]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [3]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b4  (
    .clk(clk100m),
    .d(freq1[4]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [4]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b5  (
    .clk(clk100m),
    .d(freq1[5]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [5]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b6  (
    .clk(clk100m),
    .d(freq1[6]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [6]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b7  (
    .clk(clk100m),
    .d(freq1[7]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [7]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b8  (
    .clk(clk100m),
    .d(freq1[8]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [8]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg1_b9  (
    .clk(clk100m),
    .d(freq1[9]),
    .en(\PWM1/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/FreCntr [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM1/reg2_b0  (
    .clk(clk100m),
    .d(\PWM1/n23 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[0]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b1  (
    .clk(clk100m),
    .d(\PWM1/n23 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[1]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b10  (
    .clk(clk100m),
    .d(\PWM1/n23 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[10]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b11  (
    .clk(clk100m),
    .d(\PWM1/n23 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[11]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b12  (
    .clk(clk100m),
    .d(\PWM1/n23 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[12]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b13  (
    .clk(clk100m),
    .d(\PWM1/n23 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[13]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b14  (
    .clk(clk100m),
    .d(\PWM1/n23 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[14]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b15  (
    .clk(clk100m),
    .d(\PWM1/n23 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[15]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b16  (
    .clk(clk100m),
    .d(\PWM1/n23 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[16]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b17  (
    .clk(clk100m),
    .d(\PWM1/n23 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[17]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b18  (
    .clk(clk100m),
    .d(\PWM1/n23 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[18]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b19  (
    .clk(clk100m),
    .d(\PWM1/n23 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[19]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b2  (
    .clk(clk100m),
    .d(\PWM1/n23 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[2]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b20  (
    .clk(clk100m),
    .d(\PWM1/n23 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[20]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b21  (
    .clk(clk100m),
    .d(\PWM1/n23 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[21]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b22  (
    .clk(clk100m),
    .d(\PWM1/n23 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[22]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b23  (
    .clk(clk100m),
    .d(\PWM1/n23 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[23]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b24  (
    .clk(clk100m),
    .d(\PWM1/n23 [24]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[24]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b25  (
    .clk(clk100m),
    .d(\PWM1/n23 [25]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[25]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b26  (
    .clk(clk100m),
    .d(\PWM1/n23 [26]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[26]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b27  (
    .clk(clk100m),
    .d(\PWM1/n23 [27]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[27]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b28  (
    .clk(clk100m),
    .d(\PWM1/n23 [28]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[28]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b29  (
    .clk(clk100m),
    .d(\PWM1/n23 [29]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[29]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b3  (
    .clk(clk100m),
    .d(\PWM1/n23 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[3]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b30  (
    .clk(clk100m),
    .d(\PWM1/n23 [30]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[30]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b31  (
    .clk(clk100m),
    .d(\PWM1/n23 [31]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[31]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b4  (
    .clk(clk100m),
    .d(\PWM1/n23 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[4]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b5  (
    .clk(clk100m),
    .d(\PWM1/n23 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[5]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b6  (
    .clk(clk100m),
    .d(\PWM1/n23 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[6]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b7  (
    .clk(clk100m),
    .d(\PWM1/n23 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[7]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b8  (
    .clk(clk100m),
    .d(\PWM1/n23 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[8]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg2_b9  (
    .clk(clk100m),
    .d(\PWM1/n23 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/pnumr[9]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM1/reg3_b0  (
    .clk(clk100m),
    .d(\PWM1/n31 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[0]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b1  (
    .clk(clk100m),
    .d(\PWM1/n31 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[1]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b10  (
    .clk(clk100m),
    .d(\PWM1/n31 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[10]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b11  (
    .clk(clk100m),
    .d(\PWM1/n31 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[11]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b12  (
    .clk(clk100m),
    .d(\PWM1/n31 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[12]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b13  (
    .clk(clk100m),
    .d(\PWM1/n31 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[13]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b14  (
    .clk(clk100m),
    .d(\PWM1/n31 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[14]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b15  (
    .clk(clk100m),
    .d(\PWM1/n31 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[15]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b16  (
    .clk(clk100m),
    .d(\PWM1/n31 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[16]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b17  (
    .clk(clk100m),
    .d(\PWM1/n31 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[17]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b18  (
    .clk(clk100m),
    .d(\PWM1/n31 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[18]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b19  (
    .clk(clk100m),
    .d(\PWM1/n31 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[19]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b2  (
    .clk(clk100m),
    .d(\PWM1/n31 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[2]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b20  (
    .clk(clk100m),
    .d(\PWM1/n31 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[20]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b21  (
    .clk(clk100m),
    .d(\PWM1/n31 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[21]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b22  (
    .clk(clk100m),
    .d(\PWM1/n31 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[22]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b23  (
    .clk(clk100m),
    .d(\PWM1/n31 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[23]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b3  (
    .clk(clk100m),
    .d(\PWM1/n31 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[3]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b4  (
    .clk(clk100m),
    .d(\PWM1/n31 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[4]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b5  (
    .clk(clk100m),
    .d(\PWM1/n31 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[5]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b6  (
    .clk(clk100m),
    .d(\PWM1/n31 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[6]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b7  (
    .clk(clk100m),
    .d(\PWM1/n31 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[7]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b8  (
    .clk(clk100m),
    .d(\PWM1/n31 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[8]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM1/reg3_b9  (
    .clk(clk100m),
    .d(\PWM1/n31 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM1/RemaTxNum[9]_keep ));  // src/OnePWM.v(58)
  reg_ar_ss_w1 \PWM1/stopreq_reg  (
    .clk(clk100m),
    .d(\PWM1/n1 ),
    .en(1'b1),
    .reset(1'b0),
    .set(pwm_start_stop[1]),
    .q(\PWM1/stopreq_keep ));  // src/OnePWM.v(15)
  add_pu27_mu27_o27 \PWM1/sub0  (
    .i0(\PWM1/FreCnt ),
    .i1(27'b000000000000000000000000001),
    .o(\PWM1/n12 [26:0]));  // src/OnePWM.v(32)
  add_pu24_mu24_o24 \PWM1/sub1  (
    .i0(pnumcnt1),
    .i1(24'b000000000000000000000001),
    .o(\PWM1/n26 [23:0]));  // src/OnePWM.v(55)
  AL_MUX \PWM1/u10  (
    .i0(1'b0),
    .i1(\PWM1/n9 ),
    .sel(n12),
    .o(\PWM1/n10 ));  // src/OnePWM.v(26)
  or \PWM1/u11  (\PWM1/n11 , pwm_state_read[1], pwm_start_stop[17]);  // src/OnePWM.v(30)
  and \PWM1/u14_sel_is_1  (\PWM1/u14_sel_is_1_o , pwm_state_read[1], \PWM1/n17_neg );
  and \PWM1/u15  (\PWM1/n24 , \PWM1/n0 , pwm_state_read[1]);  // src/OnePWM.v(54)
  and \PWM1/u17_sel_is_1  (\PWM1/u17_sel_is_1_o , \PWM1/n24 , \PWM1/n25_neg );
  not \PWM1/u17_sel_is_1_o_inv  (\PWM1/u17_sel_is_1_o_neg , \PWM1/u17_sel_is_1_o );
  AL_MUX \PWM1/u18  (
    .i0(\PWM1/pnumr [31]),
    .i1(dir[1]),
    .sel(\PWM1/u18_sel_is_0_o ),
    .o(\PWM1/n32 ));
  and \PWM1/u18_sel_is_0  (\PWM1/u18_sel_is_0_o , \pwm_start_stop[17]_neg , \PWM1/u17_sel_is_1_o_neg );
  AL_MUX \PWM1/u2  (
    .i0(\PWM1/stopreq ),
    .i1(1'b0),
    .sel(\PWM1/n0 ),
    .o(\PWM1/n1 ));  // src/OnePWM.v(15)
  and \PWM1/u5  (\PWM1/n4 , \PWM1/stopreq , \PWM1/n0 );  // src/OnePWM.v(23)
  and \PWM1/u6  (\PWM1/n6 , \PWM1/n5 , \PWM1/n0 );  // src/OnePWM.v(25)
  AL_MUX \PWM1/u8  (
    .i0(1'b0),
    .i1(pwm_state_read[1]),
    .sel(\PWM1/u8_sel_is_0_o ),
    .o(\PWM1/n8 ));
  and \PWM1/u8_sel_is_0  (\PWM1/u8_sel_is_0_o , \PWM1/n4_neg , \PWM1/n6_neg );
  AL_MUX \PWM1/u9  (
    .i0(\PWM1/n8 ),
    .i1(1'b1),
    .sel(pwm_start_stop[17]),
    .o(\PWM1/n9 ));  // src/OnePWM.v(26)
  reg_ar_as_w1 \PWM2/State_reg  (
    .clk(clk100m),
    .d(\PWM2/n10 ),
    .en(1'b1),
    .reset(~rstn),
    .set(1'b0),
    .q(pwm_state_read[2]));  // src/OnePWM.v(26)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[0]  (
    .i(\PWM2/RemaTxNum[0]_keep ),
    .o(pnumcnt2[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[10]  (
    .i(\PWM2/RemaTxNum[10]_keep ),
    .o(pnumcnt2[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[11]  (
    .i(\PWM2/RemaTxNum[11]_keep ),
    .o(pnumcnt2[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[12]  (
    .i(\PWM2/RemaTxNum[12]_keep ),
    .o(pnumcnt2[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[13]  (
    .i(\PWM2/RemaTxNum[13]_keep ),
    .o(pnumcnt2[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[14]  (
    .i(\PWM2/RemaTxNum[14]_keep ),
    .o(pnumcnt2[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[15]  (
    .i(\PWM2/RemaTxNum[15]_keep ),
    .o(pnumcnt2[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[16]  (
    .i(\PWM2/RemaTxNum[16]_keep ),
    .o(pnumcnt2[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[17]  (
    .i(\PWM2/RemaTxNum[17]_keep ),
    .o(pnumcnt2[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[18]  (
    .i(\PWM2/RemaTxNum[18]_keep ),
    .o(pnumcnt2[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[19]  (
    .i(\PWM2/RemaTxNum[19]_keep ),
    .o(pnumcnt2[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[1]  (
    .i(\PWM2/RemaTxNum[1]_keep ),
    .o(pnumcnt2[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[20]  (
    .i(\PWM2/RemaTxNum[20]_keep ),
    .o(pnumcnt2[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[21]  (
    .i(\PWM2/RemaTxNum[21]_keep ),
    .o(pnumcnt2[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[22]  (
    .i(\PWM2/RemaTxNum[22]_keep ),
    .o(pnumcnt2[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[23]  (
    .i(\PWM2/RemaTxNum[23]_keep ),
    .o(pnumcnt2[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[2]  (
    .i(\PWM2/RemaTxNum[2]_keep ),
    .o(pnumcnt2[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[3]  (
    .i(\PWM2/RemaTxNum[3]_keep ),
    .o(pnumcnt2[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[4]  (
    .i(\PWM2/RemaTxNum[4]_keep ),
    .o(pnumcnt2[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[5]  (
    .i(\PWM2/RemaTxNum[5]_keep ),
    .o(pnumcnt2[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[6]  (
    .i(\PWM2/RemaTxNum[6]_keep ),
    .o(pnumcnt2[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[7]  (
    .i(\PWM2/RemaTxNum[7]_keep ),
    .o(pnumcnt2[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[8]  (
    .i(\PWM2/RemaTxNum[8]_keep ),
    .o(pnumcnt2[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_RemaTxNum[9]  (
    .i(\PWM2/RemaTxNum[9]_keep ),
    .o(pnumcnt2[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_dir  (
    .i(\PWM2/dir_keep ),
    .o(dir[2]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[0]  (
    .i(\PWM2/pnumr[0]_keep ),
    .o(\PWM2/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[10]  (
    .i(\PWM2/pnumr[10]_keep ),
    .o(\PWM2/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[11]  (
    .i(\PWM2/pnumr[11]_keep ),
    .o(\PWM2/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[12]  (
    .i(\PWM2/pnumr[12]_keep ),
    .o(\PWM2/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[13]  (
    .i(\PWM2/pnumr[13]_keep ),
    .o(\PWM2/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[14]  (
    .i(\PWM2/pnumr[14]_keep ),
    .o(\PWM2/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[15]  (
    .i(\PWM2/pnumr[15]_keep ),
    .o(\PWM2/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[16]  (
    .i(\PWM2/pnumr[16]_keep ),
    .o(\PWM2/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[17]  (
    .i(\PWM2/pnumr[17]_keep ),
    .o(\PWM2/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[18]  (
    .i(\PWM2/pnumr[18]_keep ),
    .o(\PWM2/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[19]  (
    .i(\PWM2/pnumr[19]_keep ),
    .o(\PWM2/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[1]  (
    .i(\PWM2/pnumr[1]_keep ),
    .o(\PWM2/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[20]  (
    .i(\PWM2/pnumr[20]_keep ),
    .o(\PWM2/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[21]  (
    .i(\PWM2/pnumr[21]_keep ),
    .o(\PWM2/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[22]  (
    .i(\PWM2/pnumr[22]_keep ),
    .o(\PWM2/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[23]  (
    .i(\PWM2/pnumr[23]_keep ),
    .o(\PWM2/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[24]  (
    .i(\PWM2/pnumr[24]_keep ),
    .o(\PWM2/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[25]  (
    .i(\PWM2/pnumr[25]_keep ),
    .o(\PWM2/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[26]  (
    .i(\PWM2/pnumr[26]_keep ),
    .o(\PWM2/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[27]  (
    .i(\PWM2/pnumr[27]_keep ),
    .o(\PWM2/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[28]  (
    .i(\PWM2/pnumr[28]_keep ),
    .o(\PWM2/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[29]  (
    .i(\PWM2/pnumr[29]_keep ),
    .o(\PWM2/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[2]  (
    .i(\PWM2/pnumr[2]_keep ),
    .o(\PWM2/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[30]  (
    .i(\PWM2/pnumr[30]_keep ),
    .o(\PWM2/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[31]  (
    .i(\PWM2/pnumr[31]_keep ),
    .o(\PWM2/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[3]  (
    .i(\PWM2/pnumr[3]_keep ),
    .o(\PWM2/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[4]  (
    .i(\PWM2/pnumr[4]_keep ),
    .o(\PWM2/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[5]  (
    .i(\PWM2/pnumr[5]_keep ),
    .o(\PWM2/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[6]  (
    .i(\PWM2/pnumr[6]_keep ),
    .o(\PWM2/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[7]  (
    .i(\PWM2/pnumr[7]_keep ),
    .o(\PWM2/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[8]  (
    .i(\PWM2/pnumr[8]_keep ),
    .o(\PWM2/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pnumr[9]  (
    .i(\PWM2/pnumr[9]_keep ),
    .o(\PWM2/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_pwm  (
    .i(\PWM2/pwm_keep ),
    .o(pwm[2]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM2/_bufkeep_stopreq  (
    .i(\PWM2/stopreq_keep ),
    .o(\PWM2/stopreq ));  // src/OnePWM.v(14)
  reg_ar_as_w1 \PWM2/dir_reg  (
    .clk(clk100m),
    .d(\PWM2/n32 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/dir_keep ));  // src/OnePWM.v(58)
  eq_w27 \PWM2/eq0  (
    .i0(\PWM2/FreCnt ),
    .i1(27'b000000000000000000000000000),
    .o(\PWM2/n0 ));  // src/OnePWM.v(15)
  eq_w24 \PWM2/eq1  (
    .i0(pnumcnt2),
    .i1(24'b000000000000000000000001),
    .o(\PWM2/n5 ));  // src/OnePWM.v(25)
  eq_w27 \PWM2/eq2  (
    .i0(\PWM2/FreCnt ),
    .i1({1'b0,\PWM2/FreCntr [26:1]}),
    .o(\PWM2/n17 ));  // src/OnePWM.v(41)
  eq_w27 \PWM2/eq3  (
    .i0(\PWM2/FreCnt ),
    .i1(\PWM2/FreCntr ),
    .o(\PWM2/n18 ));  // src/OnePWM.v(43)
  binary_mux_s1_w1 \PWM2/mux0_b0  (
    .i0(\PWM2/n12 [0]),
    .i1(freq2[0]),
    .sel(\PWM2/n0 ),
    .o(\PWM2/n13 [0]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM2/mux0_b1  (
    .i0(\PWM2/n12 [1]),
    .i1(freq2[1]),
    .sel(\PWM2/n0 ),
    .o(\PWM2/n13 [1]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM2/mux0_b10  (
    .i0(\PWM2/n12 [10]),
    .i1(freq2[10]),
    .sel(\PWM2/n0 ),
    .o(\PWM2/n13 [10]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM2/mux0_b11  (
    .i0(\PWM2/n12 [11]),
    .i1(freq2[11]),
    .sel(\PWM2/n0 ),
    .o(\PWM2/n13 [11]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM2/mux0_b12  (
    .i0(\PWM2/n12 [12]),
    .i1(freq2[12]),
    .sel(\PWM2/n0 ),
    .o(\PWM2/n13 [12]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM2/mux0_b13  (
    .i0(\PWM2/n12 [13]),
    .i1(freq2[13]),
    .sel(\PWM2/n0 ),
    .o(\PWM2/n13 [13]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM2/mux0_b14  (
    .i0(\PWM2/n12 [14]),
    .i1(freq2[14]),
    .sel(\PWM2/n0 ),
    .o(\PWM2/n13 [14]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM2/mux0_b15  (
    .i0(\PWM2/n12 [15]),
    .i1(freq2[15]),
    .sel(\PWM2/n0 ),
    .o(\PWM2/n13 [15]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM2/mux0_b16  (
    .i0(\PWM2/n12 [16]),
    .i1(freq2[16]),
    .sel(\PWM2/n0 ),
    .o(\PWM2/n13 [16]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM2/mux0_b17  (
    .i0(\PWM2/n12 [17]),
    .i1(freq2[17]),
    .sel(\PWM2/n0 ),
    .o(\PWM2/n13 [17]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM2/mux0_b18  (
    .i0(\PWM2/n12 [18]),
    .i1(freq2[18]),
    .sel(\PWM2/n0 ),
    .o(\PWM2/n13 [18]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM2/mux0_b19  (
    .i0(\PWM2/n12 [19]),
    .i1(freq2[19]),
    .sel(\PWM2/n0 ),
    .o(\PWM2/n13 [19]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM2/mux0_b2  (
    .i0(\PWM2/n12 [2]),
    .i1(freq2[2]),
    .sel(\PWM2/n0 ),
    .o(\PWM2/n13 [2]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM2/mux0_b20  (
    .i0(\PWM2/n12 [20]),
    .i1(freq2[20]),
    .sel(\PWM2/n0 ),
    .o(\PWM2/n13 [20]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM2/mux0_b21  (
    .i0(\PWM2/n12 [21]),
    .i1(freq2[21]),
    .sel(\PWM2/n0 ),
    .o(\PWM2/n13 [21]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM2/mux0_b22  (
    .i0(\PWM2/n12 [22]),
    .i1(freq2[22]),
    .sel(\PWM2/n0 ),
    .o(\PWM2/n13 [22]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM2/mux0_b23  (
    .i0(\PWM2/n12 [23]),
    .i1(freq2[23]),
    .sel(\PWM2/n0 ),
    .o(\PWM2/n13 [23]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM2/mux0_b24  (
    .i0(\PWM2/n12 [24]),
    .i1(freq2[24]),
    .sel(\PWM2/n0 ),
    .o(\PWM2/n13 [24]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM2/mux0_b25  (
    .i0(\PWM2/n12 [25]),
    .i1(freq2[25]),
    .sel(\PWM2/n0 ),
    .o(\PWM2/n13 [25]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM2/mux0_b26  (
    .i0(\PWM2/n12 [26]),
    .i1(freq2[26]),
    .sel(\PWM2/n0 ),
    .o(\PWM2/n13 [26]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM2/mux0_b3  (
    .i0(\PWM2/n12 [3]),
    .i1(freq2[3]),
    .sel(\PWM2/n0 ),
    .o(\PWM2/n13 [3]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM2/mux0_b4  (
    .i0(\PWM2/n12 [4]),
    .i1(freq2[4]),
    .sel(\PWM2/n0 ),
    .o(\PWM2/n13 [4]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM2/mux0_b5  (
    .i0(\PWM2/n12 [5]),
    .i1(freq2[5]),
    .sel(\PWM2/n0 ),
    .o(\PWM2/n13 [5]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM2/mux0_b6  (
    .i0(\PWM2/n12 [6]),
    .i1(freq2[6]),
    .sel(\PWM2/n0 ),
    .o(\PWM2/n13 [6]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM2/mux0_b7  (
    .i0(\PWM2/n12 [7]),
    .i1(freq2[7]),
    .sel(\PWM2/n0 ),
    .o(\PWM2/n13 [7]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM2/mux0_b8  (
    .i0(\PWM2/n12 [8]),
    .i1(freq2[8]),
    .sel(\PWM2/n0 ),
    .o(\PWM2/n13 [8]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM2/mux0_b9  (
    .i0(\PWM2/n12 [9]),
    .i1(freq2[9]),
    .sel(\PWM2/n0 ),
    .o(\PWM2/n13 [9]));  // src/OnePWM.v(32)
  and \PWM2/mux3_b0_sel_is_3  (\PWM2/mux3_b0_sel_is_3_o , \PWM2/n11 , \PWM2/n0 );
  binary_mux_s1_w1 \PWM2/mux4_b0  (
    .i0(\PWM2/pnumr [0]),
    .i1(1'b0),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n22 [0]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux4_b1  (
    .i0(\PWM2/pnumr [1]),
    .i1(1'b0),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n22 [1]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux4_b10  (
    .i0(\PWM2/pnumr [10]),
    .i1(1'b0),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n22 [10]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux4_b11  (
    .i0(\PWM2/pnumr [11]),
    .i1(1'b0),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n22 [11]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux4_b12  (
    .i0(\PWM2/pnumr [12]),
    .i1(1'b0),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n22 [12]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux4_b13  (
    .i0(\PWM2/pnumr [13]),
    .i1(1'b0),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n22 [13]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux4_b14  (
    .i0(\PWM2/pnumr [14]),
    .i1(1'b0),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n22 [14]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux4_b15  (
    .i0(\PWM2/pnumr [15]),
    .i1(1'b0),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n22 [15]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux4_b16  (
    .i0(\PWM2/pnumr [16]),
    .i1(1'b0),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n22 [16]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux4_b17  (
    .i0(\PWM2/pnumr [17]),
    .i1(1'b0),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n22 [17]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux4_b18  (
    .i0(\PWM2/pnumr [18]),
    .i1(1'b0),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n22 [18]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux4_b19  (
    .i0(\PWM2/pnumr [19]),
    .i1(1'b0),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n22 [19]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux4_b2  (
    .i0(\PWM2/pnumr [2]),
    .i1(1'b0),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n22 [2]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux4_b20  (
    .i0(\PWM2/pnumr [20]),
    .i1(1'b0),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n22 [20]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux4_b21  (
    .i0(\PWM2/pnumr [21]),
    .i1(1'b0),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n22 [21]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux4_b22  (
    .i0(\PWM2/pnumr [22]),
    .i1(1'b0),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n22 [22]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux4_b23  (
    .i0(\PWM2/pnumr [23]),
    .i1(1'b0),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n22 [23]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux4_b24  (
    .i0(\PWM2/pnumr [24]),
    .i1(1'b0),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n22 [24]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux4_b25  (
    .i0(\PWM2/pnumr [25]),
    .i1(1'b0),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n22 [25]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux4_b26  (
    .i0(\PWM2/pnumr [26]),
    .i1(1'b0),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n22 [26]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux4_b27  (
    .i0(\PWM2/pnumr [27]),
    .i1(1'b0),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n22 [27]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux4_b28  (
    .i0(\PWM2/pnumr [28]),
    .i1(1'b0),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n22 [28]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux4_b29  (
    .i0(\PWM2/pnumr [29]),
    .i1(1'b0),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n22 [29]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux4_b3  (
    .i0(\PWM2/pnumr [3]),
    .i1(1'b0),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n22 [3]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux4_b30  (
    .i0(\PWM2/pnumr [30]),
    .i1(1'b0),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n22 [30]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux4_b31  (
    .i0(\PWM2/pnumr [31]),
    .i1(1'b0),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n22 [31]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux4_b4  (
    .i0(\PWM2/pnumr [4]),
    .i1(1'b0),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n22 [4]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux4_b5  (
    .i0(\PWM2/pnumr [5]),
    .i1(1'b0),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n22 [5]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux4_b6  (
    .i0(\PWM2/pnumr [6]),
    .i1(1'b0),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n22 [6]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux4_b7  (
    .i0(\PWM2/pnumr [7]),
    .i1(1'b0),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n22 [7]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux4_b8  (
    .i0(\PWM2/pnumr [8]),
    .i1(1'b0),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n22 [8]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux4_b9  (
    .i0(\PWM2/pnumr [9]),
    .i1(1'b0),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n22 [9]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux5_b0  (
    .i0(\PWM2/n22 [0]),
    .i1(pnum2[0]),
    .sel(pnum2[32]),
    .o(\PWM2/n23 [0]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux5_b1  (
    .i0(\PWM2/n22 [1]),
    .i1(pnum2[1]),
    .sel(pnum2[32]),
    .o(\PWM2/n23 [1]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux5_b10  (
    .i0(\PWM2/n22 [10]),
    .i1(pnum2[10]),
    .sel(pnum2[32]),
    .o(\PWM2/n23 [10]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux5_b11  (
    .i0(\PWM2/n22 [11]),
    .i1(pnum2[11]),
    .sel(pnum2[32]),
    .o(\PWM2/n23 [11]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux5_b12  (
    .i0(\PWM2/n22 [12]),
    .i1(pnum2[12]),
    .sel(pnum2[32]),
    .o(\PWM2/n23 [12]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux5_b13  (
    .i0(\PWM2/n22 [13]),
    .i1(pnum2[13]),
    .sel(pnum2[32]),
    .o(\PWM2/n23 [13]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux5_b14  (
    .i0(\PWM2/n22 [14]),
    .i1(pnum2[14]),
    .sel(pnum2[32]),
    .o(\PWM2/n23 [14]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux5_b15  (
    .i0(\PWM2/n22 [15]),
    .i1(pnum2[15]),
    .sel(pnum2[32]),
    .o(\PWM2/n23 [15]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux5_b16  (
    .i0(\PWM2/n22 [16]),
    .i1(pnum2[16]),
    .sel(pnum2[32]),
    .o(\PWM2/n23 [16]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux5_b17  (
    .i0(\PWM2/n22 [17]),
    .i1(pnum2[17]),
    .sel(pnum2[32]),
    .o(\PWM2/n23 [17]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux5_b18  (
    .i0(\PWM2/n22 [18]),
    .i1(pnum2[18]),
    .sel(pnum2[32]),
    .o(\PWM2/n23 [18]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux5_b19  (
    .i0(\PWM2/n22 [19]),
    .i1(pnum2[19]),
    .sel(pnum2[32]),
    .o(\PWM2/n23 [19]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux5_b2  (
    .i0(\PWM2/n22 [2]),
    .i1(pnum2[2]),
    .sel(pnum2[32]),
    .o(\PWM2/n23 [2]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux5_b20  (
    .i0(\PWM2/n22 [20]),
    .i1(pnum2[20]),
    .sel(pnum2[32]),
    .o(\PWM2/n23 [20]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux5_b21  (
    .i0(\PWM2/n22 [21]),
    .i1(pnum2[21]),
    .sel(pnum2[32]),
    .o(\PWM2/n23 [21]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux5_b22  (
    .i0(\PWM2/n22 [22]),
    .i1(pnum2[22]),
    .sel(pnum2[32]),
    .o(\PWM2/n23 [22]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux5_b23  (
    .i0(\PWM2/n22 [23]),
    .i1(pnum2[23]),
    .sel(pnum2[32]),
    .o(\PWM2/n23 [23]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux5_b24  (
    .i0(\PWM2/n22 [24]),
    .i1(pnum2[24]),
    .sel(pnum2[32]),
    .o(\PWM2/n23 [24]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux5_b25  (
    .i0(\PWM2/n22 [25]),
    .i1(pnum2[25]),
    .sel(pnum2[32]),
    .o(\PWM2/n23 [25]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux5_b26  (
    .i0(\PWM2/n22 [26]),
    .i1(pnum2[26]),
    .sel(pnum2[32]),
    .o(\PWM2/n23 [26]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux5_b27  (
    .i0(\PWM2/n22 [27]),
    .i1(pnum2[27]),
    .sel(pnum2[32]),
    .o(\PWM2/n23 [27]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux5_b28  (
    .i0(\PWM2/n22 [28]),
    .i1(pnum2[28]),
    .sel(pnum2[32]),
    .o(\PWM2/n23 [28]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux5_b29  (
    .i0(\PWM2/n22 [29]),
    .i1(pnum2[29]),
    .sel(pnum2[32]),
    .o(\PWM2/n23 [29]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux5_b3  (
    .i0(\PWM2/n22 [3]),
    .i1(pnum2[3]),
    .sel(pnum2[32]),
    .o(\PWM2/n23 [3]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux5_b30  (
    .i0(\PWM2/n22 [30]),
    .i1(pnum2[30]),
    .sel(pnum2[32]),
    .o(\PWM2/n23 [30]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux5_b31  (
    .i0(\PWM2/n22 [31]),
    .i1(pnum2[31]),
    .sel(pnum2[32]),
    .o(\PWM2/n23 [31]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux5_b4  (
    .i0(\PWM2/n22 [4]),
    .i1(pnum2[4]),
    .sel(pnum2[32]),
    .o(\PWM2/n23 [4]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux5_b5  (
    .i0(\PWM2/n22 [5]),
    .i1(pnum2[5]),
    .sel(pnum2[32]),
    .o(\PWM2/n23 [5]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux5_b6  (
    .i0(\PWM2/n22 [6]),
    .i1(pnum2[6]),
    .sel(pnum2[32]),
    .o(\PWM2/n23 [6]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux5_b7  (
    .i0(\PWM2/n22 [7]),
    .i1(pnum2[7]),
    .sel(pnum2[32]),
    .o(\PWM2/n23 [7]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux5_b8  (
    .i0(\PWM2/n22 [8]),
    .i1(pnum2[8]),
    .sel(pnum2[32]),
    .o(\PWM2/n23 [8]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux5_b9  (
    .i0(\PWM2/n22 [9]),
    .i1(pnum2[9]),
    .sel(pnum2[32]),
    .o(\PWM2/n23 [9]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM2/mux6_b0  (
    .i0(\PWM2/pnumr [0]),
    .i1(\PWM2/n26 [0]),
    .sel(\PWM2/n25 ),
    .o(\PWM2/n27 [0]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM2/mux6_b1  (
    .i0(\PWM2/pnumr [1]),
    .i1(\PWM2/n26 [1]),
    .sel(\PWM2/n25 ),
    .o(\PWM2/n27 [1]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM2/mux6_b10  (
    .i0(\PWM2/pnumr [10]),
    .i1(\PWM2/n26 [10]),
    .sel(\PWM2/n25 ),
    .o(\PWM2/n27 [10]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM2/mux6_b11  (
    .i0(\PWM2/pnumr [11]),
    .i1(\PWM2/n26 [11]),
    .sel(\PWM2/n25 ),
    .o(\PWM2/n27 [11]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM2/mux6_b12  (
    .i0(\PWM2/pnumr [12]),
    .i1(\PWM2/n26 [12]),
    .sel(\PWM2/n25 ),
    .o(\PWM2/n27 [12]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM2/mux6_b13  (
    .i0(\PWM2/pnumr [13]),
    .i1(\PWM2/n26 [13]),
    .sel(\PWM2/n25 ),
    .o(\PWM2/n27 [13]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM2/mux6_b14  (
    .i0(\PWM2/pnumr [14]),
    .i1(\PWM2/n26 [14]),
    .sel(\PWM2/n25 ),
    .o(\PWM2/n27 [14]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM2/mux6_b15  (
    .i0(\PWM2/pnumr [15]),
    .i1(\PWM2/n26 [15]),
    .sel(\PWM2/n25 ),
    .o(\PWM2/n27 [15]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM2/mux6_b16  (
    .i0(\PWM2/pnumr [16]),
    .i1(\PWM2/n26 [16]),
    .sel(\PWM2/n25 ),
    .o(\PWM2/n27 [16]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM2/mux6_b17  (
    .i0(\PWM2/pnumr [17]),
    .i1(\PWM2/n26 [17]),
    .sel(\PWM2/n25 ),
    .o(\PWM2/n27 [17]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM2/mux6_b18  (
    .i0(\PWM2/pnumr [18]),
    .i1(\PWM2/n26 [18]),
    .sel(\PWM2/n25 ),
    .o(\PWM2/n27 [18]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM2/mux6_b19  (
    .i0(\PWM2/pnumr [19]),
    .i1(\PWM2/n26 [19]),
    .sel(\PWM2/n25 ),
    .o(\PWM2/n27 [19]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM2/mux6_b2  (
    .i0(\PWM2/pnumr [2]),
    .i1(\PWM2/n26 [2]),
    .sel(\PWM2/n25 ),
    .o(\PWM2/n27 [2]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM2/mux6_b20  (
    .i0(\PWM2/pnumr [20]),
    .i1(\PWM2/n26 [20]),
    .sel(\PWM2/n25 ),
    .o(\PWM2/n27 [20]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM2/mux6_b21  (
    .i0(\PWM2/pnumr [21]),
    .i1(\PWM2/n26 [21]),
    .sel(\PWM2/n25 ),
    .o(\PWM2/n27 [21]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM2/mux6_b22  (
    .i0(\PWM2/pnumr [22]),
    .i1(\PWM2/n26 [22]),
    .sel(\PWM2/n25 ),
    .o(\PWM2/n27 [22]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM2/mux6_b23  (
    .i0(\PWM2/pnumr [23]),
    .i1(\PWM2/n26 [23]),
    .sel(\PWM2/n25 ),
    .o(\PWM2/n27 [23]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM2/mux6_b3  (
    .i0(\PWM2/pnumr [3]),
    .i1(\PWM2/n26 [3]),
    .sel(\PWM2/n25 ),
    .o(\PWM2/n27 [3]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM2/mux6_b4  (
    .i0(\PWM2/pnumr [4]),
    .i1(\PWM2/n26 [4]),
    .sel(\PWM2/n25 ),
    .o(\PWM2/n27 [4]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM2/mux6_b5  (
    .i0(\PWM2/pnumr [5]),
    .i1(\PWM2/n26 [5]),
    .sel(\PWM2/n25 ),
    .o(\PWM2/n27 [5]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM2/mux6_b6  (
    .i0(\PWM2/pnumr [6]),
    .i1(\PWM2/n26 [6]),
    .sel(\PWM2/n25 ),
    .o(\PWM2/n27 [6]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM2/mux6_b7  (
    .i0(\PWM2/pnumr [7]),
    .i1(\PWM2/n26 [7]),
    .sel(\PWM2/n25 ),
    .o(\PWM2/n27 [7]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM2/mux6_b8  (
    .i0(\PWM2/pnumr [8]),
    .i1(\PWM2/n26 [8]),
    .sel(\PWM2/n25 ),
    .o(\PWM2/n27 [8]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM2/mux6_b9  (
    .i0(\PWM2/pnumr [9]),
    .i1(\PWM2/n26 [9]),
    .sel(\PWM2/n25 ),
    .o(\PWM2/n27 [9]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM2/mux7_b0  (
    .i0(pnumcnt2[0]),
    .i1(\PWM2/n27 [0]),
    .sel(\PWM2/n24 ),
    .o(\PWM2/n29 [0]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux7_b1  (
    .i0(pnumcnt2[1]),
    .i1(\PWM2/n27 [1]),
    .sel(\PWM2/n24 ),
    .o(\PWM2/n29 [1]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux7_b10  (
    .i0(pnumcnt2[10]),
    .i1(\PWM2/n27 [10]),
    .sel(\PWM2/n24 ),
    .o(\PWM2/n29 [10]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux7_b11  (
    .i0(pnumcnt2[11]),
    .i1(\PWM2/n27 [11]),
    .sel(\PWM2/n24 ),
    .o(\PWM2/n29 [11]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux7_b12  (
    .i0(pnumcnt2[12]),
    .i1(\PWM2/n27 [12]),
    .sel(\PWM2/n24 ),
    .o(\PWM2/n29 [12]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux7_b13  (
    .i0(pnumcnt2[13]),
    .i1(\PWM2/n27 [13]),
    .sel(\PWM2/n24 ),
    .o(\PWM2/n29 [13]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux7_b14  (
    .i0(pnumcnt2[14]),
    .i1(\PWM2/n27 [14]),
    .sel(\PWM2/n24 ),
    .o(\PWM2/n29 [14]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux7_b15  (
    .i0(pnumcnt2[15]),
    .i1(\PWM2/n27 [15]),
    .sel(\PWM2/n24 ),
    .o(\PWM2/n29 [15]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux7_b16  (
    .i0(pnumcnt2[16]),
    .i1(\PWM2/n27 [16]),
    .sel(\PWM2/n24 ),
    .o(\PWM2/n29 [16]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux7_b17  (
    .i0(pnumcnt2[17]),
    .i1(\PWM2/n27 [17]),
    .sel(\PWM2/n24 ),
    .o(\PWM2/n29 [17]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux7_b18  (
    .i0(pnumcnt2[18]),
    .i1(\PWM2/n27 [18]),
    .sel(\PWM2/n24 ),
    .o(\PWM2/n29 [18]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux7_b19  (
    .i0(pnumcnt2[19]),
    .i1(\PWM2/n27 [19]),
    .sel(\PWM2/n24 ),
    .o(\PWM2/n29 [19]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux7_b2  (
    .i0(pnumcnt2[2]),
    .i1(\PWM2/n27 [2]),
    .sel(\PWM2/n24 ),
    .o(\PWM2/n29 [2]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux7_b20  (
    .i0(pnumcnt2[20]),
    .i1(\PWM2/n27 [20]),
    .sel(\PWM2/n24 ),
    .o(\PWM2/n29 [20]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux7_b21  (
    .i0(pnumcnt2[21]),
    .i1(\PWM2/n27 [21]),
    .sel(\PWM2/n24 ),
    .o(\PWM2/n29 [21]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux7_b22  (
    .i0(pnumcnt2[22]),
    .i1(\PWM2/n27 [22]),
    .sel(\PWM2/n24 ),
    .o(\PWM2/n29 [22]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux7_b23  (
    .i0(pnumcnt2[23]),
    .i1(\PWM2/n27 [23]),
    .sel(\PWM2/n24 ),
    .o(\PWM2/n29 [23]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux7_b3  (
    .i0(pnumcnt2[3]),
    .i1(\PWM2/n27 [3]),
    .sel(\PWM2/n24 ),
    .o(\PWM2/n29 [3]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux7_b4  (
    .i0(pnumcnt2[4]),
    .i1(\PWM2/n27 [4]),
    .sel(\PWM2/n24 ),
    .o(\PWM2/n29 [4]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux7_b5  (
    .i0(pnumcnt2[5]),
    .i1(\PWM2/n27 [5]),
    .sel(\PWM2/n24 ),
    .o(\PWM2/n29 [5]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux7_b6  (
    .i0(pnumcnt2[6]),
    .i1(\PWM2/n27 [6]),
    .sel(\PWM2/n24 ),
    .o(\PWM2/n29 [6]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux7_b7  (
    .i0(pnumcnt2[7]),
    .i1(\PWM2/n27 [7]),
    .sel(\PWM2/n24 ),
    .o(\PWM2/n29 [7]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux7_b8  (
    .i0(pnumcnt2[8]),
    .i1(\PWM2/n27 [8]),
    .sel(\PWM2/n24 ),
    .o(\PWM2/n29 [8]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux7_b9  (
    .i0(pnumcnt2[9]),
    .i1(\PWM2/n27 [9]),
    .sel(\PWM2/n24 ),
    .o(\PWM2/n29 [9]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux8_b0  (
    .i0(\PWM2/n29 [0]),
    .i1(\PWM2/pnumr [0]),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n31 [0]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux8_b1  (
    .i0(\PWM2/n29 [1]),
    .i1(\PWM2/pnumr [1]),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n31 [1]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux8_b10  (
    .i0(\PWM2/n29 [10]),
    .i1(\PWM2/pnumr [10]),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n31 [10]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux8_b11  (
    .i0(\PWM2/n29 [11]),
    .i1(\PWM2/pnumr [11]),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n31 [11]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux8_b12  (
    .i0(\PWM2/n29 [12]),
    .i1(\PWM2/pnumr [12]),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n31 [12]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux8_b13  (
    .i0(\PWM2/n29 [13]),
    .i1(\PWM2/pnumr [13]),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n31 [13]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux8_b14  (
    .i0(\PWM2/n29 [14]),
    .i1(\PWM2/pnumr [14]),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n31 [14]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux8_b15  (
    .i0(\PWM2/n29 [15]),
    .i1(\PWM2/pnumr [15]),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n31 [15]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux8_b16  (
    .i0(\PWM2/n29 [16]),
    .i1(\PWM2/pnumr [16]),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n31 [16]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux8_b17  (
    .i0(\PWM2/n29 [17]),
    .i1(\PWM2/pnumr [17]),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n31 [17]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux8_b18  (
    .i0(\PWM2/n29 [18]),
    .i1(\PWM2/pnumr [18]),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n31 [18]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux8_b19  (
    .i0(\PWM2/n29 [19]),
    .i1(\PWM2/pnumr [19]),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n31 [19]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux8_b2  (
    .i0(\PWM2/n29 [2]),
    .i1(\PWM2/pnumr [2]),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n31 [2]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux8_b20  (
    .i0(\PWM2/n29 [20]),
    .i1(\PWM2/pnumr [20]),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n31 [20]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux8_b21  (
    .i0(\PWM2/n29 [21]),
    .i1(\PWM2/pnumr [21]),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n31 [21]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux8_b22  (
    .i0(\PWM2/n29 [22]),
    .i1(\PWM2/pnumr [22]),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n31 [22]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux8_b23  (
    .i0(\PWM2/n29 [23]),
    .i1(\PWM2/pnumr [23]),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n31 [23]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux8_b3  (
    .i0(\PWM2/n29 [3]),
    .i1(\PWM2/pnumr [3]),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n31 [3]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux8_b4  (
    .i0(\PWM2/n29 [4]),
    .i1(\PWM2/pnumr [4]),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n31 [4]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux8_b5  (
    .i0(\PWM2/n29 [5]),
    .i1(\PWM2/pnumr [5]),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n31 [5]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux8_b6  (
    .i0(\PWM2/n29 [6]),
    .i1(\PWM2/pnumr [6]),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n31 [6]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux8_b7  (
    .i0(\PWM2/n29 [7]),
    .i1(\PWM2/pnumr [7]),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n31 [7]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux8_b8  (
    .i0(\PWM2/n29 [8]),
    .i1(\PWM2/pnumr [8]),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n31 [8]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM2/mux8_b9  (
    .i0(\PWM2/n29 [9]),
    .i1(\PWM2/pnumr [9]),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n31 [9]));  // src/OnePWM.v(57)
  not \PWM2/n17_inv  (\PWM2/n17_neg , \PWM2/n17 );
  not \PWM2/n25_inv  (\PWM2/n25_neg , \PWM2/n25 );
  not \PWM2/n4_inv  (\PWM2/n4_neg , \PWM2/n4 );
  not \PWM2/n6_inv  (\PWM2/n6_neg , \PWM2/n6 );
  ne_w24 \PWM2/neq0  (
    .i0(pnumcnt2),
    .i1(24'b000000000000000000000000),
    .o(\PWM2/n25 ));  // src/OnePWM.v(55)
  reg_sr_ss_w1 \PWM2/pwm_reg  (
    .clk(clk100m),
    .d(pwm[2]),
    .en(1'b1),
    .reset(~\PWM2/u14_sel_is_1_o ),
    .set(\PWM2/n18 ),
    .q(\PWM2/pwm_keep ));  // src/OnePWM.v(45)
  reg_sr_as_w1 \PWM2/reg0_b0  (
    .clk(clk100m),
    .d(\PWM2/n13 [0]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [0]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b1  (
    .clk(clk100m),
    .d(\PWM2/n13 [1]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [1]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b10  (
    .clk(clk100m),
    .d(\PWM2/n13 [10]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [10]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b11  (
    .clk(clk100m),
    .d(\PWM2/n13 [11]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [11]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b12  (
    .clk(clk100m),
    .d(\PWM2/n13 [12]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [12]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b13  (
    .clk(clk100m),
    .d(\PWM2/n13 [13]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [13]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b14  (
    .clk(clk100m),
    .d(\PWM2/n13 [14]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [14]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b15  (
    .clk(clk100m),
    .d(\PWM2/n13 [15]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [15]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b16  (
    .clk(clk100m),
    .d(\PWM2/n13 [16]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [16]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b17  (
    .clk(clk100m),
    .d(\PWM2/n13 [17]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [17]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b18  (
    .clk(clk100m),
    .d(\PWM2/n13 [18]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [18]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b19  (
    .clk(clk100m),
    .d(\PWM2/n13 [19]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [19]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b2  (
    .clk(clk100m),
    .d(\PWM2/n13 [2]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [2]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b20  (
    .clk(clk100m),
    .d(\PWM2/n13 [20]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [20]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b21  (
    .clk(clk100m),
    .d(\PWM2/n13 [21]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [21]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b22  (
    .clk(clk100m),
    .d(\PWM2/n13 [22]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [22]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b23  (
    .clk(clk100m),
    .d(\PWM2/n13 [23]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [23]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b24  (
    .clk(clk100m),
    .d(\PWM2/n13 [24]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [24]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b25  (
    .clk(clk100m),
    .d(\PWM2/n13 [25]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [25]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b26  (
    .clk(clk100m),
    .d(\PWM2/n13 [26]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [26]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b3  (
    .clk(clk100m),
    .d(\PWM2/n13 [3]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [3]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b4  (
    .clk(clk100m),
    .d(\PWM2/n13 [4]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [4]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b5  (
    .clk(clk100m),
    .d(\PWM2/n13 [5]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [5]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b6  (
    .clk(clk100m),
    .d(\PWM2/n13 [6]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [6]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b7  (
    .clk(clk100m),
    .d(\PWM2/n13 [7]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [7]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b8  (
    .clk(clk100m),
    .d(\PWM2/n13 [8]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [8]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM2/reg0_b9  (
    .clk(clk100m),
    .d(\PWM2/n13 [9]),
    .en(1'b1),
    .reset(~\PWM2/n11 ),
    .set(1'b0),
    .q(\PWM2/FreCnt [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b0  (
    .clk(clk100m),
    .d(freq2[0]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [0]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b1  (
    .clk(clk100m),
    .d(freq2[1]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [1]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b10  (
    .clk(clk100m),
    .d(freq2[10]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [10]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b11  (
    .clk(clk100m),
    .d(freq2[11]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [11]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b12  (
    .clk(clk100m),
    .d(freq2[12]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [12]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b13  (
    .clk(clk100m),
    .d(freq2[13]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [13]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b14  (
    .clk(clk100m),
    .d(freq2[14]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [14]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b15  (
    .clk(clk100m),
    .d(freq2[15]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [15]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b16  (
    .clk(clk100m),
    .d(freq2[16]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [16]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b17  (
    .clk(clk100m),
    .d(freq2[17]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [17]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b18  (
    .clk(clk100m),
    .d(freq2[18]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [18]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b19  (
    .clk(clk100m),
    .d(freq2[19]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [19]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b2  (
    .clk(clk100m),
    .d(freq2[2]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [2]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b20  (
    .clk(clk100m),
    .d(freq2[20]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [20]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b21  (
    .clk(clk100m),
    .d(freq2[21]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [21]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b22  (
    .clk(clk100m),
    .d(freq2[22]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [22]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b23  (
    .clk(clk100m),
    .d(freq2[23]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [23]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b24  (
    .clk(clk100m),
    .d(freq2[24]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [24]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b25  (
    .clk(clk100m),
    .d(freq2[25]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [25]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b26  (
    .clk(clk100m),
    .d(freq2[26]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [26]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b3  (
    .clk(clk100m),
    .d(freq2[3]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [3]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b4  (
    .clk(clk100m),
    .d(freq2[4]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [4]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b5  (
    .clk(clk100m),
    .d(freq2[5]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [5]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b6  (
    .clk(clk100m),
    .d(freq2[6]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [6]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b7  (
    .clk(clk100m),
    .d(freq2[7]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [7]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b8  (
    .clk(clk100m),
    .d(freq2[8]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [8]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg1_b9  (
    .clk(clk100m),
    .d(freq2[9]),
    .en(\PWM2/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/FreCntr [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM2/reg2_b0  (
    .clk(clk100m),
    .d(\PWM2/n23 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[0]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b1  (
    .clk(clk100m),
    .d(\PWM2/n23 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[1]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b10  (
    .clk(clk100m),
    .d(\PWM2/n23 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[10]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b11  (
    .clk(clk100m),
    .d(\PWM2/n23 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[11]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b12  (
    .clk(clk100m),
    .d(\PWM2/n23 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[12]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b13  (
    .clk(clk100m),
    .d(\PWM2/n23 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[13]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b14  (
    .clk(clk100m),
    .d(\PWM2/n23 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[14]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b15  (
    .clk(clk100m),
    .d(\PWM2/n23 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[15]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b16  (
    .clk(clk100m),
    .d(\PWM2/n23 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[16]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b17  (
    .clk(clk100m),
    .d(\PWM2/n23 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[17]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b18  (
    .clk(clk100m),
    .d(\PWM2/n23 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[18]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b19  (
    .clk(clk100m),
    .d(\PWM2/n23 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[19]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b2  (
    .clk(clk100m),
    .d(\PWM2/n23 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[2]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b20  (
    .clk(clk100m),
    .d(\PWM2/n23 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[20]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b21  (
    .clk(clk100m),
    .d(\PWM2/n23 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[21]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b22  (
    .clk(clk100m),
    .d(\PWM2/n23 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[22]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b23  (
    .clk(clk100m),
    .d(\PWM2/n23 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[23]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b24  (
    .clk(clk100m),
    .d(\PWM2/n23 [24]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[24]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b25  (
    .clk(clk100m),
    .d(\PWM2/n23 [25]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[25]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b26  (
    .clk(clk100m),
    .d(\PWM2/n23 [26]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[26]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b27  (
    .clk(clk100m),
    .d(\PWM2/n23 [27]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[27]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b28  (
    .clk(clk100m),
    .d(\PWM2/n23 [28]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[28]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b29  (
    .clk(clk100m),
    .d(\PWM2/n23 [29]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[29]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b3  (
    .clk(clk100m),
    .d(\PWM2/n23 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[3]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b30  (
    .clk(clk100m),
    .d(\PWM2/n23 [30]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[30]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b31  (
    .clk(clk100m),
    .d(\PWM2/n23 [31]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[31]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b4  (
    .clk(clk100m),
    .d(\PWM2/n23 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[4]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b5  (
    .clk(clk100m),
    .d(\PWM2/n23 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[5]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b6  (
    .clk(clk100m),
    .d(\PWM2/n23 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[6]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b7  (
    .clk(clk100m),
    .d(\PWM2/n23 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[7]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b8  (
    .clk(clk100m),
    .d(\PWM2/n23 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[8]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg2_b9  (
    .clk(clk100m),
    .d(\PWM2/n23 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/pnumr[9]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM2/reg3_b0  (
    .clk(clk100m),
    .d(\PWM2/n31 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[0]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b1  (
    .clk(clk100m),
    .d(\PWM2/n31 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[1]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b10  (
    .clk(clk100m),
    .d(\PWM2/n31 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[10]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b11  (
    .clk(clk100m),
    .d(\PWM2/n31 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[11]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b12  (
    .clk(clk100m),
    .d(\PWM2/n31 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[12]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b13  (
    .clk(clk100m),
    .d(\PWM2/n31 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[13]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b14  (
    .clk(clk100m),
    .d(\PWM2/n31 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[14]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b15  (
    .clk(clk100m),
    .d(\PWM2/n31 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[15]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b16  (
    .clk(clk100m),
    .d(\PWM2/n31 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[16]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b17  (
    .clk(clk100m),
    .d(\PWM2/n31 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[17]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b18  (
    .clk(clk100m),
    .d(\PWM2/n31 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[18]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b19  (
    .clk(clk100m),
    .d(\PWM2/n31 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[19]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b2  (
    .clk(clk100m),
    .d(\PWM2/n31 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[2]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b20  (
    .clk(clk100m),
    .d(\PWM2/n31 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[20]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b21  (
    .clk(clk100m),
    .d(\PWM2/n31 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[21]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b22  (
    .clk(clk100m),
    .d(\PWM2/n31 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[22]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b23  (
    .clk(clk100m),
    .d(\PWM2/n31 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[23]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b3  (
    .clk(clk100m),
    .d(\PWM2/n31 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[3]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b4  (
    .clk(clk100m),
    .d(\PWM2/n31 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[4]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b5  (
    .clk(clk100m),
    .d(\PWM2/n31 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[5]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b6  (
    .clk(clk100m),
    .d(\PWM2/n31 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[6]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b7  (
    .clk(clk100m),
    .d(\PWM2/n31 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[7]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b8  (
    .clk(clk100m),
    .d(\PWM2/n31 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[8]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM2/reg3_b9  (
    .clk(clk100m),
    .d(\PWM2/n31 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM2/RemaTxNum[9]_keep ));  // src/OnePWM.v(58)
  reg_ar_ss_w1 \PWM2/stopreq_reg  (
    .clk(clk100m),
    .d(\PWM2/n1 ),
    .en(1'b1),
    .reset(1'b0),
    .set(pwm_start_stop[2]),
    .q(\PWM2/stopreq_keep ));  // src/OnePWM.v(15)
  add_pu27_mu27_o27 \PWM2/sub0  (
    .i0(\PWM2/FreCnt ),
    .i1(27'b000000000000000000000000001),
    .o(\PWM2/n12 [26:0]));  // src/OnePWM.v(32)
  add_pu24_mu24_o24 \PWM2/sub1  (
    .i0(pnumcnt2),
    .i1(24'b000000000000000000000001),
    .o(\PWM2/n26 [23:0]));  // src/OnePWM.v(55)
  AL_MUX \PWM2/u10  (
    .i0(1'b0),
    .i1(\PWM2/n9 ),
    .sel(n13),
    .o(\PWM2/n10 ));  // src/OnePWM.v(26)
  or \PWM2/u11  (\PWM2/n11 , pwm_state_read[2], pwm_start_stop[18]);  // src/OnePWM.v(30)
  and \PWM2/u14_sel_is_1  (\PWM2/u14_sel_is_1_o , pwm_state_read[2], \PWM2/n17_neg );
  and \PWM2/u15  (\PWM2/n24 , \PWM2/n0 , pwm_state_read[2]);  // src/OnePWM.v(54)
  and \PWM2/u17_sel_is_1  (\PWM2/u17_sel_is_1_o , \PWM2/n24 , \PWM2/n25_neg );
  not \PWM2/u17_sel_is_1_o_inv  (\PWM2/u17_sel_is_1_o_neg , \PWM2/u17_sel_is_1_o );
  AL_MUX \PWM2/u18  (
    .i0(\PWM2/pnumr [31]),
    .i1(dir[2]),
    .sel(\PWM2/u18_sel_is_0_o ),
    .o(\PWM2/n32 ));
  and \PWM2/u18_sel_is_0  (\PWM2/u18_sel_is_0_o , \pwm_start_stop[18]_neg , \PWM2/u17_sel_is_1_o_neg );
  AL_MUX \PWM2/u2  (
    .i0(\PWM2/stopreq ),
    .i1(1'b0),
    .sel(\PWM2/n0 ),
    .o(\PWM2/n1 ));  // src/OnePWM.v(15)
  and \PWM2/u5  (\PWM2/n4 , \PWM2/stopreq , \PWM2/n0 );  // src/OnePWM.v(23)
  and \PWM2/u6  (\PWM2/n6 , \PWM2/n5 , \PWM2/n0 );  // src/OnePWM.v(25)
  AL_MUX \PWM2/u8  (
    .i0(1'b0),
    .i1(pwm_state_read[2]),
    .sel(\PWM2/u8_sel_is_0_o ),
    .o(\PWM2/n8 ));
  and \PWM2/u8_sel_is_0  (\PWM2/u8_sel_is_0_o , \PWM2/n4_neg , \PWM2/n6_neg );
  AL_MUX \PWM2/u9  (
    .i0(\PWM2/n8 ),
    .i1(1'b1),
    .sel(pwm_start_stop[18]),
    .o(\PWM2/n9 ));  // src/OnePWM.v(26)
  reg_ar_as_w1 \PWM3/State_reg  (
    .clk(clk100m),
    .d(\PWM3/n10 ),
    .en(1'b1),
    .reset(~rstn),
    .set(1'b0),
    .q(pwm_state_read[3]));  // src/OnePWM.v(26)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[0]  (
    .i(\PWM3/RemaTxNum[0]_keep ),
    .o(pnumcnt3[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[10]  (
    .i(\PWM3/RemaTxNum[10]_keep ),
    .o(pnumcnt3[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[11]  (
    .i(\PWM3/RemaTxNum[11]_keep ),
    .o(pnumcnt3[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[12]  (
    .i(\PWM3/RemaTxNum[12]_keep ),
    .o(pnumcnt3[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[13]  (
    .i(\PWM3/RemaTxNum[13]_keep ),
    .o(pnumcnt3[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[14]  (
    .i(\PWM3/RemaTxNum[14]_keep ),
    .o(pnumcnt3[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[15]  (
    .i(\PWM3/RemaTxNum[15]_keep ),
    .o(pnumcnt3[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[16]  (
    .i(\PWM3/RemaTxNum[16]_keep ),
    .o(pnumcnt3[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[17]  (
    .i(\PWM3/RemaTxNum[17]_keep ),
    .o(pnumcnt3[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[18]  (
    .i(\PWM3/RemaTxNum[18]_keep ),
    .o(pnumcnt3[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[19]  (
    .i(\PWM3/RemaTxNum[19]_keep ),
    .o(pnumcnt3[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[1]  (
    .i(\PWM3/RemaTxNum[1]_keep ),
    .o(pnumcnt3[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[20]  (
    .i(\PWM3/RemaTxNum[20]_keep ),
    .o(pnumcnt3[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[21]  (
    .i(\PWM3/RemaTxNum[21]_keep ),
    .o(pnumcnt3[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[22]  (
    .i(\PWM3/RemaTxNum[22]_keep ),
    .o(pnumcnt3[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[23]  (
    .i(\PWM3/RemaTxNum[23]_keep ),
    .o(pnumcnt3[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[2]  (
    .i(\PWM3/RemaTxNum[2]_keep ),
    .o(pnumcnt3[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[3]  (
    .i(\PWM3/RemaTxNum[3]_keep ),
    .o(pnumcnt3[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[4]  (
    .i(\PWM3/RemaTxNum[4]_keep ),
    .o(pnumcnt3[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[5]  (
    .i(\PWM3/RemaTxNum[5]_keep ),
    .o(pnumcnt3[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[6]  (
    .i(\PWM3/RemaTxNum[6]_keep ),
    .o(pnumcnt3[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[7]  (
    .i(\PWM3/RemaTxNum[7]_keep ),
    .o(pnumcnt3[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[8]  (
    .i(\PWM3/RemaTxNum[8]_keep ),
    .o(pnumcnt3[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_RemaTxNum[9]  (
    .i(\PWM3/RemaTxNum[9]_keep ),
    .o(pnumcnt3[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_dir  (
    .i(\PWM3/dir_keep ),
    .o(dir[3]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[0]  (
    .i(\PWM3/pnumr[0]_keep ),
    .o(\PWM3/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[10]  (
    .i(\PWM3/pnumr[10]_keep ),
    .o(\PWM3/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[11]  (
    .i(\PWM3/pnumr[11]_keep ),
    .o(\PWM3/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[12]  (
    .i(\PWM3/pnumr[12]_keep ),
    .o(\PWM3/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[13]  (
    .i(\PWM3/pnumr[13]_keep ),
    .o(\PWM3/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[14]  (
    .i(\PWM3/pnumr[14]_keep ),
    .o(\PWM3/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[15]  (
    .i(\PWM3/pnumr[15]_keep ),
    .o(\PWM3/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[16]  (
    .i(\PWM3/pnumr[16]_keep ),
    .o(\PWM3/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[17]  (
    .i(\PWM3/pnumr[17]_keep ),
    .o(\PWM3/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[18]  (
    .i(\PWM3/pnumr[18]_keep ),
    .o(\PWM3/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[19]  (
    .i(\PWM3/pnumr[19]_keep ),
    .o(\PWM3/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[1]  (
    .i(\PWM3/pnumr[1]_keep ),
    .o(\PWM3/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[20]  (
    .i(\PWM3/pnumr[20]_keep ),
    .o(\PWM3/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[21]  (
    .i(\PWM3/pnumr[21]_keep ),
    .o(\PWM3/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[22]  (
    .i(\PWM3/pnumr[22]_keep ),
    .o(\PWM3/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[23]  (
    .i(\PWM3/pnumr[23]_keep ),
    .o(\PWM3/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[24]  (
    .i(\PWM3/pnumr[24]_keep ),
    .o(\PWM3/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[25]  (
    .i(\PWM3/pnumr[25]_keep ),
    .o(\PWM3/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[26]  (
    .i(\PWM3/pnumr[26]_keep ),
    .o(\PWM3/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[27]  (
    .i(\PWM3/pnumr[27]_keep ),
    .o(\PWM3/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[28]  (
    .i(\PWM3/pnumr[28]_keep ),
    .o(\PWM3/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[29]  (
    .i(\PWM3/pnumr[29]_keep ),
    .o(\PWM3/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[2]  (
    .i(\PWM3/pnumr[2]_keep ),
    .o(\PWM3/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[30]  (
    .i(\PWM3/pnumr[30]_keep ),
    .o(\PWM3/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[31]  (
    .i(\PWM3/pnumr[31]_keep ),
    .o(\PWM3/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[3]  (
    .i(\PWM3/pnumr[3]_keep ),
    .o(\PWM3/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[4]  (
    .i(\PWM3/pnumr[4]_keep ),
    .o(\PWM3/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[5]  (
    .i(\PWM3/pnumr[5]_keep ),
    .o(\PWM3/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[6]  (
    .i(\PWM3/pnumr[6]_keep ),
    .o(\PWM3/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[7]  (
    .i(\PWM3/pnumr[7]_keep ),
    .o(\PWM3/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[8]  (
    .i(\PWM3/pnumr[8]_keep ),
    .o(\PWM3/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pnumr[9]  (
    .i(\PWM3/pnumr[9]_keep ),
    .o(\PWM3/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_pwm  (
    .i(\PWM3/pwm_keep ),
    .o(pwm[3]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM3/_bufkeep_stopreq  (
    .i(\PWM3/stopreq_keep ),
    .o(\PWM3/stopreq ));  // src/OnePWM.v(14)
  reg_ar_as_w1 \PWM3/dir_reg  (
    .clk(clk100m),
    .d(\PWM3/n32 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/dir_keep ));  // src/OnePWM.v(58)
  eq_w27 \PWM3/eq0  (
    .i0(\PWM3/FreCnt ),
    .i1(27'b000000000000000000000000000),
    .o(\PWM3/n0 ));  // src/OnePWM.v(15)
  eq_w24 \PWM3/eq1  (
    .i0(pnumcnt3),
    .i1(24'b000000000000000000000001),
    .o(\PWM3/n5 ));  // src/OnePWM.v(25)
  eq_w27 \PWM3/eq2  (
    .i0(\PWM3/FreCnt ),
    .i1({1'b0,\PWM3/FreCntr [26:1]}),
    .o(\PWM3/n17 ));  // src/OnePWM.v(41)
  eq_w27 \PWM3/eq3  (
    .i0(\PWM3/FreCnt ),
    .i1(\PWM3/FreCntr ),
    .o(\PWM3/n18 ));  // src/OnePWM.v(43)
  binary_mux_s1_w1 \PWM3/mux0_b0  (
    .i0(\PWM3/n12 [0]),
    .i1(freq3[0]),
    .sel(\PWM3/n0 ),
    .o(\PWM3/n13 [0]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM3/mux0_b1  (
    .i0(\PWM3/n12 [1]),
    .i1(freq3[1]),
    .sel(\PWM3/n0 ),
    .o(\PWM3/n13 [1]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM3/mux0_b10  (
    .i0(\PWM3/n12 [10]),
    .i1(freq3[10]),
    .sel(\PWM3/n0 ),
    .o(\PWM3/n13 [10]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM3/mux0_b11  (
    .i0(\PWM3/n12 [11]),
    .i1(freq3[11]),
    .sel(\PWM3/n0 ),
    .o(\PWM3/n13 [11]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM3/mux0_b12  (
    .i0(\PWM3/n12 [12]),
    .i1(freq3[12]),
    .sel(\PWM3/n0 ),
    .o(\PWM3/n13 [12]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM3/mux0_b13  (
    .i0(\PWM3/n12 [13]),
    .i1(freq3[13]),
    .sel(\PWM3/n0 ),
    .o(\PWM3/n13 [13]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM3/mux0_b14  (
    .i0(\PWM3/n12 [14]),
    .i1(freq3[14]),
    .sel(\PWM3/n0 ),
    .o(\PWM3/n13 [14]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM3/mux0_b15  (
    .i0(\PWM3/n12 [15]),
    .i1(freq3[15]),
    .sel(\PWM3/n0 ),
    .o(\PWM3/n13 [15]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM3/mux0_b16  (
    .i0(\PWM3/n12 [16]),
    .i1(freq3[16]),
    .sel(\PWM3/n0 ),
    .o(\PWM3/n13 [16]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM3/mux0_b17  (
    .i0(\PWM3/n12 [17]),
    .i1(freq3[17]),
    .sel(\PWM3/n0 ),
    .o(\PWM3/n13 [17]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM3/mux0_b18  (
    .i0(\PWM3/n12 [18]),
    .i1(freq3[18]),
    .sel(\PWM3/n0 ),
    .o(\PWM3/n13 [18]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM3/mux0_b19  (
    .i0(\PWM3/n12 [19]),
    .i1(freq3[19]),
    .sel(\PWM3/n0 ),
    .o(\PWM3/n13 [19]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM3/mux0_b2  (
    .i0(\PWM3/n12 [2]),
    .i1(freq3[2]),
    .sel(\PWM3/n0 ),
    .o(\PWM3/n13 [2]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM3/mux0_b20  (
    .i0(\PWM3/n12 [20]),
    .i1(freq3[20]),
    .sel(\PWM3/n0 ),
    .o(\PWM3/n13 [20]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM3/mux0_b21  (
    .i0(\PWM3/n12 [21]),
    .i1(freq3[21]),
    .sel(\PWM3/n0 ),
    .o(\PWM3/n13 [21]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM3/mux0_b22  (
    .i0(\PWM3/n12 [22]),
    .i1(freq3[22]),
    .sel(\PWM3/n0 ),
    .o(\PWM3/n13 [22]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM3/mux0_b23  (
    .i0(\PWM3/n12 [23]),
    .i1(freq3[23]),
    .sel(\PWM3/n0 ),
    .o(\PWM3/n13 [23]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM3/mux0_b24  (
    .i0(\PWM3/n12 [24]),
    .i1(freq3[24]),
    .sel(\PWM3/n0 ),
    .o(\PWM3/n13 [24]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM3/mux0_b25  (
    .i0(\PWM3/n12 [25]),
    .i1(freq3[25]),
    .sel(\PWM3/n0 ),
    .o(\PWM3/n13 [25]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM3/mux0_b26  (
    .i0(\PWM3/n12 [26]),
    .i1(freq3[26]),
    .sel(\PWM3/n0 ),
    .o(\PWM3/n13 [26]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM3/mux0_b3  (
    .i0(\PWM3/n12 [3]),
    .i1(freq3[3]),
    .sel(\PWM3/n0 ),
    .o(\PWM3/n13 [3]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM3/mux0_b4  (
    .i0(\PWM3/n12 [4]),
    .i1(freq3[4]),
    .sel(\PWM3/n0 ),
    .o(\PWM3/n13 [4]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM3/mux0_b5  (
    .i0(\PWM3/n12 [5]),
    .i1(freq3[5]),
    .sel(\PWM3/n0 ),
    .o(\PWM3/n13 [5]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM3/mux0_b6  (
    .i0(\PWM3/n12 [6]),
    .i1(freq3[6]),
    .sel(\PWM3/n0 ),
    .o(\PWM3/n13 [6]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM3/mux0_b7  (
    .i0(\PWM3/n12 [7]),
    .i1(freq3[7]),
    .sel(\PWM3/n0 ),
    .o(\PWM3/n13 [7]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM3/mux0_b8  (
    .i0(\PWM3/n12 [8]),
    .i1(freq3[8]),
    .sel(\PWM3/n0 ),
    .o(\PWM3/n13 [8]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM3/mux0_b9  (
    .i0(\PWM3/n12 [9]),
    .i1(freq3[9]),
    .sel(\PWM3/n0 ),
    .o(\PWM3/n13 [9]));  // src/OnePWM.v(32)
  and \PWM3/mux3_b0_sel_is_3  (\PWM3/mux3_b0_sel_is_3_o , \PWM3/n11 , \PWM3/n0 );
  binary_mux_s1_w1 \PWM3/mux4_b0  (
    .i0(\PWM3/pnumr [0]),
    .i1(1'b0),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n22 [0]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux4_b1  (
    .i0(\PWM3/pnumr [1]),
    .i1(1'b0),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n22 [1]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux4_b10  (
    .i0(\PWM3/pnumr [10]),
    .i1(1'b0),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n22 [10]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux4_b11  (
    .i0(\PWM3/pnumr [11]),
    .i1(1'b0),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n22 [11]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux4_b12  (
    .i0(\PWM3/pnumr [12]),
    .i1(1'b0),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n22 [12]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux4_b13  (
    .i0(\PWM3/pnumr [13]),
    .i1(1'b0),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n22 [13]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux4_b14  (
    .i0(\PWM3/pnumr [14]),
    .i1(1'b0),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n22 [14]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux4_b15  (
    .i0(\PWM3/pnumr [15]),
    .i1(1'b0),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n22 [15]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux4_b16  (
    .i0(\PWM3/pnumr [16]),
    .i1(1'b0),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n22 [16]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux4_b17  (
    .i0(\PWM3/pnumr [17]),
    .i1(1'b0),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n22 [17]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux4_b18  (
    .i0(\PWM3/pnumr [18]),
    .i1(1'b0),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n22 [18]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux4_b19  (
    .i0(\PWM3/pnumr [19]),
    .i1(1'b0),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n22 [19]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux4_b2  (
    .i0(\PWM3/pnumr [2]),
    .i1(1'b0),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n22 [2]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux4_b20  (
    .i0(\PWM3/pnumr [20]),
    .i1(1'b0),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n22 [20]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux4_b21  (
    .i0(\PWM3/pnumr [21]),
    .i1(1'b0),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n22 [21]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux4_b22  (
    .i0(\PWM3/pnumr [22]),
    .i1(1'b0),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n22 [22]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux4_b23  (
    .i0(\PWM3/pnumr [23]),
    .i1(1'b0),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n22 [23]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux4_b24  (
    .i0(\PWM3/pnumr [24]),
    .i1(1'b0),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n22 [24]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux4_b25  (
    .i0(\PWM3/pnumr [25]),
    .i1(1'b0),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n22 [25]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux4_b26  (
    .i0(\PWM3/pnumr [26]),
    .i1(1'b0),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n22 [26]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux4_b27  (
    .i0(\PWM3/pnumr [27]),
    .i1(1'b0),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n22 [27]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux4_b28  (
    .i0(\PWM3/pnumr [28]),
    .i1(1'b0),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n22 [28]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux4_b29  (
    .i0(\PWM3/pnumr [29]),
    .i1(1'b0),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n22 [29]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux4_b3  (
    .i0(\PWM3/pnumr [3]),
    .i1(1'b0),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n22 [3]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux4_b30  (
    .i0(\PWM3/pnumr [30]),
    .i1(1'b0),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n22 [30]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux4_b31  (
    .i0(\PWM3/pnumr [31]),
    .i1(1'b0),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n22 [31]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux4_b4  (
    .i0(\PWM3/pnumr [4]),
    .i1(1'b0),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n22 [4]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux4_b5  (
    .i0(\PWM3/pnumr [5]),
    .i1(1'b0),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n22 [5]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux4_b6  (
    .i0(\PWM3/pnumr [6]),
    .i1(1'b0),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n22 [6]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux4_b7  (
    .i0(\PWM3/pnumr [7]),
    .i1(1'b0),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n22 [7]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux4_b8  (
    .i0(\PWM3/pnumr [8]),
    .i1(1'b0),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n22 [8]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux4_b9  (
    .i0(\PWM3/pnumr [9]),
    .i1(1'b0),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n22 [9]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux5_b0  (
    .i0(\PWM3/n22 [0]),
    .i1(pnum3[0]),
    .sel(pnum3[32]),
    .o(\PWM3/n23 [0]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux5_b1  (
    .i0(\PWM3/n22 [1]),
    .i1(pnum3[1]),
    .sel(pnum3[32]),
    .o(\PWM3/n23 [1]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux5_b10  (
    .i0(\PWM3/n22 [10]),
    .i1(pnum3[10]),
    .sel(pnum3[32]),
    .o(\PWM3/n23 [10]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux5_b11  (
    .i0(\PWM3/n22 [11]),
    .i1(pnum3[11]),
    .sel(pnum3[32]),
    .o(\PWM3/n23 [11]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux5_b12  (
    .i0(\PWM3/n22 [12]),
    .i1(pnum3[12]),
    .sel(pnum3[32]),
    .o(\PWM3/n23 [12]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux5_b13  (
    .i0(\PWM3/n22 [13]),
    .i1(pnum3[13]),
    .sel(pnum3[32]),
    .o(\PWM3/n23 [13]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux5_b14  (
    .i0(\PWM3/n22 [14]),
    .i1(pnum3[14]),
    .sel(pnum3[32]),
    .o(\PWM3/n23 [14]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux5_b15  (
    .i0(\PWM3/n22 [15]),
    .i1(pnum3[15]),
    .sel(pnum3[32]),
    .o(\PWM3/n23 [15]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux5_b16  (
    .i0(\PWM3/n22 [16]),
    .i1(pnum3[16]),
    .sel(pnum3[32]),
    .o(\PWM3/n23 [16]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux5_b17  (
    .i0(\PWM3/n22 [17]),
    .i1(pnum3[17]),
    .sel(pnum3[32]),
    .o(\PWM3/n23 [17]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux5_b18  (
    .i0(\PWM3/n22 [18]),
    .i1(pnum3[18]),
    .sel(pnum3[32]),
    .o(\PWM3/n23 [18]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux5_b19  (
    .i0(\PWM3/n22 [19]),
    .i1(pnum3[19]),
    .sel(pnum3[32]),
    .o(\PWM3/n23 [19]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux5_b2  (
    .i0(\PWM3/n22 [2]),
    .i1(pnum3[2]),
    .sel(pnum3[32]),
    .o(\PWM3/n23 [2]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux5_b20  (
    .i0(\PWM3/n22 [20]),
    .i1(pnum3[20]),
    .sel(pnum3[32]),
    .o(\PWM3/n23 [20]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux5_b21  (
    .i0(\PWM3/n22 [21]),
    .i1(pnum3[21]),
    .sel(pnum3[32]),
    .o(\PWM3/n23 [21]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux5_b22  (
    .i0(\PWM3/n22 [22]),
    .i1(pnum3[22]),
    .sel(pnum3[32]),
    .o(\PWM3/n23 [22]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux5_b23  (
    .i0(\PWM3/n22 [23]),
    .i1(pnum3[23]),
    .sel(pnum3[32]),
    .o(\PWM3/n23 [23]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux5_b24  (
    .i0(\PWM3/n22 [24]),
    .i1(pnum3[24]),
    .sel(pnum3[32]),
    .o(\PWM3/n23 [24]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux5_b25  (
    .i0(\PWM3/n22 [25]),
    .i1(pnum3[25]),
    .sel(pnum3[32]),
    .o(\PWM3/n23 [25]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux5_b26  (
    .i0(\PWM3/n22 [26]),
    .i1(pnum3[26]),
    .sel(pnum3[32]),
    .o(\PWM3/n23 [26]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux5_b27  (
    .i0(\PWM3/n22 [27]),
    .i1(pnum3[27]),
    .sel(pnum3[32]),
    .o(\PWM3/n23 [27]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux5_b28  (
    .i0(\PWM3/n22 [28]),
    .i1(pnum3[28]),
    .sel(pnum3[32]),
    .o(\PWM3/n23 [28]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux5_b29  (
    .i0(\PWM3/n22 [29]),
    .i1(pnum3[29]),
    .sel(pnum3[32]),
    .o(\PWM3/n23 [29]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux5_b3  (
    .i0(\PWM3/n22 [3]),
    .i1(pnum3[3]),
    .sel(pnum3[32]),
    .o(\PWM3/n23 [3]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux5_b30  (
    .i0(\PWM3/n22 [30]),
    .i1(pnum3[30]),
    .sel(pnum3[32]),
    .o(\PWM3/n23 [30]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux5_b31  (
    .i0(\PWM3/n22 [31]),
    .i1(pnum3[31]),
    .sel(pnum3[32]),
    .o(\PWM3/n23 [31]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux5_b4  (
    .i0(\PWM3/n22 [4]),
    .i1(pnum3[4]),
    .sel(pnum3[32]),
    .o(\PWM3/n23 [4]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux5_b5  (
    .i0(\PWM3/n22 [5]),
    .i1(pnum3[5]),
    .sel(pnum3[32]),
    .o(\PWM3/n23 [5]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux5_b6  (
    .i0(\PWM3/n22 [6]),
    .i1(pnum3[6]),
    .sel(pnum3[32]),
    .o(\PWM3/n23 [6]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux5_b7  (
    .i0(\PWM3/n22 [7]),
    .i1(pnum3[7]),
    .sel(pnum3[32]),
    .o(\PWM3/n23 [7]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux5_b8  (
    .i0(\PWM3/n22 [8]),
    .i1(pnum3[8]),
    .sel(pnum3[32]),
    .o(\PWM3/n23 [8]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux5_b9  (
    .i0(\PWM3/n22 [9]),
    .i1(pnum3[9]),
    .sel(pnum3[32]),
    .o(\PWM3/n23 [9]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM3/mux6_b0  (
    .i0(\PWM3/pnumr [0]),
    .i1(\PWM3/n26 [0]),
    .sel(\PWM3/n25 ),
    .o(\PWM3/n27 [0]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM3/mux6_b1  (
    .i0(\PWM3/pnumr [1]),
    .i1(\PWM3/n26 [1]),
    .sel(\PWM3/n25 ),
    .o(\PWM3/n27 [1]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM3/mux6_b10  (
    .i0(\PWM3/pnumr [10]),
    .i1(\PWM3/n26 [10]),
    .sel(\PWM3/n25 ),
    .o(\PWM3/n27 [10]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM3/mux6_b11  (
    .i0(\PWM3/pnumr [11]),
    .i1(\PWM3/n26 [11]),
    .sel(\PWM3/n25 ),
    .o(\PWM3/n27 [11]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM3/mux6_b12  (
    .i0(\PWM3/pnumr [12]),
    .i1(\PWM3/n26 [12]),
    .sel(\PWM3/n25 ),
    .o(\PWM3/n27 [12]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM3/mux6_b13  (
    .i0(\PWM3/pnumr [13]),
    .i1(\PWM3/n26 [13]),
    .sel(\PWM3/n25 ),
    .o(\PWM3/n27 [13]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM3/mux6_b14  (
    .i0(\PWM3/pnumr [14]),
    .i1(\PWM3/n26 [14]),
    .sel(\PWM3/n25 ),
    .o(\PWM3/n27 [14]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM3/mux6_b15  (
    .i0(\PWM3/pnumr [15]),
    .i1(\PWM3/n26 [15]),
    .sel(\PWM3/n25 ),
    .o(\PWM3/n27 [15]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM3/mux6_b16  (
    .i0(\PWM3/pnumr [16]),
    .i1(\PWM3/n26 [16]),
    .sel(\PWM3/n25 ),
    .o(\PWM3/n27 [16]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM3/mux6_b17  (
    .i0(\PWM3/pnumr [17]),
    .i1(\PWM3/n26 [17]),
    .sel(\PWM3/n25 ),
    .o(\PWM3/n27 [17]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM3/mux6_b18  (
    .i0(\PWM3/pnumr [18]),
    .i1(\PWM3/n26 [18]),
    .sel(\PWM3/n25 ),
    .o(\PWM3/n27 [18]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM3/mux6_b19  (
    .i0(\PWM3/pnumr [19]),
    .i1(\PWM3/n26 [19]),
    .sel(\PWM3/n25 ),
    .o(\PWM3/n27 [19]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM3/mux6_b2  (
    .i0(\PWM3/pnumr [2]),
    .i1(\PWM3/n26 [2]),
    .sel(\PWM3/n25 ),
    .o(\PWM3/n27 [2]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM3/mux6_b20  (
    .i0(\PWM3/pnumr [20]),
    .i1(\PWM3/n26 [20]),
    .sel(\PWM3/n25 ),
    .o(\PWM3/n27 [20]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM3/mux6_b21  (
    .i0(\PWM3/pnumr [21]),
    .i1(\PWM3/n26 [21]),
    .sel(\PWM3/n25 ),
    .o(\PWM3/n27 [21]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM3/mux6_b22  (
    .i0(\PWM3/pnumr [22]),
    .i1(\PWM3/n26 [22]),
    .sel(\PWM3/n25 ),
    .o(\PWM3/n27 [22]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM3/mux6_b23  (
    .i0(\PWM3/pnumr [23]),
    .i1(\PWM3/n26 [23]),
    .sel(\PWM3/n25 ),
    .o(\PWM3/n27 [23]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM3/mux6_b3  (
    .i0(\PWM3/pnumr [3]),
    .i1(\PWM3/n26 [3]),
    .sel(\PWM3/n25 ),
    .o(\PWM3/n27 [3]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM3/mux6_b4  (
    .i0(\PWM3/pnumr [4]),
    .i1(\PWM3/n26 [4]),
    .sel(\PWM3/n25 ),
    .o(\PWM3/n27 [4]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM3/mux6_b5  (
    .i0(\PWM3/pnumr [5]),
    .i1(\PWM3/n26 [5]),
    .sel(\PWM3/n25 ),
    .o(\PWM3/n27 [5]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM3/mux6_b6  (
    .i0(\PWM3/pnumr [6]),
    .i1(\PWM3/n26 [6]),
    .sel(\PWM3/n25 ),
    .o(\PWM3/n27 [6]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM3/mux6_b7  (
    .i0(\PWM3/pnumr [7]),
    .i1(\PWM3/n26 [7]),
    .sel(\PWM3/n25 ),
    .o(\PWM3/n27 [7]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM3/mux6_b8  (
    .i0(\PWM3/pnumr [8]),
    .i1(\PWM3/n26 [8]),
    .sel(\PWM3/n25 ),
    .o(\PWM3/n27 [8]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM3/mux6_b9  (
    .i0(\PWM3/pnumr [9]),
    .i1(\PWM3/n26 [9]),
    .sel(\PWM3/n25 ),
    .o(\PWM3/n27 [9]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM3/mux7_b0  (
    .i0(pnumcnt3[0]),
    .i1(\PWM3/n27 [0]),
    .sel(\PWM3/n24 ),
    .o(\PWM3/n29 [0]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux7_b1  (
    .i0(pnumcnt3[1]),
    .i1(\PWM3/n27 [1]),
    .sel(\PWM3/n24 ),
    .o(\PWM3/n29 [1]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux7_b10  (
    .i0(pnumcnt3[10]),
    .i1(\PWM3/n27 [10]),
    .sel(\PWM3/n24 ),
    .o(\PWM3/n29 [10]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux7_b11  (
    .i0(pnumcnt3[11]),
    .i1(\PWM3/n27 [11]),
    .sel(\PWM3/n24 ),
    .o(\PWM3/n29 [11]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux7_b12  (
    .i0(pnumcnt3[12]),
    .i1(\PWM3/n27 [12]),
    .sel(\PWM3/n24 ),
    .o(\PWM3/n29 [12]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux7_b13  (
    .i0(pnumcnt3[13]),
    .i1(\PWM3/n27 [13]),
    .sel(\PWM3/n24 ),
    .o(\PWM3/n29 [13]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux7_b14  (
    .i0(pnumcnt3[14]),
    .i1(\PWM3/n27 [14]),
    .sel(\PWM3/n24 ),
    .o(\PWM3/n29 [14]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux7_b15  (
    .i0(pnumcnt3[15]),
    .i1(\PWM3/n27 [15]),
    .sel(\PWM3/n24 ),
    .o(\PWM3/n29 [15]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux7_b16  (
    .i0(pnumcnt3[16]),
    .i1(\PWM3/n27 [16]),
    .sel(\PWM3/n24 ),
    .o(\PWM3/n29 [16]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux7_b17  (
    .i0(pnumcnt3[17]),
    .i1(\PWM3/n27 [17]),
    .sel(\PWM3/n24 ),
    .o(\PWM3/n29 [17]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux7_b18  (
    .i0(pnumcnt3[18]),
    .i1(\PWM3/n27 [18]),
    .sel(\PWM3/n24 ),
    .o(\PWM3/n29 [18]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux7_b19  (
    .i0(pnumcnt3[19]),
    .i1(\PWM3/n27 [19]),
    .sel(\PWM3/n24 ),
    .o(\PWM3/n29 [19]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux7_b2  (
    .i0(pnumcnt3[2]),
    .i1(\PWM3/n27 [2]),
    .sel(\PWM3/n24 ),
    .o(\PWM3/n29 [2]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux7_b20  (
    .i0(pnumcnt3[20]),
    .i1(\PWM3/n27 [20]),
    .sel(\PWM3/n24 ),
    .o(\PWM3/n29 [20]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux7_b21  (
    .i0(pnumcnt3[21]),
    .i1(\PWM3/n27 [21]),
    .sel(\PWM3/n24 ),
    .o(\PWM3/n29 [21]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux7_b22  (
    .i0(pnumcnt3[22]),
    .i1(\PWM3/n27 [22]),
    .sel(\PWM3/n24 ),
    .o(\PWM3/n29 [22]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux7_b23  (
    .i0(pnumcnt3[23]),
    .i1(\PWM3/n27 [23]),
    .sel(\PWM3/n24 ),
    .o(\PWM3/n29 [23]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux7_b3  (
    .i0(pnumcnt3[3]),
    .i1(\PWM3/n27 [3]),
    .sel(\PWM3/n24 ),
    .o(\PWM3/n29 [3]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux7_b4  (
    .i0(pnumcnt3[4]),
    .i1(\PWM3/n27 [4]),
    .sel(\PWM3/n24 ),
    .o(\PWM3/n29 [4]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux7_b5  (
    .i0(pnumcnt3[5]),
    .i1(\PWM3/n27 [5]),
    .sel(\PWM3/n24 ),
    .o(\PWM3/n29 [5]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux7_b6  (
    .i0(pnumcnt3[6]),
    .i1(\PWM3/n27 [6]),
    .sel(\PWM3/n24 ),
    .o(\PWM3/n29 [6]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux7_b7  (
    .i0(pnumcnt3[7]),
    .i1(\PWM3/n27 [7]),
    .sel(\PWM3/n24 ),
    .o(\PWM3/n29 [7]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux7_b8  (
    .i0(pnumcnt3[8]),
    .i1(\PWM3/n27 [8]),
    .sel(\PWM3/n24 ),
    .o(\PWM3/n29 [8]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux7_b9  (
    .i0(pnumcnt3[9]),
    .i1(\PWM3/n27 [9]),
    .sel(\PWM3/n24 ),
    .o(\PWM3/n29 [9]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux8_b0  (
    .i0(\PWM3/n29 [0]),
    .i1(\PWM3/pnumr [0]),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n31 [0]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux8_b1  (
    .i0(\PWM3/n29 [1]),
    .i1(\PWM3/pnumr [1]),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n31 [1]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux8_b10  (
    .i0(\PWM3/n29 [10]),
    .i1(\PWM3/pnumr [10]),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n31 [10]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux8_b11  (
    .i0(\PWM3/n29 [11]),
    .i1(\PWM3/pnumr [11]),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n31 [11]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux8_b12  (
    .i0(\PWM3/n29 [12]),
    .i1(\PWM3/pnumr [12]),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n31 [12]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux8_b13  (
    .i0(\PWM3/n29 [13]),
    .i1(\PWM3/pnumr [13]),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n31 [13]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux8_b14  (
    .i0(\PWM3/n29 [14]),
    .i1(\PWM3/pnumr [14]),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n31 [14]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux8_b15  (
    .i0(\PWM3/n29 [15]),
    .i1(\PWM3/pnumr [15]),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n31 [15]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux8_b16  (
    .i0(\PWM3/n29 [16]),
    .i1(\PWM3/pnumr [16]),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n31 [16]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux8_b17  (
    .i0(\PWM3/n29 [17]),
    .i1(\PWM3/pnumr [17]),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n31 [17]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux8_b18  (
    .i0(\PWM3/n29 [18]),
    .i1(\PWM3/pnumr [18]),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n31 [18]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux8_b19  (
    .i0(\PWM3/n29 [19]),
    .i1(\PWM3/pnumr [19]),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n31 [19]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux8_b2  (
    .i0(\PWM3/n29 [2]),
    .i1(\PWM3/pnumr [2]),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n31 [2]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux8_b20  (
    .i0(\PWM3/n29 [20]),
    .i1(\PWM3/pnumr [20]),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n31 [20]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux8_b21  (
    .i0(\PWM3/n29 [21]),
    .i1(\PWM3/pnumr [21]),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n31 [21]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux8_b22  (
    .i0(\PWM3/n29 [22]),
    .i1(\PWM3/pnumr [22]),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n31 [22]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux8_b23  (
    .i0(\PWM3/n29 [23]),
    .i1(\PWM3/pnumr [23]),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n31 [23]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux8_b3  (
    .i0(\PWM3/n29 [3]),
    .i1(\PWM3/pnumr [3]),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n31 [3]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux8_b4  (
    .i0(\PWM3/n29 [4]),
    .i1(\PWM3/pnumr [4]),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n31 [4]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux8_b5  (
    .i0(\PWM3/n29 [5]),
    .i1(\PWM3/pnumr [5]),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n31 [5]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux8_b6  (
    .i0(\PWM3/n29 [6]),
    .i1(\PWM3/pnumr [6]),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n31 [6]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux8_b7  (
    .i0(\PWM3/n29 [7]),
    .i1(\PWM3/pnumr [7]),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n31 [7]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux8_b8  (
    .i0(\PWM3/n29 [8]),
    .i1(\PWM3/pnumr [8]),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n31 [8]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM3/mux8_b9  (
    .i0(\PWM3/n29 [9]),
    .i1(\PWM3/pnumr [9]),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n31 [9]));  // src/OnePWM.v(57)
  not \PWM3/n17_inv  (\PWM3/n17_neg , \PWM3/n17 );
  not \PWM3/n25_inv  (\PWM3/n25_neg , \PWM3/n25 );
  not \PWM3/n4_inv  (\PWM3/n4_neg , \PWM3/n4 );
  not \PWM3/n6_inv  (\PWM3/n6_neg , \PWM3/n6 );
  ne_w24 \PWM3/neq0  (
    .i0(pnumcnt3),
    .i1(24'b000000000000000000000000),
    .o(\PWM3/n25 ));  // src/OnePWM.v(55)
  reg_sr_ss_w1 \PWM3/pwm_reg  (
    .clk(clk100m),
    .d(pwm[3]),
    .en(1'b1),
    .reset(~\PWM3/u14_sel_is_1_o ),
    .set(\PWM3/n18 ),
    .q(\PWM3/pwm_keep ));  // src/OnePWM.v(45)
  reg_sr_as_w1 \PWM3/reg0_b0  (
    .clk(clk100m),
    .d(\PWM3/n13 [0]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [0]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b1  (
    .clk(clk100m),
    .d(\PWM3/n13 [1]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [1]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b10  (
    .clk(clk100m),
    .d(\PWM3/n13 [10]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [10]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b11  (
    .clk(clk100m),
    .d(\PWM3/n13 [11]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [11]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b12  (
    .clk(clk100m),
    .d(\PWM3/n13 [12]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [12]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b13  (
    .clk(clk100m),
    .d(\PWM3/n13 [13]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [13]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b14  (
    .clk(clk100m),
    .d(\PWM3/n13 [14]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [14]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b15  (
    .clk(clk100m),
    .d(\PWM3/n13 [15]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [15]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b16  (
    .clk(clk100m),
    .d(\PWM3/n13 [16]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [16]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b17  (
    .clk(clk100m),
    .d(\PWM3/n13 [17]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [17]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b18  (
    .clk(clk100m),
    .d(\PWM3/n13 [18]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [18]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b19  (
    .clk(clk100m),
    .d(\PWM3/n13 [19]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [19]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b2  (
    .clk(clk100m),
    .d(\PWM3/n13 [2]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [2]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b20  (
    .clk(clk100m),
    .d(\PWM3/n13 [20]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [20]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b21  (
    .clk(clk100m),
    .d(\PWM3/n13 [21]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [21]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b22  (
    .clk(clk100m),
    .d(\PWM3/n13 [22]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [22]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b23  (
    .clk(clk100m),
    .d(\PWM3/n13 [23]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [23]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b24  (
    .clk(clk100m),
    .d(\PWM3/n13 [24]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [24]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b25  (
    .clk(clk100m),
    .d(\PWM3/n13 [25]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [25]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b26  (
    .clk(clk100m),
    .d(\PWM3/n13 [26]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [26]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b3  (
    .clk(clk100m),
    .d(\PWM3/n13 [3]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [3]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b4  (
    .clk(clk100m),
    .d(\PWM3/n13 [4]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [4]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b5  (
    .clk(clk100m),
    .d(\PWM3/n13 [5]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [5]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b6  (
    .clk(clk100m),
    .d(\PWM3/n13 [6]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [6]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b7  (
    .clk(clk100m),
    .d(\PWM3/n13 [7]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [7]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b8  (
    .clk(clk100m),
    .d(\PWM3/n13 [8]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [8]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM3/reg0_b9  (
    .clk(clk100m),
    .d(\PWM3/n13 [9]),
    .en(1'b1),
    .reset(~\PWM3/n11 ),
    .set(1'b0),
    .q(\PWM3/FreCnt [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b0  (
    .clk(clk100m),
    .d(freq3[0]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [0]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b1  (
    .clk(clk100m),
    .d(freq3[1]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [1]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b10  (
    .clk(clk100m),
    .d(freq3[10]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [10]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b11  (
    .clk(clk100m),
    .d(freq3[11]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [11]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b12  (
    .clk(clk100m),
    .d(freq3[12]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [12]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b13  (
    .clk(clk100m),
    .d(freq3[13]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [13]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b14  (
    .clk(clk100m),
    .d(freq3[14]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [14]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b15  (
    .clk(clk100m),
    .d(freq3[15]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [15]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b16  (
    .clk(clk100m),
    .d(freq3[16]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [16]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b17  (
    .clk(clk100m),
    .d(freq3[17]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [17]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b18  (
    .clk(clk100m),
    .d(freq3[18]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [18]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b19  (
    .clk(clk100m),
    .d(freq3[19]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [19]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b2  (
    .clk(clk100m),
    .d(freq3[2]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [2]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b20  (
    .clk(clk100m),
    .d(freq3[20]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [20]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b21  (
    .clk(clk100m),
    .d(freq3[21]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [21]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b22  (
    .clk(clk100m),
    .d(freq3[22]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [22]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b23  (
    .clk(clk100m),
    .d(freq3[23]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [23]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b24  (
    .clk(clk100m),
    .d(freq3[24]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [24]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b25  (
    .clk(clk100m),
    .d(freq3[25]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [25]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b26  (
    .clk(clk100m),
    .d(freq3[26]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [26]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b3  (
    .clk(clk100m),
    .d(freq3[3]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [3]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b4  (
    .clk(clk100m),
    .d(freq3[4]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [4]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b5  (
    .clk(clk100m),
    .d(freq3[5]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [5]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b6  (
    .clk(clk100m),
    .d(freq3[6]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [6]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b7  (
    .clk(clk100m),
    .d(freq3[7]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [7]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b8  (
    .clk(clk100m),
    .d(freq3[8]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [8]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg1_b9  (
    .clk(clk100m),
    .d(freq3[9]),
    .en(\PWM3/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/FreCntr [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM3/reg2_b0  (
    .clk(clk100m),
    .d(\PWM3/n23 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[0]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b1  (
    .clk(clk100m),
    .d(\PWM3/n23 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[1]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b10  (
    .clk(clk100m),
    .d(\PWM3/n23 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[10]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b11  (
    .clk(clk100m),
    .d(\PWM3/n23 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[11]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b12  (
    .clk(clk100m),
    .d(\PWM3/n23 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[12]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b13  (
    .clk(clk100m),
    .d(\PWM3/n23 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[13]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b14  (
    .clk(clk100m),
    .d(\PWM3/n23 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[14]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b15  (
    .clk(clk100m),
    .d(\PWM3/n23 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[15]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b16  (
    .clk(clk100m),
    .d(\PWM3/n23 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[16]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b17  (
    .clk(clk100m),
    .d(\PWM3/n23 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[17]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b18  (
    .clk(clk100m),
    .d(\PWM3/n23 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[18]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b19  (
    .clk(clk100m),
    .d(\PWM3/n23 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[19]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b2  (
    .clk(clk100m),
    .d(\PWM3/n23 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[2]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b20  (
    .clk(clk100m),
    .d(\PWM3/n23 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[20]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b21  (
    .clk(clk100m),
    .d(\PWM3/n23 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[21]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b22  (
    .clk(clk100m),
    .d(\PWM3/n23 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[22]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b23  (
    .clk(clk100m),
    .d(\PWM3/n23 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[23]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b24  (
    .clk(clk100m),
    .d(\PWM3/n23 [24]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[24]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b25  (
    .clk(clk100m),
    .d(\PWM3/n23 [25]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[25]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b26  (
    .clk(clk100m),
    .d(\PWM3/n23 [26]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[26]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b27  (
    .clk(clk100m),
    .d(\PWM3/n23 [27]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[27]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b28  (
    .clk(clk100m),
    .d(\PWM3/n23 [28]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[28]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b29  (
    .clk(clk100m),
    .d(\PWM3/n23 [29]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[29]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b3  (
    .clk(clk100m),
    .d(\PWM3/n23 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[3]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b30  (
    .clk(clk100m),
    .d(\PWM3/n23 [30]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[30]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b31  (
    .clk(clk100m),
    .d(\PWM3/n23 [31]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[31]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b4  (
    .clk(clk100m),
    .d(\PWM3/n23 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[4]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b5  (
    .clk(clk100m),
    .d(\PWM3/n23 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[5]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b6  (
    .clk(clk100m),
    .d(\PWM3/n23 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[6]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b7  (
    .clk(clk100m),
    .d(\PWM3/n23 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[7]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b8  (
    .clk(clk100m),
    .d(\PWM3/n23 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[8]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg2_b9  (
    .clk(clk100m),
    .d(\PWM3/n23 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/pnumr[9]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM3/reg3_b0  (
    .clk(clk100m),
    .d(\PWM3/n31 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[0]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b1  (
    .clk(clk100m),
    .d(\PWM3/n31 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[1]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b10  (
    .clk(clk100m),
    .d(\PWM3/n31 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[10]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b11  (
    .clk(clk100m),
    .d(\PWM3/n31 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[11]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b12  (
    .clk(clk100m),
    .d(\PWM3/n31 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[12]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b13  (
    .clk(clk100m),
    .d(\PWM3/n31 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[13]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b14  (
    .clk(clk100m),
    .d(\PWM3/n31 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[14]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b15  (
    .clk(clk100m),
    .d(\PWM3/n31 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[15]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b16  (
    .clk(clk100m),
    .d(\PWM3/n31 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[16]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b17  (
    .clk(clk100m),
    .d(\PWM3/n31 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[17]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b18  (
    .clk(clk100m),
    .d(\PWM3/n31 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[18]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b19  (
    .clk(clk100m),
    .d(\PWM3/n31 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[19]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b2  (
    .clk(clk100m),
    .d(\PWM3/n31 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[2]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b20  (
    .clk(clk100m),
    .d(\PWM3/n31 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[20]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b21  (
    .clk(clk100m),
    .d(\PWM3/n31 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[21]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b22  (
    .clk(clk100m),
    .d(\PWM3/n31 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[22]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b23  (
    .clk(clk100m),
    .d(\PWM3/n31 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[23]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b3  (
    .clk(clk100m),
    .d(\PWM3/n31 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[3]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b4  (
    .clk(clk100m),
    .d(\PWM3/n31 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[4]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b5  (
    .clk(clk100m),
    .d(\PWM3/n31 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[5]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b6  (
    .clk(clk100m),
    .d(\PWM3/n31 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[6]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b7  (
    .clk(clk100m),
    .d(\PWM3/n31 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[7]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b8  (
    .clk(clk100m),
    .d(\PWM3/n31 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[8]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM3/reg3_b9  (
    .clk(clk100m),
    .d(\PWM3/n31 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM3/RemaTxNum[9]_keep ));  // src/OnePWM.v(58)
  reg_ar_ss_w1 \PWM3/stopreq_reg  (
    .clk(clk100m),
    .d(\PWM3/n1 ),
    .en(1'b1),
    .reset(1'b0),
    .set(pwm_start_stop[3]),
    .q(\PWM3/stopreq_keep ));  // src/OnePWM.v(15)
  add_pu27_mu27_o27 \PWM3/sub0  (
    .i0(\PWM3/FreCnt ),
    .i1(27'b000000000000000000000000001),
    .o(\PWM3/n12 [26:0]));  // src/OnePWM.v(32)
  add_pu24_mu24_o24 \PWM3/sub1  (
    .i0(pnumcnt3),
    .i1(24'b000000000000000000000001),
    .o(\PWM3/n26 [23:0]));  // src/OnePWM.v(55)
  AL_MUX \PWM3/u10  (
    .i0(1'b0),
    .i1(\PWM3/n9 ),
    .sel(n14),
    .o(\PWM3/n10 ));  // src/OnePWM.v(26)
  or \PWM3/u11  (\PWM3/n11 , pwm_state_read[3], pwm_start_stop[19]);  // src/OnePWM.v(30)
  and \PWM3/u14_sel_is_1  (\PWM3/u14_sel_is_1_o , pwm_state_read[3], \PWM3/n17_neg );
  and \PWM3/u15  (\PWM3/n24 , \PWM3/n0 , pwm_state_read[3]);  // src/OnePWM.v(54)
  and \PWM3/u17_sel_is_1  (\PWM3/u17_sel_is_1_o , \PWM3/n24 , \PWM3/n25_neg );
  not \PWM3/u17_sel_is_1_o_inv  (\PWM3/u17_sel_is_1_o_neg , \PWM3/u17_sel_is_1_o );
  AL_MUX \PWM3/u18  (
    .i0(\PWM3/pnumr [31]),
    .i1(dir[3]),
    .sel(\PWM3/u18_sel_is_0_o ),
    .o(\PWM3/n32 ));
  and \PWM3/u18_sel_is_0  (\PWM3/u18_sel_is_0_o , \pwm_start_stop[19]_neg , \PWM3/u17_sel_is_1_o_neg );
  AL_MUX \PWM3/u2  (
    .i0(\PWM3/stopreq ),
    .i1(1'b0),
    .sel(\PWM3/n0 ),
    .o(\PWM3/n1 ));  // src/OnePWM.v(15)
  and \PWM3/u5  (\PWM3/n4 , \PWM3/stopreq , \PWM3/n0 );  // src/OnePWM.v(23)
  and \PWM3/u6  (\PWM3/n6 , \PWM3/n5 , \PWM3/n0 );  // src/OnePWM.v(25)
  AL_MUX \PWM3/u8  (
    .i0(1'b0),
    .i1(pwm_state_read[3]),
    .sel(\PWM3/u8_sel_is_0_o ),
    .o(\PWM3/n8 ));
  and \PWM3/u8_sel_is_0  (\PWM3/u8_sel_is_0_o , \PWM3/n4_neg , \PWM3/n6_neg );
  AL_MUX \PWM3/u9  (
    .i0(\PWM3/n8 ),
    .i1(1'b1),
    .sel(pwm_start_stop[19]),
    .o(\PWM3/n9 ));  // src/OnePWM.v(26)
  reg_ar_as_w1 \PWM4/State_reg  (
    .clk(clk100m),
    .d(\PWM4/n10 ),
    .en(1'b1),
    .reset(~rstn),
    .set(1'b0),
    .q(pwm_state_read[4]));  // src/OnePWM.v(26)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[0]  (
    .i(\PWM4/RemaTxNum[0]_keep ),
    .o(pnumcnt4[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[10]  (
    .i(\PWM4/RemaTxNum[10]_keep ),
    .o(pnumcnt4[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[11]  (
    .i(\PWM4/RemaTxNum[11]_keep ),
    .o(pnumcnt4[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[12]  (
    .i(\PWM4/RemaTxNum[12]_keep ),
    .o(pnumcnt4[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[13]  (
    .i(\PWM4/RemaTxNum[13]_keep ),
    .o(pnumcnt4[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[14]  (
    .i(\PWM4/RemaTxNum[14]_keep ),
    .o(pnumcnt4[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[15]  (
    .i(\PWM4/RemaTxNum[15]_keep ),
    .o(pnumcnt4[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[16]  (
    .i(\PWM4/RemaTxNum[16]_keep ),
    .o(pnumcnt4[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[17]  (
    .i(\PWM4/RemaTxNum[17]_keep ),
    .o(pnumcnt4[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[18]  (
    .i(\PWM4/RemaTxNum[18]_keep ),
    .o(pnumcnt4[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[19]  (
    .i(\PWM4/RemaTxNum[19]_keep ),
    .o(pnumcnt4[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[1]  (
    .i(\PWM4/RemaTxNum[1]_keep ),
    .o(pnumcnt4[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[20]  (
    .i(\PWM4/RemaTxNum[20]_keep ),
    .o(pnumcnt4[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[21]  (
    .i(\PWM4/RemaTxNum[21]_keep ),
    .o(pnumcnt4[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[22]  (
    .i(\PWM4/RemaTxNum[22]_keep ),
    .o(pnumcnt4[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[23]  (
    .i(\PWM4/RemaTxNum[23]_keep ),
    .o(pnumcnt4[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[2]  (
    .i(\PWM4/RemaTxNum[2]_keep ),
    .o(pnumcnt4[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[3]  (
    .i(\PWM4/RemaTxNum[3]_keep ),
    .o(pnumcnt4[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[4]  (
    .i(\PWM4/RemaTxNum[4]_keep ),
    .o(pnumcnt4[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[5]  (
    .i(\PWM4/RemaTxNum[5]_keep ),
    .o(pnumcnt4[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[6]  (
    .i(\PWM4/RemaTxNum[6]_keep ),
    .o(pnumcnt4[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[7]  (
    .i(\PWM4/RemaTxNum[7]_keep ),
    .o(pnumcnt4[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[8]  (
    .i(\PWM4/RemaTxNum[8]_keep ),
    .o(pnumcnt4[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_RemaTxNum[9]  (
    .i(\PWM4/RemaTxNum[9]_keep ),
    .o(pnumcnt4[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_dir  (
    .i(\PWM4/dir_keep ),
    .o(dir[4]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[0]  (
    .i(\PWM4/pnumr[0]_keep ),
    .o(\PWM4/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[10]  (
    .i(\PWM4/pnumr[10]_keep ),
    .o(\PWM4/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[11]  (
    .i(\PWM4/pnumr[11]_keep ),
    .o(\PWM4/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[12]  (
    .i(\PWM4/pnumr[12]_keep ),
    .o(\PWM4/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[13]  (
    .i(\PWM4/pnumr[13]_keep ),
    .o(\PWM4/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[14]  (
    .i(\PWM4/pnumr[14]_keep ),
    .o(\PWM4/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[15]  (
    .i(\PWM4/pnumr[15]_keep ),
    .o(\PWM4/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[16]  (
    .i(\PWM4/pnumr[16]_keep ),
    .o(\PWM4/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[17]  (
    .i(\PWM4/pnumr[17]_keep ),
    .o(\PWM4/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[18]  (
    .i(\PWM4/pnumr[18]_keep ),
    .o(\PWM4/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[19]  (
    .i(\PWM4/pnumr[19]_keep ),
    .o(\PWM4/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[1]  (
    .i(\PWM4/pnumr[1]_keep ),
    .o(\PWM4/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[20]  (
    .i(\PWM4/pnumr[20]_keep ),
    .o(\PWM4/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[21]  (
    .i(\PWM4/pnumr[21]_keep ),
    .o(\PWM4/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[22]  (
    .i(\PWM4/pnumr[22]_keep ),
    .o(\PWM4/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[23]  (
    .i(\PWM4/pnumr[23]_keep ),
    .o(\PWM4/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[24]  (
    .i(\PWM4/pnumr[24]_keep ),
    .o(\PWM4/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[25]  (
    .i(\PWM4/pnumr[25]_keep ),
    .o(\PWM4/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[26]  (
    .i(\PWM4/pnumr[26]_keep ),
    .o(\PWM4/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[27]  (
    .i(\PWM4/pnumr[27]_keep ),
    .o(\PWM4/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[28]  (
    .i(\PWM4/pnumr[28]_keep ),
    .o(\PWM4/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[29]  (
    .i(\PWM4/pnumr[29]_keep ),
    .o(\PWM4/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[2]  (
    .i(\PWM4/pnumr[2]_keep ),
    .o(\PWM4/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[30]  (
    .i(\PWM4/pnumr[30]_keep ),
    .o(\PWM4/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[31]  (
    .i(\PWM4/pnumr[31]_keep ),
    .o(\PWM4/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[3]  (
    .i(\PWM4/pnumr[3]_keep ),
    .o(\PWM4/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[4]  (
    .i(\PWM4/pnumr[4]_keep ),
    .o(\PWM4/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[5]  (
    .i(\PWM4/pnumr[5]_keep ),
    .o(\PWM4/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[6]  (
    .i(\PWM4/pnumr[6]_keep ),
    .o(\PWM4/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[7]  (
    .i(\PWM4/pnumr[7]_keep ),
    .o(\PWM4/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[8]  (
    .i(\PWM4/pnumr[8]_keep ),
    .o(\PWM4/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pnumr[9]  (
    .i(\PWM4/pnumr[9]_keep ),
    .o(\PWM4/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_pwm  (
    .i(\PWM4/pwm_keep ),
    .o(pwm[4]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM4/_bufkeep_stopreq  (
    .i(\PWM4/stopreq_keep ),
    .o(\PWM4/stopreq ));  // src/OnePWM.v(14)
  reg_ar_as_w1 \PWM4/dir_reg  (
    .clk(clk100m),
    .d(\PWM4/n32 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/dir_keep ));  // src/OnePWM.v(58)
  eq_w27 \PWM4/eq0  (
    .i0(\PWM4/FreCnt ),
    .i1(27'b000000000000000000000000000),
    .o(\PWM4/n0 ));  // src/OnePWM.v(15)
  eq_w24 \PWM4/eq1  (
    .i0(pnumcnt4),
    .i1(24'b000000000000000000000001),
    .o(\PWM4/n5 ));  // src/OnePWM.v(25)
  eq_w27 \PWM4/eq2  (
    .i0(\PWM4/FreCnt ),
    .i1({1'b0,\PWM4/FreCntr [26:1]}),
    .o(\PWM4/n17 ));  // src/OnePWM.v(41)
  eq_w27 \PWM4/eq3  (
    .i0(\PWM4/FreCnt ),
    .i1(\PWM4/FreCntr ),
    .o(\PWM4/n18 ));  // src/OnePWM.v(43)
  binary_mux_s1_w1 \PWM4/mux0_b0  (
    .i0(\PWM4/n12 [0]),
    .i1(freq4[0]),
    .sel(\PWM4/n0 ),
    .o(\PWM4/n13 [0]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM4/mux0_b1  (
    .i0(\PWM4/n12 [1]),
    .i1(freq4[1]),
    .sel(\PWM4/n0 ),
    .o(\PWM4/n13 [1]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM4/mux0_b10  (
    .i0(\PWM4/n12 [10]),
    .i1(freq4[10]),
    .sel(\PWM4/n0 ),
    .o(\PWM4/n13 [10]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM4/mux0_b11  (
    .i0(\PWM4/n12 [11]),
    .i1(freq4[11]),
    .sel(\PWM4/n0 ),
    .o(\PWM4/n13 [11]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM4/mux0_b12  (
    .i0(\PWM4/n12 [12]),
    .i1(freq4[12]),
    .sel(\PWM4/n0 ),
    .o(\PWM4/n13 [12]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM4/mux0_b13  (
    .i0(\PWM4/n12 [13]),
    .i1(freq4[13]),
    .sel(\PWM4/n0 ),
    .o(\PWM4/n13 [13]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM4/mux0_b14  (
    .i0(\PWM4/n12 [14]),
    .i1(freq4[14]),
    .sel(\PWM4/n0 ),
    .o(\PWM4/n13 [14]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM4/mux0_b15  (
    .i0(\PWM4/n12 [15]),
    .i1(freq4[15]),
    .sel(\PWM4/n0 ),
    .o(\PWM4/n13 [15]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM4/mux0_b16  (
    .i0(\PWM4/n12 [16]),
    .i1(freq4[16]),
    .sel(\PWM4/n0 ),
    .o(\PWM4/n13 [16]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM4/mux0_b17  (
    .i0(\PWM4/n12 [17]),
    .i1(freq4[17]),
    .sel(\PWM4/n0 ),
    .o(\PWM4/n13 [17]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM4/mux0_b18  (
    .i0(\PWM4/n12 [18]),
    .i1(freq4[18]),
    .sel(\PWM4/n0 ),
    .o(\PWM4/n13 [18]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM4/mux0_b19  (
    .i0(\PWM4/n12 [19]),
    .i1(freq4[19]),
    .sel(\PWM4/n0 ),
    .o(\PWM4/n13 [19]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM4/mux0_b2  (
    .i0(\PWM4/n12 [2]),
    .i1(freq4[2]),
    .sel(\PWM4/n0 ),
    .o(\PWM4/n13 [2]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM4/mux0_b20  (
    .i0(\PWM4/n12 [20]),
    .i1(freq4[20]),
    .sel(\PWM4/n0 ),
    .o(\PWM4/n13 [20]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM4/mux0_b21  (
    .i0(\PWM4/n12 [21]),
    .i1(freq4[21]),
    .sel(\PWM4/n0 ),
    .o(\PWM4/n13 [21]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM4/mux0_b22  (
    .i0(\PWM4/n12 [22]),
    .i1(freq4[22]),
    .sel(\PWM4/n0 ),
    .o(\PWM4/n13 [22]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM4/mux0_b23  (
    .i0(\PWM4/n12 [23]),
    .i1(freq4[23]),
    .sel(\PWM4/n0 ),
    .o(\PWM4/n13 [23]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM4/mux0_b24  (
    .i0(\PWM4/n12 [24]),
    .i1(freq4[24]),
    .sel(\PWM4/n0 ),
    .o(\PWM4/n13 [24]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM4/mux0_b25  (
    .i0(\PWM4/n12 [25]),
    .i1(freq4[25]),
    .sel(\PWM4/n0 ),
    .o(\PWM4/n13 [25]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM4/mux0_b26  (
    .i0(\PWM4/n12 [26]),
    .i1(freq4[26]),
    .sel(\PWM4/n0 ),
    .o(\PWM4/n13 [26]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM4/mux0_b3  (
    .i0(\PWM4/n12 [3]),
    .i1(freq4[3]),
    .sel(\PWM4/n0 ),
    .o(\PWM4/n13 [3]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM4/mux0_b4  (
    .i0(\PWM4/n12 [4]),
    .i1(freq4[4]),
    .sel(\PWM4/n0 ),
    .o(\PWM4/n13 [4]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM4/mux0_b5  (
    .i0(\PWM4/n12 [5]),
    .i1(freq4[5]),
    .sel(\PWM4/n0 ),
    .o(\PWM4/n13 [5]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM4/mux0_b6  (
    .i0(\PWM4/n12 [6]),
    .i1(freq4[6]),
    .sel(\PWM4/n0 ),
    .o(\PWM4/n13 [6]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM4/mux0_b7  (
    .i0(\PWM4/n12 [7]),
    .i1(freq4[7]),
    .sel(\PWM4/n0 ),
    .o(\PWM4/n13 [7]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM4/mux0_b8  (
    .i0(\PWM4/n12 [8]),
    .i1(freq4[8]),
    .sel(\PWM4/n0 ),
    .o(\PWM4/n13 [8]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM4/mux0_b9  (
    .i0(\PWM4/n12 [9]),
    .i1(freq4[9]),
    .sel(\PWM4/n0 ),
    .o(\PWM4/n13 [9]));  // src/OnePWM.v(32)
  and \PWM4/mux3_b0_sel_is_3  (\PWM4/mux3_b0_sel_is_3_o , \PWM4/n11 , \PWM4/n0 );
  binary_mux_s1_w1 \PWM4/mux4_b0  (
    .i0(\PWM4/pnumr [0]),
    .i1(1'b0),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n22 [0]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux4_b1  (
    .i0(\PWM4/pnumr [1]),
    .i1(1'b0),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n22 [1]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux4_b10  (
    .i0(\PWM4/pnumr [10]),
    .i1(1'b0),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n22 [10]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux4_b11  (
    .i0(\PWM4/pnumr [11]),
    .i1(1'b0),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n22 [11]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux4_b12  (
    .i0(\PWM4/pnumr [12]),
    .i1(1'b0),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n22 [12]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux4_b13  (
    .i0(\PWM4/pnumr [13]),
    .i1(1'b0),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n22 [13]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux4_b14  (
    .i0(\PWM4/pnumr [14]),
    .i1(1'b0),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n22 [14]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux4_b15  (
    .i0(\PWM4/pnumr [15]),
    .i1(1'b0),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n22 [15]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux4_b16  (
    .i0(\PWM4/pnumr [16]),
    .i1(1'b0),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n22 [16]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux4_b17  (
    .i0(\PWM4/pnumr [17]),
    .i1(1'b0),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n22 [17]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux4_b18  (
    .i0(\PWM4/pnumr [18]),
    .i1(1'b0),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n22 [18]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux4_b19  (
    .i0(\PWM4/pnumr [19]),
    .i1(1'b0),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n22 [19]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux4_b2  (
    .i0(\PWM4/pnumr [2]),
    .i1(1'b0),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n22 [2]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux4_b20  (
    .i0(\PWM4/pnumr [20]),
    .i1(1'b0),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n22 [20]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux4_b21  (
    .i0(\PWM4/pnumr [21]),
    .i1(1'b0),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n22 [21]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux4_b22  (
    .i0(\PWM4/pnumr [22]),
    .i1(1'b0),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n22 [22]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux4_b23  (
    .i0(\PWM4/pnumr [23]),
    .i1(1'b0),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n22 [23]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux4_b24  (
    .i0(\PWM4/pnumr [24]),
    .i1(1'b0),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n22 [24]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux4_b25  (
    .i0(\PWM4/pnumr [25]),
    .i1(1'b0),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n22 [25]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux4_b26  (
    .i0(\PWM4/pnumr [26]),
    .i1(1'b0),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n22 [26]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux4_b27  (
    .i0(\PWM4/pnumr [27]),
    .i1(1'b0),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n22 [27]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux4_b28  (
    .i0(\PWM4/pnumr [28]),
    .i1(1'b0),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n22 [28]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux4_b29  (
    .i0(\PWM4/pnumr [29]),
    .i1(1'b0),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n22 [29]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux4_b3  (
    .i0(\PWM4/pnumr [3]),
    .i1(1'b0),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n22 [3]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux4_b30  (
    .i0(\PWM4/pnumr [30]),
    .i1(1'b0),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n22 [30]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux4_b31  (
    .i0(\PWM4/pnumr [31]),
    .i1(1'b0),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n22 [31]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux4_b4  (
    .i0(\PWM4/pnumr [4]),
    .i1(1'b0),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n22 [4]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux4_b5  (
    .i0(\PWM4/pnumr [5]),
    .i1(1'b0),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n22 [5]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux4_b6  (
    .i0(\PWM4/pnumr [6]),
    .i1(1'b0),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n22 [6]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux4_b7  (
    .i0(\PWM4/pnumr [7]),
    .i1(1'b0),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n22 [7]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux4_b8  (
    .i0(\PWM4/pnumr [8]),
    .i1(1'b0),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n22 [8]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux4_b9  (
    .i0(\PWM4/pnumr [9]),
    .i1(1'b0),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n22 [9]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux5_b0  (
    .i0(\PWM4/n22 [0]),
    .i1(pnum4[0]),
    .sel(pnum4[32]),
    .o(\PWM4/n23 [0]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux5_b1  (
    .i0(\PWM4/n22 [1]),
    .i1(pnum4[1]),
    .sel(pnum4[32]),
    .o(\PWM4/n23 [1]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux5_b10  (
    .i0(\PWM4/n22 [10]),
    .i1(pnum4[10]),
    .sel(pnum4[32]),
    .o(\PWM4/n23 [10]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux5_b11  (
    .i0(\PWM4/n22 [11]),
    .i1(pnum4[11]),
    .sel(pnum4[32]),
    .o(\PWM4/n23 [11]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux5_b12  (
    .i0(\PWM4/n22 [12]),
    .i1(pnum4[12]),
    .sel(pnum4[32]),
    .o(\PWM4/n23 [12]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux5_b13  (
    .i0(\PWM4/n22 [13]),
    .i1(pnum4[13]),
    .sel(pnum4[32]),
    .o(\PWM4/n23 [13]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux5_b14  (
    .i0(\PWM4/n22 [14]),
    .i1(pnum4[14]),
    .sel(pnum4[32]),
    .o(\PWM4/n23 [14]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux5_b15  (
    .i0(\PWM4/n22 [15]),
    .i1(pnum4[15]),
    .sel(pnum4[32]),
    .o(\PWM4/n23 [15]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux5_b16  (
    .i0(\PWM4/n22 [16]),
    .i1(pnum4[16]),
    .sel(pnum4[32]),
    .o(\PWM4/n23 [16]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux5_b17  (
    .i0(\PWM4/n22 [17]),
    .i1(pnum4[17]),
    .sel(pnum4[32]),
    .o(\PWM4/n23 [17]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux5_b18  (
    .i0(\PWM4/n22 [18]),
    .i1(pnum4[18]),
    .sel(pnum4[32]),
    .o(\PWM4/n23 [18]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux5_b19  (
    .i0(\PWM4/n22 [19]),
    .i1(pnum4[19]),
    .sel(pnum4[32]),
    .o(\PWM4/n23 [19]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux5_b2  (
    .i0(\PWM4/n22 [2]),
    .i1(pnum4[2]),
    .sel(pnum4[32]),
    .o(\PWM4/n23 [2]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux5_b20  (
    .i0(\PWM4/n22 [20]),
    .i1(pnum4[20]),
    .sel(pnum4[32]),
    .o(\PWM4/n23 [20]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux5_b21  (
    .i0(\PWM4/n22 [21]),
    .i1(pnum4[21]),
    .sel(pnum4[32]),
    .o(\PWM4/n23 [21]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux5_b22  (
    .i0(\PWM4/n22 [22]),
    .i1(pnum4[22]),
    .sel(pnum4[32]),
    .o(\PWM4/n23 [22]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux5_b23  (
    .i0(\PWM4/n22 [23]),
    .i1(pnum4[23]),
    .sel(pnum4[32]),
    .o(\PWM4/n23 [23]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux5_b24  (
    .i0(\PWM4/n22 [24]),
    .i1(pnum4[24]),
    .sel(pnum4[32]),
    .o(\PWM4/n23 [24]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux5_b25  (
    .i0(\PWM4/n22 [25]),
    .i1(pnum4[25]),
    .sel(pnum4[32]),
    .o(\PWM4/n23 [25]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux5_b26  (
    .i0(\PWM4/n22 [26]),
    .i1(pnum4[26]),
    .sel(pnum4[32]),
    .o(\PWM4/n23 [26]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux5_b27  (
    .i0(\PWM4/n22 [27]),
    .i1(pnum4[27]),
    .sel(pnum4[32]),
    .o(\PWM4/n23 [27]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux5_b28  (
    .i0(\PWM4/n22 [28]),
    .i1(pnum4[28]),
    .sel(pnum4[32]),
    .o(\PWM4/n23 [28]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux5_b29  (
    .i0(\PWM4/n22 [29]),
    .i1(pnum4[29]),
    .sel(pnum4[32]),
    .o(\PWM4/n23 [29]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux5_b3  (
    .i0(\PWM4/n22 [3]),
    .i1(pnum4[3]),
    .sel(pnum4[32]),
    .o(\PWM4/n23 [3]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux5_b30  (
    .i0(\PWM4/n22 [30]),
    .i1(pnum4[30]),
    .sel(pnum4[32]),
    .o(\PWM4/n23 [30]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux5_b31  (
    .i0(\PWM4/n22 [31]),
    .i1(pnum4[31]),
    .sel(pnum4[32]),
    .o(\PWM4/n23 [31]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux5_b4  (
    .i0(\PWM4/n22 [4]),
    .i1(pnum4[4]),
    .sel(pnum4[32]),
    .o(\PWM4/n23 [4]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux5_b5  (
    .i0(\PWM4/n22 [5]),
    .i1(pnum4[5]),
    .sel(pnum4[32]),
    .o(\PWM4/n23 [5]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux5_b6  (
    .i0(\PWM4/n22 [6]),
    .i1(pnum4[6]),
    .sel(pnum4[32]),
    .o(\PWM4/n23 [6]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux5_b7  (
    .i0(\PWM4/n22 [7]),
    .i1(pnum4[7]),
    .sel(pnum4[32]),
    .o(\PWM4/n23 [7]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux5_b8  (
    .i0(\PWM4/n22 [8]),
    .i1(pnum4[8]),
    .sel(pnum4[32]),
    .o(\PWM4/n23 [8]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux5_b9  (
    .i0(\PWM4/n22 [9]),
    .i1(pnum4[9]),
    .sel(pnum4[32]),
    .o(\PWM4/n23 [9]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM4/mux6_b0  (
    .i0(\PWM4/pnumr [0]),
    .i1(\PWM4/n26 [0]),
    .sel(\PWM4/n25 ),
    .o(\PWM4/n27 [0]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM4/mux6_b1  (
    .i0(\PWM4/pnumr [1]),
    .i1(\PWM4/n26 [1]),
    .sel(\PWM4/n25 ),
    .o(\PWM4/n27 [1]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM4/mux6_b10  (
    .i0(\PWM4/pnumr [10]),
    .i1(\PWM4/n26 [10]),
    .sel(\PWM4/n25 ),
    .o(\PWM4/n27 [10]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM4/mux6_b11  (
    .i0(\PWM4/pnumr [11]),
    .i1(\PWM4/n26 [11]),
    .sel(\PWM4/n25 ),
    .o(\PWM4/n27 [11]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM4/mux6_b12  (
    .i0(\PWM4/pnumr [12]),
    .i1(\PWM4/n26 [12]),
    .sel(\PWM4/n25 ),
    .o(\PWM4/n27 [12]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM4/mux6_b13  (
    .i0(\PWM4/pnumr [13]),
    .i1(\PWM4/n26 [13]),
    .sel(\PWM4/n25 ),
    .o(\PWM4/n27 [13]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM4/mux6_b14  (
    .i0(\PWM4/pnumr [14]),
    .i1(\PWM4/n26 [14]),
    .sel(\PWM4/n25 ),
    .o(\PWM4/n27 [14]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM4/mux6_b15  (
    .i0(\PWM4/pnumr [15]),
    .i1(\PWM4/n26 [15]),
    .sel(\PWM4/n25 ),
    .o(\PWM4/n27 [15]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM4/mux6_b16  (
    .i0(\PWM4/pnumr [16]),
    .i1(\PWM4/n26 [16]),
    .sel(\PWM4/n25 ),
    .o(\PWM4/n27 [16]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM4/mux6_b17  (
    .i0(\PWM4/pnumr [17]),
    .i1(\PWM4/n26 [17]),
    .sel(\PWM4/n25 ),
    .o(\PWM4/n27 [17]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM4/mux6_b18  (
    .i0(\PWM4/pnumr [18]),
    .i1(\PWM4/n26 [18]),
    .sel(\PWM4/n25 ),
    .o(\PWM4/n27 [18]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM4/mux6_b19  (
    .i0(\PWM4/pnumr [19]),
    .i1(\PWM4/n26 [19]),
    .sel(\PWM4/n25 ),
    .o(\PWM4/n27 [19]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM4/mux6_b2  (
    .i0(\PWM4/pnumr [2]),
    .i1(\PWM4/n26 [2]),
    .sel(\PWM4/n25 ),
    .o(\PWM4/n27 [2]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM4/mux6_b20  (
    .i0(\PWM4/pnumr [20]),
    .i1(\PWM4/n26 [20]),
    .sel(\PWM4/n25 ),
    .o(\PWM4/n27 [20]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM4/mux6_b21  (
    .i0(\PWM4/pnumr [21]),
    .i1(\PWM4/n26 [21]),
    .sel(\PWM4/n25 ),
    .o(\PWM4/n27 [21]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM4/mux6_b22  (
    .i0(\PWM4/pnumr [22]),
    .i1(\PWM4/n26 [22]),
    .sel(\PWM4/n25 ),
    .o(\PWM4/n27 [22]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM4/mux6_b23  (
    .i0(\PWM4/pnumr [23]),
    .i1(\PWM4/n26 [23]),
    .sel(\PWM4/n25 ),
    .o(\PWM4/n27 [23]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM4/mux6_b3  (
    .i0(\PWM4/pnumr [3]),
    .i1(\PWM4/n26 [3]),
    .sel(\PWM4/n25 ),
    .o(\PWM4/n27 [3]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM4/mux6_b4  (
    .i0(\PWM4/pnumr [4]),
    .i1(\PWM4/n26 [4]),
    .sel(\PWM4/n25 ),
    .o(\PWM4/n27 [4]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM4/mux6_b5  (
    .i0(\PWM4/pnumr [5]),
    .i1(\PWM4/n26 [5]),
    .sel(\PWM4/n25 ),
    .o(\PWM4/n27 [5]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM4/mux6_b6  (
    .i0(\PWM4/pnumr [6]),
    .i1(\PWM4/n26 [6]),
    .sel(\PWM4/n25 ),
    .o(\PWM4/n27 [6]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM4/mux6_b7  (
    .i0(\PWM4/pnumr [7]),
    .i1(\PWM4/n26 [7]),
    .sel(\PWM4/n25 ),
    .o(\PWM4/n27 [7]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM4/mux6_b8  (
    .i0(\PWM4/pnumr [8]),
    .i1(\PWM4/n26 [8]),
    .sel(\PWM4/n25 ),
    .o(\PWM4/n27 [8]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM4/mux6_b9  (
    .i0(\PWM4/pnumr [9]),
    .i1(\PWM4/n26 [9]),
    .sel(\PWM4/n25 ),
    .o(\PWM4/n27 [9]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM4/mux7_b0  (
    .i0(pnumcnt4[0]),
    .i1(\PWM4/n27 [0]),
    .sel(\PWM4/n24 ),
    .o(\PWM4/n29 [0]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux7_b1  (
    .i0(pnumcnt4[1]),
    .i1(\PWM4/n27 [1]),
    .sel(\PWM4/n24 ),
    .o(\PWM4/n29 [1]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux7_b10  (
    .i0(pnumcnt4[10]),
    .i1(\PWM4/n27 [10]),
    .sel(\PWM4/n24 ),
    .o(\PWM4/n29 [10]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux7_b11  (
    .i0(pnumcnt4[11]),
    .i1(\PWM4/n27 [11]),
    .sel(\PWM4/n24 ),
    .o(\PWM4/n29 [11]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux7_b12  (
    .i0(pnumcnt4[12]),
    .i1(\PWM4/n27 [12]),
    .sel(\PWM4/n24 ),
    .o(\PWM4/n29 [12]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux7_b13  (
    .i0(pnumcnt4[13]),
    .i1(\PWM4/n27 [13]),
    .sel(\PWM4/n24 ),
    .o(\PWM4/n29 [13]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux7_b14  (
    .i0(pnumcnt4[14]),
    .i1(\PWM4/n27 [14]),
    .sel(\PWM4/n24 ),
    .o(\PWM4/n29 [14]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux7_b15  (
    .i0(pnumcnt4[15]),
    .i1(\PWM4/n27 [15]),
    .sel(\PWM4/n24 ),
    .o(\PWM4/n29 [15]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux7_b16  (
    .i0(pnumcnt4[16]),
    .i1(\PWM4/n27 [16]),
    .sel(\PWM4/n24 ),
    .o(\PWM4/n29 [16]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux7_b17  (
    .i0(pnumcnt4[17]),
    .i1(\PWM4/n27 [17]),
    .sel(\PWM4/n24 ),
    .o(\PWM4/n29 [17]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux7_b18  (
    .i0(pnumcnt4[18]),
    .i1(\PWM4/n27 [18]),
    .sel(\PWM4/n24 ),
    .o(\PWM4/n29 [18]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux7_b19  (
    .i0(pnumcnt4[19]),
    .i1(\PWM4/n27 [19]),
    .sel(\PWM4/n24 ),
    .o(\PWM4/n29 [19]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux7_b2  (
    .i0(pnumcnt4[2]),
    .i1(\PWM4/n27 [2]),
    .sel(\PWM4/n24 ),
    .o(\PWM4/n29 [2]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux7_b20  (
    .i0(pnumcnt4[20]),
    .i1(\PWM4/n27 [20]),
    .sel(\PWM4/n24 ),
    .o(\PWM4/n29 [20]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux7_b21  (
    .i0(pnumcnt4[21]),
    .i1(\PWM4/n27 [21]),
    .sel(\PWM4/n24 ),
    .o(\PWM4/n29 [21]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux7_b22  (
    .i0(pnumcnt4[22]),
    .i1(\PWM4/n27 [22]),
    .sel(\PWM4/n24 ),
    .o(\PWM4/n29 [22]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux7_b23  (
    .i0(pnumcnt4[23]),
    .i1(\PWM4/n27 [23]),
    .sel(\PWM4/n24 ),
    .o(\PWM4/n29 [23]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux7_b3  (
    .i0(pnumcnt4[3]),
    .i1(\PWM4/n27 [3]),
    .sel(\PWM4/n24 ),
    .o(\PWM4/n29 [3]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux7_b4  (
    .i0(pnumcnt4[4]),
    .i1(\PWM4/n27 [4]),
    .sel(\PWM4/n24 ),
    .o(\PWM4/n29 [4]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux7_b5  (
    .i0(pnumcnt4[5]),
    .i1(\PWM4/n27 [5]),
    .sel(\PWM4/n24 ),
    .o(\PWM4/n29 [5]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux7_b6  (
    .i0(pnumcnt4[6]),
    .i1(\PWM4/n27 [6]),
    .sel(\PWM4/n24 ),
    .o(\PWM4/n29 [6]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux7_b7  (
    .i0(pnumcnt4[7]),
    .i1(\PWM4/n27 [7]),
    .sel(\PWM4/n24 ),
    .o(\PWM4/n29 [7]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux7_b8  (
    .i0(pnumcnt4[8]),
    .i1(\PWM4/n27 [8]),
    .sel(\PWM4/n24 ),
    .o(\PWM4/n29 [8]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux7_b9  (
    .i0(pnumcnt4[9]),
    .i1(\PWM4/n27 [9]),
    .sel(\PWM4/n24 ),
    .o(\PWM4/n29 [9]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux8_b0  (
    .i0(\PWM4/n29 [0]),
    .i1(\PWM4/pnumr [0]),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n31 [0]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux8_b1  (
    .i0(\PWM4/n29 [1]),
    .i1(\PWM4/pnumr [1]),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n31 [1]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux8_b10  (
    .i0(\PWM4/n29 [10]),
    .i1(\PWM4/pnumr [10]),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n31 [10]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux8_b11  (
    .i0(\PWM4/n29 [11]),
    .i1(\PWM4/pnumr [11]),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n31 [11]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux8_b12  (
    .i0(\PWM4/n29 [12]),
    .i1(\PWM4/pnumr [12]),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n31 [12]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux8_b13  (
    .i0(\PWM4/n29 [13]),
    .i1(\PWM4/pnumr [13]),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n31 [13]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux8_b14  (
    .i0(\PWM4/n29 [14]),
    .i1(\PWM4/pnumr [14]),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n31 [14]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux8_b15  (
    .i0(\PWM4/n29 [15]),
    .i1(\PWM4/pnumr [15]),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n31 [15]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux8_b16  (
    .i0(\PWM4/n29 [16]),
    .i1(\PWM4/pnumr [16]),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n31 [16]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux8_b17  (
    .i0(\PWM4/n29 [17]),
    .i1(\PWM4/pnumr [17]),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n31 [17]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux8_b18  (
    .i0(\PWM4/n29 [18]),
    .i1(\PWM4/pnumr [18]),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n31 [18]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux8_b19  (
    .i0(\PWM4/n29 [19]),
    .i1(\PWM4/pnumr [19]),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n31 [19]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux8_b2  (
    .i0(\PWM4/n29 [2]),
    .i1(\PWM4/pnumr [2]),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n31 [2]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux8_b20  (
    .i0(\PWM4/n29 [20]),
    .i1(\PWM4/pnumr [20]),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n31 [20]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux8_b21  (
    .i0(\PWM4/n29 [21]),
    .i1(\PWM4/pnumr [21]),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n31 [21]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux8_b22  (
    .i0(\PWM4/n29 [22]),
    .i1(\PWM4/pnumr [22]),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n31 [22]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux8_b23  (
    .i0(\PWM4/n29 [23]),
    .i1(\PWM4/pnumr [23]),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n31 [23]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux8_b3  (
    .i0(\PWM4/n29 [3]),
    .i1(\PWM4/pnumr [3]),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n31 [3]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux8_b4  (
    .i0(\PWM4/n29 [4]),
    .i1(\PWM4/pnumr [4]),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n31 [4]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux8_b5  (
    .i0(\PWM4/n29 [5]),
    .i1(\PWM4/pnumr [5]),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n31 [5]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux8_b6  (
    .i0(\PWM4/n29 [6]),
    .i1(\PWM4/pnumr [6]),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n31 [6]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux8_b7  (
    .i0(\PWM4/n29 [7]),
    .i1(\PWM4/pnumr [7]),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n31 [7]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux8_b8  (
    .i0(\PWM4/n29 [8]),
    .i1(\PWM4/pnumr [8]),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n31 [8]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM4/mux8_b9  (
    .i0(\PWM4/n29 [9]),
    .i1(\PWM4/pnumr [9]),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n31 [9]));  // src/OnePWM.v(57)
  not \PWM4/n17_inv  (\PWM4/n17_neg , \PWM4/n17 );
  not \PWM4/n25_inv  (\PWM4/n25_neg , \PWM4/n25 );
  not \PWM4/n4_inv  (\PWM4/n4_neg , \PWM4/n4 );
  not \PWM4/n6_inv  (\PWM4/n6_neg , \PWM4/n6 );
  ne_w24 \PWM4/neq0  (
    .i0(pnumcnt4),
    .i1(24'b000000000000000000000000),
    .o(\PWM4/n25 ));  // src/OnePWM.v(55)
  reg_sr_ss_w1 \PWM4/pwm_reg  (
    .clk(clk100m),
    .d(pwm[4]),
    .en(1'b1),
    .reset(~\PWM4/u14_sel_is_1_o ),
    .set(\PWM4/n18 ),
    .q(\PWM4/pwm_keep ));  // src/OnePWM.v(45)
  reg_sr_as_w1 \PWM4/reg0_b0  (
    .clk(clk100m),
    .d(\PWM4/n13 [0]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [0]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b1  (
    .clk(clk100m),
    .d(\PWM4/n13 [1]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [1]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b10  (
    .clk(clk100m),
    .d(\PWM4/n13 [10]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [10]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b11  (
    .clk(clk100m),
    .d(\PWM4/n13 [11]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [11]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b12  (
    .clk(clk100m),
    .d(\PWM4/n13 [12]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [12]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b13  (
    .clk(clk100m),
    .d(\PWM4/n13 [13]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [13]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b14  (
    .clk(clk100m),
    .d(\PWM4/n13 [14]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [14]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b15  (
    .clk(clk100m),
    .d(\PWM4/n13 [15]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [15]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b16  (
    .clk(clk100m),
    .d(\PWM4/n13 [16]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [16]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b17  (
    .clk(clk100m),
    .d(\PWM4/n13 [17]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [17]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b18  (
    .clk(clk100m),
    .d(\PWM4/n13 [18]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [18]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b19  (
    .clk(clk100m),
    .d(\PWM4/n13 [19]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [19]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b2  (
    .clk(clk100m),
    .d(\PWM4/n13 [2]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [2]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b20  (
    .clk(clk100m),
    .d(\PWM4/n13 [20]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [20]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b21  (
    .clk(clk100m),
    .d(\PWM4/n13 [21]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [21]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b22  (
    .clk(clk100m),
    .d(\PWM4/n13 [22]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [22]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b23  (
    .clk(clk100m),
    .d(\PWM4/n13 [23]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [23]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b24  (
    .clk(clk100m),
    .d(\PWM4/n13 [24]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [24]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b25  (
    .clk(clk100m),
    .d(\PWM4/n13 [25]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [25]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b26  (
    .clk(clk100m),
    .d(\PWM4/n13 [26]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [26]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b3  (
    .clk(clk100m),
    .d(\PWM4/n13 [3]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [3]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b4  (
    .clk(clk100m),
    .d(\PWM4/n13 [4]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [4]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b5  (
    .clk(clk100m),
    .d(\PWM4/n13 [5]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [5]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b6  (
    .clk(clk100m),
    .d(\PWM4/n13 [6]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [6]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b7  (
    .clk(clk100m),
    .d(\PWM4/n13 [7]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [7]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b8  (
    .clk(clk100m),
    .d(\PWM4/n13 [8]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [8]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM4/reg0_b9  (
    .clk(clk100m),
    .d(\PWM4/n13 [9]),
    .en(1'b1),
    .reset(~\PWM4/n11 ),
    .set(1'b0),
    .q(\PWM4/FreCnt [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b0  (
    .clk(clk100m),
    .d(freq4[0]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [0]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b1  (
    .clk(clk100m),
    .d(freq4[1]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [1]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b10  (
    .clk(clk100m),
    .d(freq4[10]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [10]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b11  (
    .clk(clk100m),
    .d(freq4[11]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [11]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b12  (
    .clk(clk100m),
    .d(freq4[12]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [12]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b13  (
    .clk(clk100m),
    .d(freq4[13]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [13]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b14  (
    .clk(clk100m),
    .d(freq4[14]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [14]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b15  (
    .clk(clk100m),
    .d(freq4[15]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [15]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b16  (
    .clk(clk100m),
    .d(freq4[16]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [16]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b17  (
    .clk(clk100m),
    .d(freq4[17]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [17]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b18  (
    .clk(clk100m),
    .d(freq4[18]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [18]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b19  (
    .clk(clk100m),
    .d(freq4[19]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [19]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b2  (
    .clk(clk100m),
    .d(freq4[2]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [2]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b20  (
    .clk(clk100m),
    .d(freq4[20]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [20]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b21  (
    .clk(clk100m),
    .d(freq4[21]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [21]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b22  (
    .clk(clk100m),
    .d(freq4[22]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [22]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b23  (
    .clk(clk100m),
    .d(freq4[23]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [23]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b24  (
    .clk(clk100m),
    .d(freq4[24]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [24]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b25  (
    .clk(clk100m),
    .d(freq4[25]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [25]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b26  (
    .clk(clk100m),
    .d(freq4[26]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [26]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b3  (
    .clk(clk100m),
    .d(freq4[3]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [3]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b4  (
    .clk(clk100m),
    .d(freq4[4]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [4]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b5  (
    .clk(clk100m),
    .d(freq4[5]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [5]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b6  (
    .clk(clk100m),
    .d(freq4[6]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [6]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b7  (
    .clk(clk100m),
    .d(freq4[7]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [7]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b8  (
    .clk(clk100m),
    .d(freq4[8]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [8]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg1_b9  (
    .clk(clk100m),
    .d(freq4[9]),
    .en(\PWM4/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/FreCntr [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM4/reg2_b0  (
    .clk(clk100m),
    .d(\PWM4/n23 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[0]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b1  (
    .clk(clk100m),
    .d(\PWM4/n23 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[1]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b10  (
    .clk(clk100m),
    .d(\PWM4/n23 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[10]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b11  (
    .clk(clk100m),
    .d(\PWM4/n23 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[11]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b12  (
    .clk(clk100m),
    .d(\PWM4/n23 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[12]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b13  (
    .clk(clk100m),
    .d(\PWM4/n23 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[13]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b14  (
    .clk(clk100m),
    .d(\PWM4/n23 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[14]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b15  (
    .clk(clk100m),
    .d(\PWM4/n23 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[15]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b16  (
    .clk(clk100m),
    .d(\PWM4/n23 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[16]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b17  (
    .clk(clk100m),
    .d(\PWM4/n23 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[17]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b18  (
    .clk(clk100m),
    .d(\PWM4/n23 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[18]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b19  (
    .clk(clk100m),
    .d(\PWM4/n23 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[19]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b2  (
    .clk(clk100m),
    .d(\PWM4/n23 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[2]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b20  (
    .clk(clk100m),
    .d(\PWM4/n23 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[20]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b21  (
    .clk(clk100m),
    .d(\PWM4/n23 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[21]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b22  (
    .clk(clk100m),
    .d(\PWM4/n23 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[22]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b23  (
    .clk(clk100m),
    .d(\PWM4/n23 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[23]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b24  (
    .clk(clk100m),
    .d(\PWM4/n23 [24]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[24]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b25  (
    .clk(clk100m),
    .d(\PWM4/n23 [25]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[25]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b26  (
    .clk(clk100m),
    .d(\PWM4/n23 [26]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[26]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b27  (
    .clk(clk100m),
    .d(\PWM4/n23 [27]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[27]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b28  (
    .clk(clk100m),
    .d(\PWM4/n23 [28]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[28]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b29  (
    .clk(clk100m),
    .d(\PWM4/n23 [29]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[29]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b3  (
    .clk(clk100m),
    .d(\PWM4/n23 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[3]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b30  (
    .clk(clk100m),
    .d(\PWM4/n23 [30]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[30]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b31  (
    .clk(clk100m),
    .d(\PWM4/n23 [31]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[31]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b4  (
    .clk(clk100m),
    .d(\PWM4/n23 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[4]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b5  (
    .clk(clk100m),
    .d(\PWM4/n23 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[5]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b6  (
    .clk(clk100m),
    .d(\PWM4/n23 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[6]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b7  (
    .clk(clk100m),
    .d(\PWM4/n23 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[7]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b8  (
    .clk(clk100m),
    .d(\PWM4/n23 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[8]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg2_b9  (
    .clk(clk100m),
    .d(\PWM4/n23 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/pnumr[9]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM4/reg3_b0  (
    .clk(clk100m),
    .d(\PWM4/n31 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[0]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b1  (
    .clk(clk100m),
    .d(\PWM4/n31 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[1]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b10  (
    .clk(clk100m),
    .d(\PWM4/n31 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[10]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b11  (
    .clk(clk100m),
    .d(\PWM4/n31 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[11]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b12  (
    .clk(clk100m),
    .d(\PWM4/n31 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[12]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b13  (
    .clk(clk100m),
    .d(\PWM4/n31 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[13]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b14  (
    .clk(clk100m),
    .d(\PWM4/n31 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[14]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b15  (
    .clk(clk100m),
    .d(\PWM4/n31 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[15]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b16  (
    .clk(clk100m),
    .d(\PWM4/n31 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[16]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b17  (
    .clk(clk100m),
    .d(\PWM4/n31 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[17]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b18  (
    .clk(clk100m),
    .d(\PWM4/n31 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[18]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b19  (
    .clk(clk100m),
    .d(\PWM4/n31 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[19]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b2  (
    .clk(clk100m),
    .d(\PWM4/n31 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[2]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b20  (
    .clk(clk100m),
    .d(\PWM4/n31 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[20]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b21  (
    .clk(clk100m),
    .d(\PWM4/n31 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[21]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b22  (
    .clk(clk100m),
    .d(\PWM4/n31 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[22]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b23  (
    .clk(clk100m),
    .d(\PWM4/n31 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[23]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b3  (
    .clk(clk100m),
    .d(\PWM4/n31 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[3]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b4  (
    .clk(clk100m),
    .d(\PWM4/n31 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[4]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b5  (
    .clk(clk100m),
    .d(\PWM4/n31 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[5]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b6  (
    .clk(clk100m),
    .d(\PWM4/n31 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[6]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b7  (
    .clk(clk100m),
    .d(\PWM4/n31 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[7]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b8  (
    .clk(clk100m),
    .d(\PWM4/n31 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[8]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM4/reg3_b9  (
    .clk(clk100m),
    .d(\PWM4/n31 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM4/RemaTxNum[9]_keep ));  // src/OnePWM.v(58)
  reg_ar_ss_w1 \PWM4/stopreq_reg  (
    .clk(clk100m),
    .d(\PWM4/n1 ),
    .en(1'b1),
    .reset(1'b0),
    .set(pwm_start_stop[4]),
    .q(\PWM4/stopreq_keep ));  // src/OnePWM.v(15)
  add_pu27_mu27_o27 \PWM4/sub0  (
    .i0(\PWM4/FreCnt ),
    .i1(27'b000000000000000000000000001),
    .o(\PWM4/n12 [26:0]));  // src/OnePWM.v(32)
  add_pu24_mu24_o24 \PWM4/sub1  (
    .i0(pnumcnt4),
    .i1(24'b000000000000000000000001),
    .o(\PWM4/n26 [23:0]));  // src/OnePWM.v(55)
  AL_MUX \PWM4/u10  (
    .i0(1'b0),
    .i1(\PWM4/n9 ),
    .sel(n15),
    .o(\PWM4/n10 ));  // src/OnePWM.v(26)
  or \PWM4/u11  (\PWM4/n11 , pwm_state_read[4], pwm_start_stop[20]);  // src/OnePWM.v(30)
  and \PWM4/u14_sel_is_1  (\PWM4/u14_sel_is_1_o , pwm_state_read[4], \PWM4/n17_neg );
  and \PWM4/u15  (\PWM4/n24 , \PWM4/n0 , pwm_state_read[4]);  // src/OnePWM.v(54)
  and \PWM4/u17_sel_is_1  (\PWM4/u17_sel_is_1_o , \PWM4/n24 , \PWM4/n25_neg );
  not \PWM4/u17_sel_is_1_o_inv  (\PWM4/u17_sel_is_1_o_neg , \PWM4/u17_sel_is_1_o );
  AL_MUX \PWM4/u18  (
    .i0(\PWM4/pnumr [31]),
    .i1(dir[4]),
    .sel(\PWM4/u18_sel_is_0_o ),
    .o(\PWM4/n32 ));
  and \PWM4/u18_sel_is_0  (\PWM4/u18_sel_is_0_o , \pwm_start_stop[20]_neg , \PWM4/u17_sel_is_1_o_neg );
  AL_MUX \PWM4/u2  (
    .i0(\PWM4/stopreq ),
    .i1(1'b0),
    .sel(\PWM4/n0 ),
    .o(\PWM4/n1 ));  // src/OnePWM.v(15)
  and \PWM4/u5  (\PWM4/n4 , \PWM4/stopreq , \PWM4/n0 );  // src/OnePWM.v(23)
  and \PWM4/u6  (\PWM4/n6 , \PWM4/n5 , \PWM4/n0 );  // src/OnePWM.v(25)
  AL_MUX \PWM4/u8  (
    .i0(1'b0),
    .i1(pwm_state_read[4]),
    .sel(\PWM4/u8_sel_is_0_o ),
    .o(\PWM4/n8 ));
  and \PWM4/u8_sel_is_0  (\PWM4/u8_sel_is_0_o , \PWM4/n4_neg , \PWM4/n6_neg );
  AL_MUX \PWM4/u9  (
    .i0(\PWM4/n8 ),
    .i1(1'b1),
    .sel(pwm_start_stop[20]),
    .o(\PWM4/n9 ));  // src/OnePWM.v(26)
  reg_ar_as_w1 \PWM5/State_reg  (
    .clk(clk100m),
    .d(\PWM5/n10 ),
    .en(1'b1),
    .reset(~rstn),
    .set(1'b0),
    .q(pwm_state_read[5]));  // src/OnePWM.v(26)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[0]  (
    .i(\PWM5/RemaTxNum[0]_keep ),
    .o(pnumcnt5[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[10]  (
    .i(\PWM5/RemaTxNum[10]_keep ),
    .o(pnumcnt5[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[11]  (
    .i(\PWM5/RemaTxNum[11]_keep ),
    .o(pnumcnt5[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[12]  (
    .i(\PWM5/RemaTxNum[12]_keep ),
    .o(pnumcnt5[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[13]  (
    .i(\PWM5/RemaTxNum[13]_keep ),
    .o(pnumcnt5[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[14]  (
    .i(\PWM5/RemaTxNum[14]_keep ),
    .o(pnumcnt5[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[15]  (
    .i(\PWM5/RemaTxNum[15]_keep ),
    .o(pnumcnt5[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[16]  (
    .i(\PWM5/RemaTxNum[16]_keep ),
    .o(pnumcnt5[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[17]  (
    .i(\PWM5/RemaTxNum[17]_keep ),
    .o(pnumcnt5[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[18]  (
    .i(\PWM5/RemaTxNum[18]_keep ),
    .o(pnumcnt5[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[19]  (
    .i(\PWM5/RemaTxNum[19]_keep ),
    .o(pnumcnt5[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[1]  (
    .i(\PWM5/RemaTxNum[1]_keep ),
    .o(pnumcnt5[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[20]  (
    .i(\PWM5/RemaTxNum[20]_keep ),
    .o(pnumcnt5[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[21]  (
    .i(\PWM5/RemaTxNum[21]_keep ),
    .o(pnumcnt5[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[22]  (
    .i(\PWM5/RemaTxNum[22]_keep ),
    .o(pnumcnt5[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[23]  (
    .i(\PWM5/RemaTxNum[23]_keep ),
    .o(pnumcnt5[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[2]  (
    .i(\PWM5/RemaTxNum[2]_keep ),
    .o(pnumcnt5[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[3]  (
    .i(\PWM5/RemaTxNum[3]_keep ),
    .o(pnumcnt5[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[4]  (
    .i(\PWM5/RemaTxNum[4]_keep ),
    .o(pnumcnt5[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[5]  (
    .i(\PWM5/RemaTxNum[5]_keep ),
    .o(pnumcnt5[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[6]  (
    .i(\PWM5/RemaTxNum[6]_keep ),
    .o(pnumcnt5[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[7]  (
    .i(\PWM5/RemaTxNum[7]_keep ),
    .o(pnumcnt5[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[8]  (
    .i(\PWM5/RemaTxNum[8]_keep ),
    .o(pnumcnt5[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_RemaTxNum[9]  (
    .i(\PWM5/RemaTxNum[9]_keep ),
    .o(pnumcnt5[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_dir  (
    .i(\PWM5/dir_keep ),
    .o(dir[5]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[0]  (
    .i(\PWM5/pnumr[0]_keep ),
    .o(\PWM5/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[10]  (
    .i(\PWM5/pnumr[10]_keep ),
    .o(\PWM5/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[11]  (
    .i(\PWM5/pnumr[11]_keep ),
    .o(\PWM5/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[12]  (
    .i(\PWM5/pnumr[12]_keep ),
    .o(\PWM5/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[13]  (
    .i(\PWM5/pnumr[13]_keep ),
    .o(\PWM5/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[14]  (
    .i(\PWM5/pnumr[14]_keep ),
    .o(\PWM5/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[15]  (
    .i(\PWM5/pnumr[15]_keep ),
    .o(\PWM5/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[16]  (
    .i(\PWM5/pnumr[16]_keep ),
    .o(\PWM5/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[17]  (
    .i(\PWM5/pnumr[17]_keep ),
    .o(\PWM5/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[18]  (
    .i(\PWM5/pnumr[18]_keep ),
    .o(\PWM5/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[19]  (
    .i(\PWM5/pnumr[19]_keep ),
    .o(\PWM5/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[1]  (
    .i(\PWM5/pnumr[1]_keep ),
    .o(\PWM5/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[20]  (
    .i(\PWM5/pnumr[20]_keep ),
    .o(\PWM5/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[21]  (
    .i(\PWM5/pnumr[21]_keep ),
    .o(\PWM5/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[22]  (
    .i(\PWM5/pnumr[22]_keep ),
    .o(\PWM5/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[23]  (
    .i(\PWM5/pnumr[23]_keep ),
    .o(\PWM5/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[24]  (
    .i(\PWM5/pnumr[24]_keep ),
    .o(\PWM5/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[25]  (
    .i(\PWM5/pnumr[25]_keep ),
    .o(\PWM5/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[26]  (
    .i(\PWM5/pnumr[26]_keep ),
    .o(\PWM5/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[27]  (
    .i(\PWM5/pnumr[27]_keep ),
    .o(\PWM5/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[28]  (
    .i(\PWM5/pnumr[28]_keep ),
    .o(\PWM5/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[29]  (
    .i(\PWM5/pnumr[29]_keep ),
    .o(\PWM5/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[2]  (
    .i(\PWM5/pnumr[2]_keep ),
    .o(\PWM5/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[30]  (
    .i(\PWM5/pnumr[30]_keep ),
    .o(\PWM5/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[31]  (
    .i(\PWM5/pnumr[31]_keep ),
    .o(\PWM5/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[3]  (
    .i(\PWM5/pnumr[3]_keep ),
    .o(\PWM5/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[4]  (
    .i(\PWM5/pnumr[4]_keep ),
    .o(\PWM5/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[5]  (
    .i(\PWM5/pnumr[5]_keep ),
    .o(\PWM5/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[6]  (
    .i(\PWM5/pnumr[6]_keep ),
    .o(\PWM5/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[7]  (
    .i(\PWM5/pnumr[7]_keep ),
    .o(\PWM5/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[8]  (
    .i(\PWM5/pnumr[8]_keep ),
    .o(\PWM5/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pnumr[9]  (
    .i(\PWM5/pnumr[9]_keep ),
    .o(\PWM5/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_pwm  (
    .i(\PWM5/pwm_keep ),
    .o(pwm[5]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM5/_bufkeep_stopreq  (
    .i(\PWM5/stopreq_keep ),
    .o(\PWM5/stopreq ));  // src/OnePWM.v(14)
  reg_ar_as_w1 \PWM5/dir_reg  (
    .clk(clk100m),
    .d(\PWM5/n32 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/dir_keep ));  // src/OnePWM.v(58)
  eq_w27 \PWM5/eq0  (
    .i0(\PWM5/FreCnt ),
    .i1(27'b000000000000000000000000000),
    .o(\PWM5/n0 ));  // src/OnePWM.v(15)
  eq_w24 \PWM5/eq1  (
    .i0(pnumcnt5),
    .i1(24'b000000000000000000000001),
    .o(\PWM5/n5 ));  // src/OnePWM.v(25)
  eq_w27 \PWM5/eq2  (
    .i0(\PWM5/FreCnt ),
    .i1({1'b0,\PWM5/FreCntr [26:1]}),
    .o(\PWM5/n17 ));  // src/OnePWM.v(41)
  eq_w27 \PWM5/eq3  (
    .i0(\PWM5/FreCnt ),
    .i1(\PWM5/FreCntr ),
    .o(\PWM5/n18 ));  // src/OnePWM.v(43)
  binary_mux_s1_w1 \PWM5/mux0_b0  (
    .i0(\PWM5/n12 [0]),
    .i1(freq5[0]),
    .sel(\PWM5/n0 ),
    .o(\PWM5/n13 [0]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM5/mux0_b1  (
    .i0(\PWM5/n12 [1]),
    .i1(freq5[1]),
    .sel(\PWM5/n0 ),
    .o(\PWM5/n13 [1]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM5/mux0_b10  (
    .i0(\PWM5/n12 [10]),
    .i1(freq5[10]),
    .sel(\PWM5/n0 ),
    .o(\PWM5/n13 [10]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM5/mux0_b11  (
    .i0(\PWM5/n12 [11]),
    .i1(freq5[11]),
    .sel(\PWM5/n0 ),
    .o(\PWM5/n13 [11]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM5/mux0_b12  (
    .i0(\PWM5/n12 [12]),
    .i1(freq5[12]),
    .sel(\PWM5/n0 ),
    .o(\PWM5/n13 [12]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM5/mux0_b13  (
    .i0(\PWM5/n12 [13]),
    .i1(freq5[13]),
    .sel(\PWM5/n0 ),
    .o(\PWM5/n13 [13]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM5/mux0_b14  (
    .i0(\PWM5/n12 [14]),
    .i1(freq5[14]),
    .sel(\PWM5/n0 ),
    .o(\PWM5/n13 [14]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM5/mux0_b15  (
    .i0(\PWM5/n12 [15]),
    .i1(freq5[15]),
    .sel(\PWM5/n0 ),
    .o(\PWM5/n13 [15]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM5/mux0_b16  (
    .i0(\PWM5/n12 [16]),
    .i1(freq5[16]),
    .sel(\PWM5/n0 ),
    .o(\PWM5/n13 [16]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM5/mux0_b17  (
    .i0(\PWM5/n12 [17]),
    .i1(freq5[17]),
    .sel(\PWM5/n0 ),
    .o(\PWM5/n13 [17]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM5/mux0_b18  (
    .i0(\PWM5/n12 [18]),
    .i1(freq5[18]),
    .sel(\PWM5/n0 ),
    .o(\PWM5/n13 [18]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM5/mux0_b19  (
    .i0(\PWM5/n12 [19]),
    .i1(freq5[19]),
    .sel(\PWM5/n0 ),
    .o(\PWM5/n13 [19]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM5/mux0_b2  (
    .i0(\PWM5/n12 [2]),
    .i1(freq5[2]),
    .sel(\PWM5/n0 ),
    .o(\PWM5/n13 [2]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM5/mux0_b20  (
    .i0(\PWM5/n12 [20]),
    .i1(freq5[20]),
    .sel(\PWM5/n0 ),
    .o(\PWM5/n13 [20]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM5/mux0_b21  (
    .i0(\PWM5/n12 [21]),
    .i1(freq5[21]),
    .sel(\PWM5/n0 ),
    .o(\PWM5/n13 [21]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM5/mux0_b22  (
    .i0(\PWM5/n12 [22]),
    .i1(freq5[22]),
    .sel(\PWM5/n0 ),
    .o(\PWM5/n13 [22]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM5/mux0_b23  (
    .i0(\PWM5/n12 [23]),
    .i1(freq5[23]),
    .sel(\PWM5/n0 ),
    .o(\PWM5/n13 [23]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM5/mux0_b24  (
    .i0(\PWM5/n12 [24]),
    .i1(freq5[24]),
    .sel(\PWM5/n0 ),
    .o(\PWM5/n13 [24]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM5/mux0_b25  (
    .i0(\PWM5/n12 [25]),
    .i1(freq5[25]),
    .sel(\PWM5/n0 ),
    .o(\PWM5/n13 [25]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM5/mux0_b26  (
    .i0(\PWM5/n12 [26]),
    .i1(freq5[26]),
    .sel(\PWM5/n0 ),
    .o(\PWM5/n13 [26]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM5/mux0_b3  (
    .i0(\PWM5/n12 [3]),
    .i1(freq5[3]),
    .sel(\PWM5/n0 ),
    .o(\PWM5/n13 [3]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM5/mux0_b4  (
    .i0(\PWM5/n12 [4]),
    .i1(freq5[4]),
    .sel(\PWM5/n0 ),
    .o(\PWM5/n13 [4]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM5/mux0_b5  (
    .i0(\PWM5/n12 [5]),
    .i1(freq5[5]),
    .sel(\PWM5/n0 ),
    .o(\PWM5/n13 [5]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM5/mux0_b6  (
    .i0(\PWM5/n12 [6]),
    .i1(freq5[6]),
    .sel(\PWM5/n0 ),
    .o(\PWM5/n13 [6]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM5/mux0_b7  (
    .i0(\PWM5/n12 [7]),
    .i1(freq5[7]),
    .sel(\PWM5/n0 ),
    .o(\PWM5/n13 [7]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM5/mux0_b8  (
    .i0(\PWM5/n12 [8]),
    .i1(freq5[8]),
    .sel(\PWM5/n0 ),
    .o(\PWM5/n13 [8]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM5/mux0_b9  (
    .i0(\PWM5/n12 [9]),
    .i1(freq5[9]),
    .sel(\PWM5/n0 ),
    .o(\PWM5/n13 [9]));  // src/OnePWM.v(32)
  and \PWM5/mux3_b0_sel_is_3  (\PWM5/mux3_b0_sel_is_3_o , \PWM5/n11 , \PWM5/n0 );
  binary_mux_s1_w1 \PWM5/mux4_b0  (
    .i0(\PWM5/pnumr [0]),
    .i1(1'b0),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n22 [0]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux4_b1  (
    .i0(\PWM5/pnumr [1]),
    .i1(1'b0),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n22 [1]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux4_b10  (
    .i0(\PWM5/pnumr [10]),
    .i1(1'b0),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n22 [10]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux4_b11  (
    .i0(\PWM5/pnumr [11]),
    .i1(1'b0),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n22 [11]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux4_b12  (
    .i0(\PWM5/pnumr [12]),
    .i1(1'b0),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n22 [12]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux4_b13  (
    .i0(\PWM5/pnumr [13]),
    .i1(1'b0),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n22 [13]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux4_b14  (
    .i0(\PWM5/pnumr [14]),
    .i1(1'b0),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n22 [14]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux4_b15  (
    .i0(\PWM5/pnumr [15]),
    .i1(1'b0),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n22 [15]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux4_b16  (
    .i0(\PWM5/pnumr [16]),
    .i1(1'b0),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n22 [16]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux4_b17  (
    .i0(\PWM5/pnumr [17]),
    .i1(1'b0),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n22 [17]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux4_b18  (
    .i0(\PWM5/pnumr [18]),
    .i1(1'b0),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n22 [18]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux4_b19  (
    .i0(\PWM5/pnumr [19]),
    .i1(1'b0),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n22 [19]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux4_b2  (
    .i0(\PWM5/pnumr [2]),
    .i1(1'b0),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n22 [2]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux4_b20  (
    .i0(\PWM5/pnumr [20]),
    .i1(1'b0),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n22 [20]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux4_b21  (
    .i0(\PWM5/pnumr [21]),
    .i1(1'b0),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n22 [21]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux4_b22  (
    .i0(\PWM5/pnumr [22]),
    .i1(1'b0),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n22 [22]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux4_b23  (
    .i0(\PWM5/pnumr [23]),
    .i1(1'b0),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n22 [23]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux4_b24  (
    .i0(\PWM5/pnumr [24]),
    .i1(1'b0),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n22 [24]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux4_b25  (
    .i0(\PWM5/pnumr [25]),
    .i1(1'b0),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n22 [25]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux4_b26  (
    .i0(\PWM5/pnumr [26]),
    .i1(1'b0),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n22 [26]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux4_b27  (
    .i0(\PWM5/pnumr [27]),
    .i1(1'b0),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n22 [27]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux4_b28  (
    .i0(\PWM5/pnumr [28]),
    .i1(1'b0),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n22 [28]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux4_b29  (
    .i0(\PWM5/pnumr [29]),
    .i1(1'b0),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n22 [29]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux4_b3  (
    .i0(\PWM5/pnumr [3]),
    .i1(1'b0),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n22 [3]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux4_b30  (
    .i0(\PWM5/pnumr [30]),
    .i1(1'b0),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n22 [30]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux4_b31  (
    .i0(\PWM5/pnumr [31]),
    .i1(1'b0),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n22 [31]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux4_b4  (
    .i0(\PWM5/pnumr [4]),
    .i1(1'b0),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n22 [4]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux4_b5  (
    .i0(\PWM5/pnumr [5]),
    .i1(1'b0),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n22 [5]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux4_b6  (
    .i0(\PWM5/pnumr [6]),
    .i1(1'b0),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n22 [6]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux4_b7  (
    .i0(\PWM5/pnumr [7]),
    .i1(1'b0),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n22 [7]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux4_b8  (
    .i0(\PWM5/pnumr [8]),
    .i1(1'b0),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n22 [8]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux4_b9  (
    .i0(\PWM5/pnumr [9]),
    .i1(1'b0),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n22 [9]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux5_b0  (
    .i0(\PWM5/n22 [0]),
    .i1(pnum5[0]),
    .sel(pnum5[32]),
    .o(\PWM5/n23 [0]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux5_b1  (
    .i0(\PWM5/n22 [1]),
    .i1(pnum5[1]),
    .sel(pnum5[32]),
    .o(\PWM5/n23 [1]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux5_b10  (
    .i0(\PWM5/n22 [10]),
    .i1(pnum5[10]),
    .sel(pnum5[32]),
    .o(\PWM5/n23 [10]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux5_b11  (
    .i0(\PWM5/n22 [11]),
    .i1(pnum5[11]),
    .sel(pnum5[32]),
    .o(\PWM5/n23 [11]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux5_b12  (
    .i0(\PWM5/n22 [12]),
    .i1(pnum5[12]),
    .sel(pnum5[32]),
    .o(\PWM5/n23 [12]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux5_b13  (
    .i0(\PWM5/n22 [13]),
    .i1(pnum5[13]),
    .sel(pnum5[32]),
    .o(\PWM5/n23 [13]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux5_b14  (
    .i0(\PWM5/n22 [14]),
    .i1(pnum5[14]),
    .sel(pnum5[32]),
    .o(\PWM5/n23 [14]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux5_b15  (
    .i0(\PWM5/n22 [15]),
    .i1(pnum5[15]),
    .sel(pnum5[32]),
    .o(\PWM5/n23 [15]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux5_b16  (
    .i0(\PWM5/n22 [16]),
    .i1(pnum5[16]),
    .sel(pnum5[32]),
    .o(\PWM5/n23 [16]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux5_b17  (
    .i0(\PWM5/n22 [17]),
    .i1(pnum5[17]),
    .sel(pnum5[32]),
    .o(\PWM5/n23 [17]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux5_b18  (
    .i0(\PWM5/n22 [18]),
    .i1(pnum5[18]),
    .sel(pnum5[32]),
    .o(\PWM5/n23 [18]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux5_b19  (
    .i0(\PWM5/n22 [19]),
    .i1(pnum5[19]),
    .sel(pnum5[32]),
    .o(\PWM5/n23 [19]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux5_b2  (
    .i0(\PWM5/n22 [2]),
    .i1(pnum5[2]),
    .sel(pnum5[32]),
    .o(\PWM5/n23 [2]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux5_b20  (
    .i0(\PWM5/n22 [20]),
    .i1(pnum5[20]),
    .sel(pnum5[32]),
    .o(\PWM5/n23 [20]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux5_b21  (
    .i0(\PWM5/n22 [21]),
    .i1(pnum5[21]),
    .sel(pnum5[32]),
    .o(\PWM5/n23 [21]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux5_b22  (
    .i0(\PWM5/n22 [22]),
    .i1(pnum5[22]),
    .sel(pnum5[32]),
    .o(\PWM5/n23 [22]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux5_b23  (
    .i0(\PWM5/n22 [23]),
    .i1(pnum5[23]),
    .sel(pnum5[32]),
    .o(\PWM5/n23 [23]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux5_b24  (
    .i0(\PWM5/n22 [24]),
    .i1(pnum5[24]),
    .sel(pnum5[32]),
    .o(\PWM5/n23 [24]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux5_b25  (
    .i0(\PWM5/n22 [25]),
    .i1(pnum5[25]),
    .sel(pnum5[32]),
    .o(\PWM5/n23 [25]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux5_b26  (
    .i0(\PWM5/n22 [26]),
    .i1(pnum5[26]),
    .sel(pnum5[32]),
    .o(\PWM5/n23 [26]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux5_b27  (
    .i0(\PWM5/n22 [27]),
    .i1(pnum5[27]),
    .sel(pnum5[32]),
    .o(\PWM5/n23 [27]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux5_b28  (
    .i0(\PWM5/n22 [28]),
    .i1(pnum5[28]),
    .sel(pnum5[32]),
    .o(\PWM5/n23 [28]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux5_b29  (
    .i0(\PWM5/n22 [29]),
    .i1(pnum5[29]),
    .sel(pnum5[32]),
    .o(\PWM5/n23 [29]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux5_b3  (
    .i0(\PWM5/n22 [3]),
    .i1(pnum5[3]),
    .sel(pnum5[32]),
    .o(\PWM5/n23 [3]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux5_b30  (
    .i0(\PWM5/n22 [30]),
    .i1(pnum5[30]),
    .sel(pnum5[32]),
    .o(\PWM5/n23 [30]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux5_b31  (
    .i0(\PWM5/n22 [31]),
    .i1(pnum5[31]),
    .sel(pnum5[32]),
    .o(\PWM5/n23 [31]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux5_b4  (
    .i0(\PWM5/n22 [4]),
    .i1(pnum5[4]),
    .sel(pnum5[32]),
    .o(\PWM5/n23 [4]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux5_b5  (
    .i0(\PWM5/n22 [5]),
    .i1(pnum5[5]),
    .sel(pnum5[32]),
    .o(\PWM5/n23 [5]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux5_b6  (
    .i0(\PWM5/n22 [6]),
    .i1(pnum5[6]),
    .sel(pnum5[32]),
    .o(\PWM5/n23 [6]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux5_b7  (
    .i0(\PWM5/n22 [7]),
    .i1(pnum5[7]),
    .sel(pnum5[32]),
    .o(\PWM5/n23 [7]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux5_b8  (
    .i0(\PWM5/n22 [8]),
    .i1(pnum5[8]),
    .sel(pnum5[32]),
    .o(\PWM5/n23 [8]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux5_b9  (
    .i0(\PWM5/n22 [9]),
    .i1(pnum5[9]),
    .sel(pnum5[32]),
    .o(\PWM5/n23 [9]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM5/mux6_b0  (
    .i0(\PWM5/pnumr [0]),
    .i1(\PWM5/n26 [0]),
    .sel(\PWM5/n25 ),
    .o(\PWM5/n27 [0]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM5/mux6_b1  (
    .i0(\PWM5/pnumr [1]),
    .i1(\PWM5/n26 [1]),
    .sel(\PWM5/n25 ),
    .o(\PWM5/n27 [1]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM5/mux6_b10  (
    .i0(\PWM5/pnumr [10]),
    .i1(\PWM5/n26 [10]),
    .sel(\PWM5/n25 ),
    .o(\PWM5/n27 [10]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM5/mux6_b11  (
    .i0(\PWM5/pnumr [11]),
    .i1(\PWM5/n26 [11]),
    .sel(\PWM5/n25 ),
    .o(\PWM5/n27 [11]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM5/mux6_b12  (
    .i0(\PWM5/pnumr [12]),
    .i1(\PWM5/n26 [12]),
    .sel(\PWM5/n25 ),
    .o(\PWM5/n27 [12]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM5/mux6_b13  (
    .i0(\PWM5/pnumr [13]),
    .i1(\PWM5/n26 [13]),
    .sel(\PWM5/n25 ),
    .o(\PWM5/n27 [13]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM5/mux6_b14  (
    .i0(\PWM5/pnumr [14]),
    .i1(\PWM5/n26 [14]),
    .sel(\PWM5/n25 ),
    .o(\PWM5/n27 [14]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM5/mux6_b15  (
    .i0(\PWM5/pnumr [15]),
    .i1(\PWM5/n26 [15]),
    .sel(\PWM5/n25 ),
    .o(\PWM5/n27 [15]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM5/mux6_b16  (
    .i0(\PWM5/pnumr [16]),
    .i1(\PWM5/n26 [16]),
    .sel(\PWM5/n25 ),
    .o(\PWM5/n27 [16]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM5/mux6_b17  (
    .i0(\PWM5/pnumr [17]),
    .i1(\PWM5/n26 [17]),
    .sel(\PWM5/n25 ),
    .o(\PWM5/n27 [17]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM5/mux6_b18  (
    .i0(\PWM5/pnumr [18]),
    .i1(\PWM5/n26 [18]),
    .sel(\PWM5/n25 ),
    .o(\PWM5/n27 [18]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM5/mux6_b19  (
    .i0(\PWM5/pnumr [19]),
    .i1(\PWM5/n26 [19]),
    .sel(\PWM5/n25 ),
    .o(\PWM5/n27 [19]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM5/mux6_b2  (
    .i0(\PWM5/pnumr [2]),
    .i1(\PWM5/n26 [2]),
    .sel(\PWM5/n25 ),
    .o(\PWM5/n27 [2]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM5/mux6_b20  (
    .i0(\PWM5/pnumr [20]),
    .i1(\PWM5/n26 [20]),
    .sel(\PWM5/n25 ),
    .o(\PWM5/n27 [20]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM5/mux6_b21  (
    .i0(\PWM5/pnumr [21]),
    .i1(\PWM5/n26 [21]),
    .sel(\PWM5/n25 ),
    .o(\PWM5/n27 [21]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM5/mux6_b22  (
    .i0(\PWM5/pnumr [22]),
    .i1(\PWM5/n26 [22]),
    .sel(\PWM5/n25 ),
    .o(\PWM5/n27 [22]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM5/mux6_b23  (
    .i0(\PWM5/pnumr [23]),
    .i1(\PWM5/n26 [23]),
    .sel(\PWM5/n25 ),
    .o(\PWM5/n27 [23]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM5/mux6_b3  (
    .i0(\PWM5/pnumr [3]),
    .i1(\PWM5/n26 [3]),
    .sel(\PWM5/n25 ),
    .o(\PWM5/n27 [3]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM5/mux6_b4  (
    .i0(\PWM5/pnumr [4]),
    .i1(\PWM5/n26 [4]),
    .sel(\PWM5/n25 ),
    .o(\PWM5/n27 [4]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM5/mux6_b5  (
    .i0(\PWM5/pnumr [5]),
    .i1(\PWM5/n26 [5]),
    .sel(\PWM5/n25 ),
    .o(\PWM5/n27 [5]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM5/mux6_b6  (
    .i0(\PWM5/pnumr [6]),
    .i1(\PWM5/n26 [6]),
    .sel(\PWM5/n25 ),
    .o(\PWM5/n27 [6]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM5/mux6_b7  (
    .i0(\PWM5/pnumr [7]),
    .i1(\PWM5/n26 [7]),
    .sel(\PWM5/n25 ),
    .o(\PWM5/n27 [7]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM5/mux6_b8  (
    .i0(\PWM5/pnumr [8]),
    .i1(\PWM5/n26 [8]),
    .sel(\PWM5/n25 ),
    .o(\PWM5/n27 [8]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM5/mux6_b9  (
    .i0(\PWM5/pnumr [9]),
    .i1(\PWM5/n26 [9]),
    .sel(\PWM5/n25 ),
    .o(\PWM5/n27 [9]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM5/mux7_b0  (
    .i0(pnumcnt5[0]),
    .i1(\PWM5/n27 [0]),
    .sel(\PWM5/n24 ),
    .o(\PWM5/n29 [0]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux7_b1  (
    .i0(pnumcnt5[1]),
    .i1(\PWM5/n27 [1]),
    .sel(\PWM5/n24 ),
    .o(\PWM5/n29 [1]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux7_b10  (
    .i0(pnumcnt5[10]),
    .i1(\PWM5/n27 [10]),
    .sel(\PWM5/n24 ),
    .o(\PWM5/n29 [10]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux7_b11  (
    .i0(pnumcnt5[11]),
    .i1(\PWM5/n27 [11]),
    .sel(\PWM5/n24 ),
    .o(\PWM5/n29 [11]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux7_b12  (
    .i0(pnumcnt5[12]),
    .i1(\PWM5/n27 [12]),
    .sel(\PWM5/n24 ),
    .o(\PWM5/n29 [12]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux7_b13  (
    .i0(pnumcnt5[13]),
    .i1(\PWM5/n27 [13]),
    .sel(\PWM5/n24 ),
    .o(\PWM5/n29 [13]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux7_b14  (
    .i0(pnumcnt5[14]),
    .i1(\PWM5/n27 [14]),
    .sel(\PWM5/n24 ),
    .o(\PWM5/n29 [14]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux7_b15  (
    .i0(pnumcnt5[15]),
    .i1(\PWM5/n27 [15]),
    .sel(\PWM5/n24 ),
    .o(\PWM5/n29 [15]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux7_b16  (
    .i0(pnumcnt5[16]),
    .i1(\PWM5/n27 [16]),
    .sel(\PWM5/n24 ),
    .o(\PWM5/n29 [16]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux7_b17  (
    .i0(pnumcnt5[17]),
    .i1(\PWM5/n27 [17]),
    .sel(\PWM5/n24 ),
    .o(\PWM5/n29 [17]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux7_b18  (
    .i0(pnumcnt5[18]),
    .i1(\PWM5/n27 [18]),
    .sel(\PWM5/n24 ),
    .o(\PWM5/n29 [18]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux7_b19  (
    .i0(pnumcnt5[19]),
    .i1(\PWM5/n27 [19]),
    .sel(\PWM5/n24 ),
    .o(\PWM5/n29 [19]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux7_b2  (
    .i0(pnumcnt5[2]),
    .i1(\PWM5/n27 [2]),
    .sel(\PWM5/n24 ),
    .o(\PWM5/n29 [2]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux7_b20  (
    .i0(pnumcnt5[20]),
    .i1(\PWM5/n27 [20]),
    .sel(\PWM5/n24 ),
    .o(\PWM5/n29 [20]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux7_b21  (
    .i0(pnumcnt5[21]),
    .i1(\PWM5/n27 [21]),
    .sel(\PWM5/n24 ),
    .o(\PWM5/n29 [21]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux7_b22  (
    .i0(pnumcnt5[22]),
    .i1(\PWM5/n27 [22]),
    .sel(\PWM5/n24 ),
    .o(\PWM5/n29 [22]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux7_b23  (
    .i0(pnumcnt5[23]),
    .i1(\PWM5/n27 [23]),
    .sel(\PWM5/n24 ),
    .o(\PWM5/n29 [23]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux7_b3  (
    .i0(pnumcnt5[3]),
    .i1(\PWM5/n27 [3]),
    .sel(\PWM5/n24 ),
    .o(\PWM5/n29 [3]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux7_b4  (
    .i0(pnumcnt5[4]),
    .i1(\PWM5/n27 [4]),
    .sel(\PWM5/n24 ),
    .o(\PWM5/n29 [4]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux7_b5  (
    .i0(pnumcnt5[5]),
    .i1(\PWM5/n27 [5]),
    .sel(\PWM5/n24 ),
    .o(\PWM5/n29 [5]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux7_b6  (
    .i0(pnumcnt5[6]),
    .i1(\PWM5/n27 [6]),
    .sel(\PWM5/n24 ),
    .o(\PWM5/n29 [6]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux7_b7  (
    .i0(pnumcnt5[7]),
    .i1(\PWM5/n27 [7]),
    .sel(\PWM5/n24 ),
    .o(\PWM5/n29 [7]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux7_b8  (
    .i0(pnumcnt5[8]),
    .i1(\PWM5/n27 [8]),
    .sel(\PWM5/n24 ),
    .o(\PWM5/n29 [8]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux7_b9  (
    .i0(pnumcnt5[9]),
    .i1(\PWM5/n27 [9]),
    .sel(\PWM5/n24 ),
    .o(\PWM5/n29 [9]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux8_b0  (
    .i0(\PWM5/n29 [0]),
    .i1(\PWM5/pnumr [0]),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n31 [0]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux8_b1  (
    .i0(\PWM5/n29 [1]),
    .i1(\PWM5/pnumr [1]),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n31 [1]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux8_b10  (
    .i0(\PWM5/n29 [10]),
    .i1(\PWM5/pnumr [10]),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n31 [10]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux8_b11  (
    .i0(\PWM5/n29 [11]),
    .i1(\PWM5/pnumr [11]),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n31 [11]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux8_b12  (
    .i0(\PWM5/n29 [12]),
    .i1(\PWM5/pnumr [12]),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n31 [12]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux8_b13  (
    .i0(\PWM5/n29 [13]),
    .i1(\PWM5/pnumr [13]),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n31 [13]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux8_b14  (
    .i0(\PWM5/n29 [14]),
    .i1(\PWM5/pnumr [14]),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n31 [14]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux8_b15  (
    .i0(\PWM5/n29 [15]),
    .i1(\PWM5/pnumr [15]),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n31 [15]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux8_b16  (
    .i0(\PWM5/n29 [16]),
    .i1(\PWM5/pnumr [16]),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n31 [16]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux8_b17  (
    .i0(\PWM5/n29 [17]),
    .i1(\PWM5/pnumr [17]),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n31 [17]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux8_b18  (
    .i0(\PWM5/n29 [18]),
    .i1(\PWM5/pnumr [18]),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n31 [18]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux8_b19  (
    .i0(\PWM5/n29 [19]),
    .i1(\PWM5/pnumr [19]),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n31 [19]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux8_b2  (
    .i0(\PWM5/n29 [2]),
    .i1(\PWM5/pnumr [2]),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n31 [2]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux8_b20  (
    .i0(\PWM5/n29 [20]),
    .i1(\PWM5/pnumr [20]),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n31 [20]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux8_b21  (
    .i0(\PWM5/n29 [21]),
    .i1(\PWM5/pnumr [21]),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n31 [21]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux8_b22  (
    .i0(\PWM5/n29 [22]),
    .i1(\PWM5/pnumr [22]),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n31 [22]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux8_b23  (
    .i0(\PWM5/n29 [23]),
    .i1(\PWM5/pnumr [23]),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n31 [23]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux8_b3  (
    .i0(\PWM5/n29 [3]),
    .i1(\PWM5/pnumr [3]),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n31 [3]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux8_b4  (
    .i0(\PWM5/n29 [4]),
    .i1(\PWM5/pnumr [4]),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n31 [4]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux8_b5  (
    .i0(\PWM5/n29 [5]),
    .i1(\PWM5/pnumr [5]),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n31 [5]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux8_b6  (
    .i0(\PWM5/n29 [6]),
    .i1(\PWM5/pnumr [6]),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n31 [6]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux8_b7  (
    .i0(\PWM5/n29 [7]),
    .i1(\PWM5/pnumr [7]),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n31 [7]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux8_b8  (
    .i0(\PWM5/n29 [8]),
    .i1(\PWM5/pnumr [8]),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n31 [8]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM5/mux8_b9  (
    .i0(\PWM5/n29 [9]),
    .i1(\PWM5/pnumr [9]),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n31 [9]));  // src/OnePWM.v(57)
  not \PWM5/n17_inv  (\PWM5/n17_neg , \PWM5/n17 );
  not \PWM5/n25_inv  (\PWM5/n25_neg , \PWM5/n25 );
  not \PWM5/n4_inv  (\PWM5/n4_neg , \PWM5/n4 );
  not \PWM5/n6_inv  (\PWM5/n6_neg , \PWM5/n6 );
  ne_w24 \PWM5/neq0  (
    .i0(pnumcnt5),
    .i1(24'b000000000000000000000000),
    .o(\PWM5/n25 ));  // src/OnePWM.v(55)
  reg_sr_ss_w1 \PWM5/pwm_reg  (
    .clk(clk100m),
    .d(pwm[5]),
    .en(1'b1),
    .reset(~\PWM5/u14_sel_is_1_o ),
    .set(\PWM5/n18 ),
    .q(\PWM5/pwm_keep ));  // src/OnePWM.v(45)
  reg_sr_as_w1 \PWM5/reg0_b0  (
    .clk(clk100m),
    .d(\PWM5/n13 [0]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [0]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b1  (
    .clk(clk100m),
    .d(\PWM5/n13 [1]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [1]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b10  (
    .clk(clk100m),
    .d(\PWM5/n13 [10]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [10]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b11  (
    .clk(clk100m),
    .d(\PWM5/n13 [11]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [11]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b12  (
    .clk(clk100m),
    .d(\PWM5/n13 [12]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [12]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b13  (
    .clk(clk100m),
    .d(\PWM5/n13 [13]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [13]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b14  (
    .clk(clk100m),
    .d(\PWM5/n13 [14]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [14]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b15  (
    .clk(clk100m),
    .d(\PWM5/n13 [15]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [15]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b16  (
    .clk(clk100m),
    .d(\PWM5/n13 [16]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [16]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b17  (
    .clk(clk100m),
    .d(\PWM5/n13 [17]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [17]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b18  (
    .clk(clk100m),
    .d(\PWM5/n13 [18]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [18]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b19  (
    .clk(clk100m),
    .d(\PWM5/n13 [19]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [19]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b2  (
    .clk(clk100m),
    .d(\PWM5/n13 [2]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [2]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b20  (
    .clk(clk100m),
    .d(\PWM5/n13 [20]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [20]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b21  (
    .clk(clk100m),
    .d(\PWM5/n13 [21]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [21]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b22  (
    .clk(clk100m),
    .d(\PWM5/n13 [22]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [22]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b23  (
    .clk(clk100m),
    .d(\PWM5/n13 [23]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [23]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b24  (
    .clk(clk100m),
    .d(\PWM5/n13 [24]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [24]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b25  (
    .clk(clk100m),
    .d(\PWM5/n13 [25]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [25]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b26  (
    .clk(clk100m),
    .d(\PWM5/n13 [26]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [26]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b3  (
    .clk(clk100m),
    .d(\PWM5/n13 [3]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [3]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b4  (
    .clk(clk100m),
    .d(\PWM5/n13 [4]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [4]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b5  (
    .clk(clk100m),
    .d(\PWM5/n13 [5]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [5]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b6  (
    .clk(clk100m),
    .d(\PWM5/n13 [6]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [6]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b7  (
    .clk(clk100m),
    .d(\PWM5/n13 [7]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [7]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b8  (
    .clk(clk100m),
    .d(\PWM5/n13 [8]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [8]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM5/reg0_b9  (
    .clk(clk100m),
    .d(\PWM5/n13 [9]),
    .en(1'b1),
    .reset(~\PWM5/n11 ),
    .set(1'b0),
    .q(\PWM5/FreCnt [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b0  (
    .clk(clk100m),
    .d(freq5[0]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [0]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b1  (
    .clk(clk100m),
    .d(freq5[1]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [1]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b10  (
    .clk(clk100m),
    .d(freq5[10]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [10]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b11  (
    .clk(clk100m),
    .d(freq5[11]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [11]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b12  (
    .clk(clk100m),
    .d(freq5[12]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [12]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b13  (
    .clk(clk100m),
    .d(freq5[13]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [13]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b14  (
    .clk(clk100m),
    .d(freq5[14]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [14]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b15  (
    .clk(clk100m),
    .d(freq5[15]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [15]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b16  (
    .clk(clk100m),
    .d(freq5[16]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [16]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b17  (
    .clk(clk100m),
    .d(freq5[17]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [17]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b18  (
    .clk(clk100m),
    .d(freq5[18]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [18]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b19  (
    .clk(clk100m),
    .d(freq5[19]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [19]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b2  (
    .clk(clk100m),
    .d(freq5[2]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [2]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b20  (
    .clk(clk100m),
    .d(freq5[20]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [20]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b21  (
    .clk(clk100m),
    .d(freq5[21]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [21]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b22  (
    .clk(clk100m),
    .d(freq5[22]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [22]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b23  (
    .clk(clk100m),
    .d(freq5[23]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [23]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b24  (
    .clk(clk100m),
    .d(freq5[24]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [24]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b25  (
    .clk(clk100m),
    .d(freq5[25]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [25]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b26  (
    .clk(clk100m),
    .d(freq5[26]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [26]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b3  (
    .clk(clk100m),
    .d(freq5[3]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [3]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b4  (
    .clk(clk100m),
    .d(freq5[4]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [4]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b5  (
    .clk(clk100m),
    .d(freq5[5]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [5]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b6  (
    .clk(clk100m),
    .d(freq5[6]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [6]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b7  (
    .clk(clk100m),
    .d(freq5[7]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [7]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b8  (
    .clk(clk100m),
    .d(freq5[8]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [8]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg1_b9  (
    .clk(clk100m),
    .d(freq5[9]),
    .en(\PWM5/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/FreCntr [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM5/reg2_b0  (
    .clk(clk100m),
    .d(\PWM5/n23 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[0]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b1  (
    .clk(clk100m),
    .d(\PWM5/n23 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[1]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b10  (
    .clk(clk100m),
    .d(\PWM5/n23 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[10]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b11  (
    .clk(clk100m),
    .d(\PWM5/n23 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[11]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b12  (
    .clk(clk100m),
    .d(\PWM5/n23 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[12]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b13  (
    .clk(clk100m),
    .d(\PWM5/n23 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[13]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b14  (
    .clk(clk100m),
    .d(\PWM5/n23 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[14]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b15  (
    .clk(clk100m),
    .d(\PWM5/n23 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[15]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b16  (
    .clk(clk100m),
    .d(\PWM5/n23 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[16]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b17  (
    .clk(clk100m),
    .d(\PWM5/n23 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[17]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b18  (
    .clk(clk100m),
    .d(\PWM5/n23 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[18]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b19  (
    .clk(clk100m),
    .d(\PWM5/n23 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[19]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b2  (
    .clk(clk100m),
    .d(\PWM5/n23 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[2]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b20  (
    .clk(clk100m),
    .d(\PWM5/n23 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[20]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b21  (
    .clk(clk100m),
    .d(\PWM5/n23 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[21]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b22  (
    .clk(clk100m),
    .d(\PWM5/n23 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[22]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b23  (
    .clk(clk100m),
    .d(\PWM5/n23 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[23]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b24  (
    .clk(clk100m),
    .d(\PWM5/n23 [24]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[24]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b25  (
    .clk(clk100m),
    .d(\PWM5/n23 [25]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[25]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b26  (
    .clk(clk100m),
    .d(\PWM5/n23 [26]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[26]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b27  (
    .clk(clk100m),
    .d(\PWM5/n23 [27]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[27]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b28  (
    .clk(clk100m),
    .d(\PWM5/n23 [28]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[28]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b29  (
    .clk(clk100m),
    .d(\PWM5/n23 [29]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[29]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b3  (
    .clk(clk100m),
    .d(\PWM5/n23 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[3]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b30  (
    .clk(clk100m),
    .d(\PWM5/n23 [30]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[30]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b31  (
    .clk(clk100m),
    .d(\PWM5/n23 [31]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[31]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b4  (
    .clk(clk100m),
    .d(\PWM5/n23 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[4]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b5  (
    .clk(clk100m),
    .d(\PWM5/n23 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[5]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b6  (
    .clk(clk100m),
    .d(\PWM5/n23 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[6]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b7  (
    .clk(clk100m),
    .d(\PWM5/n23 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[7]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b8  (
    .clk(clk100m),
    .d(\PWM5/n23 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[8]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg2_b9  (
    .clk(clk100m),
    .d(\PWM5/n23 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/pnumr[9]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM5/reg3_b0  (
    .clk(clk100m),
    .d(\PWM5/n31 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[0]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b1  (
    .clk(clk100m),
    .d(\PWM5/n31 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[1]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b10  (
    .clk(clk100m),
    .d(\PWM5/n31 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[10]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b11  (
    .clk(clk100m),
    .d(\PWM5/n31 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[11]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b12  (
    .clk(clk100m),
    .d(\PWM5/n31 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[12]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b13  (
    .clk(clk100m),
    .d(\PWM5/n31 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[13]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b14  (
    .clk(clk100m),
    .d(\PWM5/n31 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[14]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b15  (
    .clk(clk100m),
    .d(\PWM5/n31 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[15]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b16  (
    .clk(clk100m),
    .d(\PWM5/n31 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[16]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b17  (
    .clk(clk100m),
    .d(\PWM5/n31 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[17]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b18  (
    .clk(clk100m),
    .d(\PWM5/n31 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[18]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b19  (
    .clk(clk100m),
    .d(\PWM5/n31 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[19]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b2  (
    .clk(clk100m),
    .d(\PWM5/n31 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[2]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b20  (
    .clk(clk100m),
    .d(\PWM5/n31 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[20]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b21  (
    .clk(clk100m),
    .d(\PWM5/n31 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[21]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b22  (
    .clk(clk100m),
    .d(\PWM5/n31 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[22]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b23  (
    .clk(clk100m),
    .d(\PWM5/n31 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[23]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b3  (
    .clk(clk100m),
    .d(\PWM5/n31 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[3]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b4  (
    .clk(clk100m),
    .d(\PWM5/n31 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[4]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b5  (
    .clk(clk100m),
    .d(\PWM5/n31 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[5]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b6  (
    .clk(clk100m),
    .d(\PWM5/n31 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[6]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b7  (
    .clk(clk100m),
    .d(\PWM5/n31 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[7]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b8  (
    .clk(clk100m),
    .d(\PWM5/n31 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[8]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM5/reg3_b9  (
    .clk(clk100m),
    .d(\PWM5/n31 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM5/RemaTxNum[9]_keep ));  // src/OnePWM.v(58)
  reg_ar_ss_w1 \PWM5/stopreq_reg  (
    .clk(clk100m),
    .d(\PWM5/n1 ),
    .en(1'b1),
    .reset(1'b0),
    .set(pwm_start_stop[5]),
    .q(\PWM5/stopreq_keep ));  // src/OnePWM.v(15)
  add_pu27_mu27_o27 \PWM5/sub0  (
    .i0(\PWM5/FreCnt ),
    .i1(27'b000000000000000000000000001),
    .o(\PWM5/n12 [26:0]));  // src/OnePWM.v(32)
  add_pu24_mu24_o24 \PWM5/sub1  (
    .i0(pnumcnt5),
    .i1(24'b000000000000000000000001),
    .o(\PWM5/n26 [23:0]));  // src/OnePWM.v(55)
  AL_MUX \PWM5/u10  (
    .i0(1'b0),
    .i1(\PWM5/n9 ),
    .sel(n16),
    .o(\PWM5/n10 ));  // src/OnePWM.v(26)
  or \PWM5/u11  (\PWM5/n11 , pwm_state_read[5], pwm_start_stop[21]);  // src/OnePWM.v(30)
  and \PWM5/u14_sel_is_1  (\PWM5/u14_sel_is_1_o , pwm_state_read[5], \PWM5/n17_neg );
  and \PWM5/u15  (\PWM5/n24 , \PWM5/n0 , pwm_state_read[5]);  // src/OnePWM.v(54)
  and \PWM5/u17_sel_is_1  (\PWM5/u17_sel_is_1_o , \PWM5/n24 , \PWM5/n25_neg );
  not \PWM5/u17_sel_is_1_o_inv  (\PWM5/u17_sel_is_1_o_neg , \PWM5/u17_sel_is_1_o );
  AL_MUX \PWM5/u18  (
    .i0(\PWM5/pnumr [31]),
    .i1(dir[5]),
    .sel(\PWM5/u18_sel_is_0_o ),
    .o(\PWM5/n32 ));
  and \PWM5/u18_sel_is_0  (\PWM5/u18_sel_is_0_o , \pwm_start_stop[21]_neg , \PWM5/u17_sel_is_1_o_neg );
  AL_MUX \PWM5/u2  (
    .i0(\PWM5/stopreq ),
    .i1(1'b0),
    .sel(\PWM5/n0 ),
    .o(\PWM5/n1 ));  // src/OnePWM.v(15)
  and \PWM5/u5  (\PWM5/n4 , \PWM5/stopreq , \PWM5/n0 );  // src/OnePWM.v(23)
  and \PWM5/u6  (\PWM5/n6 , \PWM5/n5 , \PWM5/n0 );  // src/OnePWM.v(25)
  AL_MUX \PWM5/u8  (
    .i0(1'b0),
    .i1(pwm_state_read[5]),
    .sel(\PWM5/u8_sel_is_0_o ),
    .o(\PWM5/n8 ));
  and \PWM5/u8_sel_is_0  (\PWM5/u8_sel_is_0_o , \PWM5/n4_neg , \PWM5/n6_neg );
  AL_MUX \PWM5/u9  (
    .i0(\PWM5/n8 ),
    .i1(1'b1),
    .sel(pwm_start_stop[21]),
    .o(\PWM5/n9 ));  // src/OnePWM.v(26)
  reg_ar_as_w1 \PWM6/State_reg  (
    .clk(clk100m),
    .d(\PWM6/n10 ),
    .en(1'b1),
    .reset(~rstn),
    .set(1'b0),
    .q(pwm_state_read[6]));  // src/OnePWM.v(26)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[0]  (
    .i(\PWM6/RemaTxNum[0]_keep ),
    .o(pnumcnt6[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[10]  (
    .i(\PWM6/RemaTxNum[10]_keep ),
    .o(pnumcnt6[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[11]  (
    .i(\PWM6/RemaTxNum[11]_keep ),
    .o(pnumcnt6[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[12]  (
    .i(\PWM6/RemaTxNum[12]_keep ),
    .o(pnumcnt6[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[13]  (
    .i(\PWM6/RemaTxNum[13]_keep ),
    .o(pnumcnt6[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[14]  (
    .i(\PWM6/RemaTxNum[14]_keep ),
    .o(pnumcnt6[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[15]  (
    .i(\PWM6/RemaTxNum[15]_keep ),
    .o(pnumcnt6[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[16]  (
    .i(\PWM6/RemaTxNum[16]_keep ),
    .o(pnumcnt6[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[17]  (
    .i(\PWM6/RemaTxNum[17]_keep ),
    .o(pnumcnt6[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[18]  (
    .i(\PWM6/RemaTxNum[18]_keep ),
    .o(pnumcnt6[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[19]  (
    .i(\PWM6/RemaTxNum[19]_keep ),
    .o(pnumcnt6[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[1]  (
    .i(\PWM6/RemaTxNum[1]_keep ),
    .o(pnumcnt6[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[20]  (
    .i(\PWM6/RemaTxNum[20]_keep ),
    .o(pnumcnt6[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[21]  (
    .i(\PWM6/RemaTxNum[21]_keep ),
    .o(pnumcnt6[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[22]  (
    .i(\PWM6/RemaTxNum[22]_keep ),
    .o(pnumcnt6[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[23]  (
    .i(\PWM6/RemaTxNum[23]_keep ),
    .o(pnumcnt6[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[2]  (
    .i(\PWM6/RemaTxNum[2]_keep ),
    .o(pnumcnt6[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[3]  (
    .i(\PWM6/RemaTxNum[3]_keep ),
    .o(pnumcnt6[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[4]  (
    .i(\PWM6/RemaTxNum[4]_keep ),
    .o(pnumcnt6[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[5]  (
    .i(\PWM6/RemaTxNum[5]_keep ),
    .o(pnumcnt6[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[6]  (
    .i(\PWM6/RemaTxNum[6]_keep ),
    .o(pnumcnt6[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[7]  (
    .i(\PWM6/RemaTxNum[7]_keep ),
    .o(pnumcnt6[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[8]  (
    .i(\PWM6/RemaTxNum[8]_keep ),
    .o(pnumcnt6[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_RemaTxNum[9]  (
    .i(\PWM6/RemaTxNum[9]_keep ),
    .o(pnumcnt6[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_dir  (
    .i(\PWM6/dir_keep ),
    .o(dir[6]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[0]  (
    .i(\PWM6/pnumr[0]_keep ),
    .o(\PWM6/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[10]  (
    .i(\PWM6/pnumr[10]_keep ),
    .o(\PWM6/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[11]  (
    .i(\PWM6/pnumr[11]_keep ),
    .o(\PWM6/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[12]  (
    .i(\PWM6/pnumr[12]_keep ),
    .o(\PWM6/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[13]  (
    .i(\PWM6/pnumr[13]_keep ),
    .o(\PWM6/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[14]  (
    .i(\PWM6/pnumr[14]_keep ),
    .o(\PWM6/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[15]  (
    .i(\PWM6/pnumr[15]_keep ),
    .o(\PWM6/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[16]  (
    .i(\PWM6/pnumr[16]_keep ),
    .o(\PWM6/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[17]  (
    .i(\PWM6/pnumr[17]_keep ),
    .o(\PWM6/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[18]  (
    .i(\PWM6/pnumr[18]_keep ),
    .o(\PWM6/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[19]  (
    .i(\PWM6/pnumr[19]_keep ),
    .o(\PWM6/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[1]  (
    .i(\PWM6/pnumr[1]_keep ),
    .o(\PWM6/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[20]  (
    .i(\PWM6/pnumr[20]_keep ),
    .o(\PWM6/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[21]  (
    .i(\PWM6/pnumr[21]_keep ),
    .o(\PWM6/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[22]  (
    .i(\PWM6/pnumr[22]_keep ),
    .o(\PWM6/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[23]  (
    .i(\PWM6/pnumr[23]_keep ),
    .o(\PWM6/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[24]  (
    .i(\PWM6/pnumr[24]_keep ),
    .o(\PWM6/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[25]  (
    .i(\PWM6/pnumr[25]_keep ),
    .o(\PWM6/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[26]  (
    .i(\PWM6/pnumr[26]_keep ),
    .o(\PWM6/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[27]  (
    .i(\PWM6/pnumr[27]_keep ),
    .o(\PWM6/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[28]  (
    .i(\PWM6/pnumr[28]_keep ),
    .o(\PWM6/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[29]  (
    .i(\PWM6/pnumr[29]_keep ),
    .o(\PWM6/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[2]  (
    .i(\PWM6/pnumr[2]_keep ),
    .o(\PWM6/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[30]  (
    .i(\PWM6/pnumr[30]_keep ),
    .o(\PWM6/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[31]  (
    .i(\PWM6/pnumr[31]_keep ),
    .o(\PWM6/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[3]  (
    .i(\PWM6/pnumr[3]_keep ),
    .o(\PWM6/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[4]  (
    .i(\PWM6/pnumr[4]_keep ),
    .o(\PWM6/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[5]  (
    .i(\PWM6/pnumr[5]_keep ),
    .o(\PWM6/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[6]  (
    .i(\PWM6/pnumr[6]_keep ),
    .o(\PWM6/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[7]  (
    .i(\PWM6/pnumr[7]_keep ),
    .o(\PWM6/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[8]  (
    .i(\PWM6/pnumr[8]_keep ),
    .o(\PWM6/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pnumr[9]  (
    .i(\PWM6/pnumr[9]_keep ),
    .o(\PWM6/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_pwm  (
    .i(\PWM6/pwm_keep ),
    .o(pwm[6]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM6/_bufkeep_stopreq  (
    .i(\PWM6/stopreq_keep ),
    .o(\PWM6/stopreq ));  // src/OnePWM.v(14)
  reg_ar_as_w1 \PWM6/dir_reg  (
    .clk(clk100m),
    .d(\PWM6/n32 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/dir_keep ));  // src/OnePWM.v(58)
  eq_w27 \PWM6/eq0  (
    .i0(\PWM6/FreCnt ),
    .i1(27'b000000000000000000000000000),
    .o(\PWM6/n0 ));  // src/OnePWM.v(15)
  eq_w24 \PWM6/eq1  (
    .i0(pnumcnt6),
    .i1(24'b000000000000000000000001),
    .o(\PWM6/n5 ));  // src/OnePWM.v(25)
  eq_w27 \PWM6/eq2  (
    .i0(\PWM6/FreCnt ),
    .i1({1'b0,\PWM6/FreCntr [26:1]}),
    .o(\PWM6/n17 ));  // src/OnePWM.v(41)
  eq_w27 \PWM6/eq3  (
    .i0(\PWM6/FreCnt ),
    .i1(\PWM6/FreCntr ),
    .o(\PWM6/n18 ));  // src/OnePWM.v(43)
  binary_mux_s1_w1 \PWM6/mux0_b0  (
    .i0(\PWM6/n12 [0]),
    .i1(freq6[0]),
    .sel(\PWM6/n0 ),
    .o(\PWM6/n13 [0]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM6/mux0_b1  (
    .i0(\PWM6/n12 [1]),
    .i1(freq6[1]),
    .sel(\PWM6/n0 ),
    .o(\PWM6/n13 [1]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM6/mux0_b10  (
    .i0(\PWM6/n12 [10]),
    .i1(freq6[10]),
    .sel(\PWM6/n0 ),
    .o(\PWM6/n13 [10]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM6/mux0_b11  (
    .i0(\PWM6/n12 [11]),
    .i1(freq6[11]),
    .sel(\PWM6/n0 ),
    .o(\PWM6/n13 [11]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM6/mux0_b12  (
    .i0(\PWM6/n12 [12]),
    .i1(freq6[12]),
    .sel(\PWM6/n0 ),
    .o(\PWM6/n13 [12]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM6/mux0_b13  (
    .i0(\PWM6/n12 [13]),
    .i1(freq6[13]),
    .sel(\PWM6/n0 ),
    .o(\PWM6/n13 [13]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM6/mux0_b14  (
    .i0(\PWM6/n12 [14]),
    .i1(freq6[14]),
    .sel(\PWM6/n0 ),
    .o(\PWM6/n13 [14]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM6/mux0_b15  (
    .i0(\PWM6/n12 [15]),
    .i1(freq6[15]),
    .sel(\PWM6/n0 ),
    .o(\PWM6/n13 [15]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM6/mux0_b16  (
    .i0(\PWM6/n12 [16]),
    .i1(freq6[16]),
    .sel(\PWM6/n0 ),
    .o(\PWM6/n13 [16]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM6/mux0_b17  (
    .i0(\PWM6/n12 [17]),
    .i1(freq6[17]),
    .sel(\PWM6/n0 ),
    .o(\PWM6/n13 [17]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM6/mux0_b18  (
    .i0(\PWM6/n12 [18]),
    .i1(freq6[18]),
    .sel(\PWM6/n0 ),
    .o(\PWM6/n13 [18]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM6/mux0_b19  (
    .i0(\PWM6/n12 [19]),
    .i1(freq6[19]),
    .sel(\PWM6/n0 ),
    .o(\PWM6/n13 [19]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM6/mux0_b2  (
    .i0(\PWM6/n12 [2]),
    .i1(freq6[2]),
    .sel(\PWM6/n0 ),
    .o(\PWM6/n13 [2]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM6/mux0_b20  (
    .i0(\PWM6/n12 [20]),
    .i1(freq6[20]),
    .sel(\PWM6/n0 ),
    .o(\PWM6/n13 [20]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM6/mux0_b21  (
    .i0(\PWM6/n12 [21]),
    .i1(freq6[21]),
    .sel(\PWM6/n0 ),
    .o(\PWM6/n13 [21]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM6/mux0_b22  (
    .i0(\PWM6/n12 [22]),
    .i1(freq6[22]),
    .sel(\PWM6/n0 ),
    .o(\PWM6/n13 [22]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM6/mux0_b23  (
    .i0(\PWM6/n12 [23]),
    .i1(freq6[23]),
    .sel(\PWM6/n0 ),
    .o(\PWM6/n13 [23]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM6/mux0_b24  (
    .i0(\PWM6/n12 [24]),
    .i1(freq6[24]),
    .sel(\PWM6/n0 ),
    .o(\PWM6/n13 [24]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM6/mux0_b25  (
    .i0(\PWM6/n12 [25]),
    .i1(freq6[25]),
    .sel(\PWM6/n0 ),
    .o(\PWM6/n13 [25]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM6/mux0_b26  (
    .i0(\PWM6/n12 [26]),
    .i1(freq6[26]),
    .sel(\PWM6/n0 ),
    .o(\PWM6/n13 [26]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM6/mux0_b3  (
    .i0(\PWM6/n12 [3]),
    .i1(freq6[3]),
    .sel(\PWM6/n0 ),
    .o(\PWM6/n13 [3]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM6/mux0_b4  (
    .i0(\PWM6/n12 [4]),
    .i1(freq6[4]),
    .sel(\PWM6/n0 ),
    .o(\PWM6/n13 [4]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM6/mux0_b5  (
    .i0(\PWM6/n12 [5]),
    .i1(freq6[5]),
    .sel(\PWM6/n0 ),
    .o(\PWM6/n13 [5]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM6/mux0_b6  (
    .i0(\PWM6/n12 [6]),
    .i1(freq6[6]),
    .sel(\PWM6/n0 ),
    .o(\PWM6/n13 [6]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM6/mux0_b7  (
    .i0(\PWM6/n12 [7]),
    .i1(freq6[7]),
    .sel(\PWM6/n0 ),
    .o(\PWM6/n13 [7]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM6/mux0_b8  (
    .i0(\PWM6/n12 [8]),
    .i1(freq6[8]),
    .sel(\PWM6/n0 ),
    .o(\PWM6/n13 [8]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM6/mux0_b9  (
    .i0(\PWM6/n12 [9]),
    .i1(freq6[9]),
    .sel(\PWM6/n0 ),
    .o(\PWM6/n13 [9]));  // src/OnePWM.v(32)
  and \PWM6/mux3_b0_sel_is_3  (\PWM6/mux3_b0_sel_is_3_o , \PWM6/n11 , \PWM6/n0 );
  binary_mux_s1_w1 \PWM6/mux4_b0  (
    .i0(\PWM6/pnumr [0]),
    .i1(1'b0),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n22 [0]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux4_b1  (
    .i0(\PWM6/pnumr [1]),
    .i1(1'b0),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n22 [1]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux4_b10  (
    .i0(\PWM6/pnumr [10]),
    .i1(1'b0),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n22 [10]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux4_b11  (
    .i0(\PWM6/pnumr [11]),
    .i1(1'b0),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n22 [11]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux4_b12  (
    .i0(\PWM6/pnumr [12]),
    .i1(1'b0),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n22 [12]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux4_b13  (
    .i0(\PWM6/pnumr [13]),
    .i1(1'b0),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n22 [13]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux4_b14  (
    .i0(\PWM6/pnumr [14]),
    .i1(1'b0),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n22 [14]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux4_b15  (
    .i0(\PWM6/pnumr [15]),
    .i1(1'b0),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n22 [15]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux4_b16  (
    .i0(\PWM6/pnumr [16]),
    .i1(1'b0),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n22 [16]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux4_b17  (
    .i0(\PWM6/pnumr [17]),
    .i1(1'b0),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n22 [17]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux4_b18  (
    .i0(\PWM6/pnumr [18]),
    .i1(1'b0),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n22 [18]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux4_b19  (
    .i0(\PWM6/pnumr [19]),
    .i1(1'b0),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n22 [19]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux4_b2  (
    .i0(\PWM6/pnumr [2]),
    .i1(1'b0),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n22 [2]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux4_b20  (
    .i0(\PWM6/pnumr [20]),
    .i1(1'b0),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n22 [20]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux4_b21  (
    .i0(\PWM6/pnumr [21]),
    .i1(1'b0),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n22 [21]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux4_b22  (
    .i0(\PWM6/pnumr [22]),
    .i1(1'b0),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n22 [22]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux4_b23  (
    .i0(\PWM6/pnumr [23]),
    .i1(1'b0),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n22 [23]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux4_b24  (
    .i0(\PWM6/pnumr [24]),
    .i1(1'b0),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n22 [24]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux4_b25  (
    .i0(\PWM6/pnumr [25]),
    .i1(1'b0),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n22 [25]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux4_b26  (
    .i0(\PWM6/pnumr [26]),
    .i1(1'b0),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n22 [26]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux4_b27  (
    .i0(\PWM6/pnumr [27]),
    .i1(1'b0),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n22 [27]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux4_b28  (
    .i0(\PWM6/pnumr [28]),
    .i1(1'b0),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n22 [28]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux4_b29  (
    .i0(\PWM6/pnumr [29]),
    .i1(1'b0),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n22 [29]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux4_b3  (
    .i0(\PWM6/pnumr [3]),
    .i1(1'b0),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n22 [3]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux4_b30  (
    .i0(\PWM6/pnumr [30]),
    .i1(1'b0),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n22 [30]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux4_b31  (
    .i0(\PWM6/pnumr [31]),
    .i1(1'b0),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n22 [31]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux4_b4  (
    .i0(\PWM6/pnumr [4]),
    .i1(1'b0),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n22 [4]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux4_b5  (
    .i0(\PWM6/pnumr [5]),
    .i1(1'b0),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n22 [5]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux4_b6  (
    .i0(\PWM6/pnumr [6]),
    .i1(1'b0),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n22 [6]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux4_b7  (
    .i0(\PWM6/pnumr [7]),
    .i1(1'b0),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n22 [7]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux4_b8  (
    .i0(\PWM6/pnumr [8]),
    .i1(1'b0),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n22 [8]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux4_b9  (
    .i0(\PWM6/pnumr [9]),
    .i1(1'b0),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n22 [9]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux5_b0  (
    .i0(\PWM6/n22 [0]),
    .i1(pnum6[0]),
    .sel(pnum6[32]),
    .o(\PWM6/n23 [0]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux5_b1  (
    .i0(\PWM6/n22 [1]),
    .i1(pnum6[1]),
    .sel(pnum6[32]),
    .o(\PWM6/n23 [1]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux5_b10  (
    .i0(\PWM6/n22 [10]),
    .i1(pnum6[10]),
    .sel(pnum6[32]),
    .o(\PWM6/n23 [10]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux5_b11  (
    .i0(\PWM6/n22 [11]),
    .i1(pnum6[11]),
    .sel(pnum6[32]),
    .o(\PWM6/n23 [11]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux5_b12  (
    .i0(\PWM6/n22 [12]),
    .i1(pnum6[12]),
    .sel(pnum6[32]),
    .o(\PWM6/n23 [12]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux5_b13  (
    .i0(\PWM6/n22 [13]),
    .i1(pnum6[13]),
    .sel(pnum6[32]),
    .o(\PWM6/n23 [13]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux5_b14  (
    .i0(\PWM6/n22 [14]),
    .i1(pnum6[14]),
    .sel(pnum6[32]),
    .o(\PWM6/n23 [14]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux5_b15  (
    .i0(\PWM6/n22 [15]),
    .i1(pnum6[15]),
    .sel(pnum6[32]),
    .o(\PWM6/n23 [15]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux5_b16  (
    .i0(\PWM6/n22 [16]),
    .i1(pnum6[16]),
    .sel(pnum6[32]),
    .o(\PWM6/n23 [16]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux5_b17  (
    .i0(\PWM6/n22 [17]),
    .i1(pnum6[17]),
    .sel(pnum6[32]),
    .o(\PWM6/n23 [17]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux5_b18  (
    .i0(\PWM6/n22 [18]),
    .i1(pnum6[18]),
    .sel(pnum6[32]),
    .o(\PWM6/n23 [18]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux5_b19  (
    .i0(\PWM6/n22 [19]),
    .i1(pnum6[19]),
    .sel(pnum6[32]),
    .o(\PWM6/n23 [19]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux5_b2  (
    .i0(\PWM6/n22 [2]),
    .i1(pnum6[2]),
    .sel(pnum6[32]),
    .o(\PWM6/n23 [2]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux5_b20  (
    .i0(\PWM6/n22 [20]),
    .i1(pnum6[20]),
    .sel(pnum6[32]),
    .o(\PWM6/n23 [20]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux5_b21  (
    .i0(\PWM6/n22 [21]),
    .i1(pnum6[21]),
    .sel(pnum6[32]),
    .o(\PWM6/n23 [21]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux5_b22  (
    .i0(\PWM6/n22 [22]),
    .i1(pnum6[22]),
    .sel(pnum6[32]),
    .o(\PWM6/n23 [22]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux5_b23  (
    .i0(\PWM6/n22 [23]),
    .i1(pnum6[23]),
    .sel(pnum6[32]),
    .o(\PWM6/n23 [23]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux5_b24  (
    .i0(\PWM6/n22 [24]),
    .i1(pnum6[24]),
    .sel(pnum6[32]),
    .o(\PWM6/n23 [24]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux5_b25  (
    .i0(\PWM6/n22 [25]),
    .i1(pnum6[25]),
    .sel(pnum6[32]),
    .o(\PWM6/n23 [25]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux5_b26  (
    .i0(\PWM6/n22 [26]),
    .i1(pnum6[26]),
    .sel(pnum6[32]),
    .o(\PWM6/n23 [26]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux5_b27  (
    .i0(\PWM6/n22 [27]),
    .i1(pnum6[27]),
    .sel(pnum6[32]),
    .o(\PWM6/n23 [27]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux5_b28  (
    .i0(\PWM6/n22 [28]),
    .i1(pnum6[28]),
    .sel(pnum6[32]),
    .o(\PWM6/n23 [28]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux5_b29  (
    .i0(\PWM6/n22 [29]),
    .i1(pnum6[29]),
    .sel(pnum6[32]),
    .o(\PWM6/n23 [29]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux5_b3  (
    .i0(\PWM6/n22 [3]),
    .i1(pnum6[3]),
    .sel(pnum6[32]),
    .o(\PWM6/n23 [3]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux5_b30  (
    .i0(\PWM6/n22 [30]),
    .i1(pnum6[30]),
    .sel(pnum6[32]),
    .o(\PWM6/n23 [30]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux5_b31  (
    .i0(\PWM6/n22 [31]),
    .i1(pnum6[31]),
    .sel(pnum6[32]),
    .o(\PWM6/n23 [31]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux5_b4  (
    .i0(\PWM6/n22 [4]),
    .i1(pnum6[4]),
    .sel(pnum6[32]),
    .o(\PWM6/n23 [4]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux5_b5  (
    .i0(\PWM6/n22 [5]),
    .i1(pnum6[5]),
    .sel(pnum6[32]),
    .o(\PWM6/n23 [5]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux5_b6  (
    .i0(\PWM6/n22 [6]),
    .i1(pnum6[6]),
    .sel(pnum6[32]),
    .o(\PWM6/n23 [6]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux5_b7  (
    .i0(\PWM6/n22 [7]),
    .i1(pnum6[7]),
    .sel(pnum6[32]),
    .o(\PWM6/n23 [7]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux5_b8  (
    .i0(\PWM6/n22 [8]),
    .i1(pnum6[8]),
    .sel(pnum6[32]),
    .o(\PWM6/n23 [8]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux5_b9  (
    .i0(\PWM6/n22 [9]),
    .i1(pnum6[9]),
    .sel(pnum6[32]),
    .o(\PWM6/n23 [9]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM6/mux6_b0  (
    .i0(\PWM6/pnumr [0]),
    .i1(\PWM6/n26 [0]),
    .sel(\PWM6/n25 ),
    .o(\PWM6/n27 [0]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM6/mux6_b1  (
    .i0(\PWM6/pnumr [1]),
    .i1(\PWM6/n26 [1]),
    .sel(\PWM6/n25 ),
    .o(\PWM6/n27 [1]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM6/mux6_b10  (
    .i0(\PWM6/pnumr [10]),
    .i1(\PWM6/n26 [10]),
    .sel(\PWM6/n25 ),
    .o(\PWM6/n27 [10]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM6/mux6_b11  (
    .i0(\PWM6/pnumr [11]),
    .i1(\PWM6/n26 [11]),
    .sel(\PWM6/n25 ),
    .o(\PWM6/n27 [11]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM6/mux6_b12  (
    .i0(\PWM6/pnumr [12]),
    .i1(\PWM6/n26 [12]),
    .sel(\PWM6/n25 ),
    .o(\PWM6/n27 [12]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM6/mux6_b13  (
    .i0(\PWM6/pnumr [13]),
    .i1(\PWM6/n26 [13]),
    .sel(\PWM6/n25 ),
    .o(\PWM6/n27 [13]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM6/mux6_b14  (
    .i0(\PWM6/pnumr [14]),
    .i1(\PWM6/n26 [14]),
    .sel(\PWM6/n25 ),
    .o(\PWM6/n27 [14]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM6/mux6_b15  (
    .i0(\PWM6/pnumr [15]),
    .i1(\PWM6/n26 [15]),
    .sel(\PWM6/n25 ),
    .o(\PWM6/n27 [15]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM6/mux6_b16  (
    .i0(\PWM6/pnumr [16]),
    .i1(\PWM6/n26 [16]),
    .sel(\PWM6/n25 ),
    .o(\PWM6/n27 [16]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM6/mux6_b17  (
    .i0(\PWM6/pnumr [17]),
    .i1(\PWM6/n26 [17]),
    .sel(\PWM6/n25 ),
    .o(\PWM6/n27 [17]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM6/mux6_b18  (
    .i0(\PWM6/pnumr [18]),
    .i1(\PWM6/n26 [18]),
    .sel(\PWM6/n25 ),
    .o(\PWM6/n27 [18]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM6/mux6_b19  (
    .i0(\PWM6/pnumr [19]),
    .i1(\PWM6/n26 [19]),
    .sel(\PWM6/n25 ),
    .o(\PWM6/n27 [19]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM6/mux6_b2  (
    .i0(\PWM6/pnumr [2]),
    .i1(\PWM6/n26 [2]),
    .sel(\PWM6/n25 ),
    .o(\PWM6/n27 [2]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM6/mux6_b20  (
    .i0(\PWM6/pnumr [20]),
    .i1(\PWM6/n26 [20]),
    .sel(\PWM6/n25 ),
    .o(\PWM6/n27 [20]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM6/mux6_b21  (
    .i0(\PWM6/pnumr [21]),
    .i1(\PWM6/n26 [21]),
    .sel(\PWM6/n25 ),
    .o(\PWM6/n27 [21]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM6/mux6_b22  (
    .i0(\PWM6/pnumr [22]),
    .i1(\PWM6/n26 [22]),
    .sel(\PWM6/n25 ),
    .o(\PWM6/n27 [22]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM6/mux6_b23  (
    .i0(\PWM6/pnumr [23]),
    .i1(\PWM6/n26 [23]),
    .sel(\PWM6/n25 ),
    .o(\PWM6/n27 [23]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM6/mux6_b3  (
    .i0(\PWM6/pnumr [3]),
    .i1(\PWM6/n26 [3]),
    .sel(\PWM6/n25 ),
    .o(\PWM6/n27 [3]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM6/mux6_b4  (
    .i0(\PWM6/pnumr [4]),
    .i1(\PWM6/n26 [4]),
    .sel(\PWM6/n25 ),
    .o(\PWM6/n27 [4]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM6/mux6_b5  (
    .i0(\PWM6/pnumr [5]),
    .i1(\PWM6/n26 [5]),
    .sel(\PWM6/n25 ),
    .o(\PWM6/n27 [5]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM6/mux6_b6  (
    .i0(\PWM6/pnumr [6]),
    .i1(\PWM6/n26 [6]),
    .sel(\PWM6/n25 ),
    .o(\PWM6/n27 [6]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM6/mux6_b7  (
    .i0(\PWM6/pnumr [7]),
    .i1(\PWM6/n26 [7]),
    .sel(\PWM6/n25 ),
    .o(\PWM6/n27 [7]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM6/mux6_b8  (
    .i0(\PWM6/pnumr [8]),
    .i1(\PWM6/n26 [8]),
    .sel(\PWM6/n25 ),
    .o(\PWM6/n27 [8]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM6/mux6_b9  (
    .i0(\PWM6/pnumr [9]),
    .i1(\PWM6/n26 [9]),
    .sel(\PWM6/n25 ),
    .o(\PWM6/n27 [9]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM6/mux7_b0  (
    .i0(pnumcnt6[0]),
    .i1(\PWM6/n27 [0]),
    .sel(\PWM6/n24 ),
    .o(\PWM6/n29 [0]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux7_b1  (
    .i0(pnumcnt6[1]),
    .i1(\PWM6/n27 [1]),
    .sel(\PWM6/n24 ),
    .o(\PWM6/n29 [1]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux7_b10  (
    .i0(pnumcnt6[10]),
    .i1(\PWM6/n27 [10]),
    .sel(\PWM6/n24 ),
    .o(\PWM6/n29 [10]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux7_b11  (
    .i0(pnumcnt6[11]),
    .i1(\PWM6/n27 [11]),
    .sel(\PWM6/n24 ),
    .o(\PWM6/n29 [11]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux7_b12  (
    .i0(pnumcnt6[12]),
    .i1(\PWM6/n27 [12]),
    .sel(\PWM6/n24 ),
    .o(\PWM6/n29 [12]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux7_b13  (
    .i0(pnumcnt6[13]),
    .i1(\PWM6/n27 [13]),
    .sel(\PWM6/n24 ),
    .o(\PWM6/n29 [13]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux7_b14  (
    .i0(pnumcnt6[14]),
    .i1(\PWM6/n27 [14]),
    .sel(\PWM6/n24 ),
    .o(\PWM6/n29 [14]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux7_b15  (
    .i0(pnumcnt6[15]),
    .i1(\PWM6/n27 [15]),
    .sel(\PWM6/n24 ),
    .o(\PWM6/n29 [15]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux7_b16  (
    .i0(pnumcnt6[16]),
    .i1(\PWM6/n27 [16]),
    .sel(\PWM6/n24 ),
    .o(\PWM6/n29 [16]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux7_b17  (
    .i0(pnumcnt6[17]),
    .i1(\PWM6/n27 [17]),
    .sel(\PWM6/n24 ),
    .o(\PWM6/n29 [17]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux7_b18  (
    .i0(pnumcnt6[18]),
    .i1(\PWM6/n27 [18]),
    .sel(\PWM6/n24 ),
    .o(\PWM6/n29 [18]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux7_b19  (
    .i0(pnumcnt6[19]),
    .i1(\PWM6/n27 [19]),
    .sel(\PWM6/n24 ),
    .o(\PWM6/n29 [19]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux7_b2  (
    .i0(pnumcnt6[2]),
    .i1(\PWM6/n27 [2]),
    .sel(\PWM6/n24 ),
    .o(\PWM6/n29 [2]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux7_b20  (
    .i0(pnumcnt6[20]),
    .i1(\PWM6/n27 [20]),
    .sel(\PWM6/n24 ),
    .o(\PWM6/n29 [20]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux7_b21  (
    .i0(pnumcnt6[21]),
    .i1(\PWM6/n27 [21]),
    .sel(\PWM6/n24 ),
    .o(\PWM6/n29 [21]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux7_b22  (
    .i0(pnumcnt6[22]),
    .i1(\PWM6/n27 [22]),
    .sel(\PWM6/n24 ),
    .o(\PWM6/n29 [22]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux7_b23  (
    .i0(pnumcnt6[23]),
    .i1(\PWM6/n27 [23]),
    .sel(\PWM6/n24 ),
    .o(\PWM6/n29 [23]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux7_b3  (
    .i0(pnumcnt6[3]),
    .i1(\PWM6/n27 [3]),
    .sel(\PWM6/n24 ),
    .o(\PWM6/n29 [3]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux7_b4  (
    .i0(pnumcnt6[4]),
    .i1(\PWM6/n27 [4]),
    .sel(\PWM6/n24 ),
    .o(\PWM6/n29 [4]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux7_b5  (
    .i0(pnumcnt6[5]),
    .i1(\PWM6/n27 [5]),
    .sel(\PWM6/n24 ),
    .o(\PWM6/n29 [5]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux7_b6  (
    .i0(pnumcnt6[6]),
    .i1(\PWM6/n27 [6]),
    .sel(\PWM6/n24 ),
    .o(\PWM6/n29 [6]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux7_b7  (
    .i0(pnumcnt6[7]),
    .i1(\PWM6/n27 [7]),
    .sel(\PWM6/n24 ),
    .o(\PWM6/n29 [7]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux7_b8  (
    .i0(pnumcnt6[8]),
    .i1(\PWM6/n27 [8]),
    .sel(\PWM6/n24 ),
    .o(\PWM6/n29 [8]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux7_b9  (
    .i0(pnumcnt6[9]),
    .i1(\PWM6/n27 [9]),
    .sel(\PWM6/n24 ),
    .o(\PWM6/n29 [9]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux8_b0  (
    .i0(\PWM6/n29 [0]),
    .i1(\PWM6/pnumr [0]),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n31 [0]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux8_b1  (
    .i0(\PWM6/n29 [1]),
    .i1(\PWM6/pnumr [1]),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n31 [1]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux8_b10  (
    .i0(\PWM6/n29 [10]),
    .i1(\PWM6/pnumr [10]),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n31 [10]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux8_b11  (
    .i0(\PWM6/n29 [11]),
    .i1(\PWM6/pnumr [11]),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n31 [11]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux8_b12  (
    .i0(\PWM6/n29 [12]),
    .i1(\PWM6/pnumr [12]),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n31 [12]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux8_b13  (
    .i0(\PWM6/n29 [13]),
    .i1(\PWM6/pnumr [13]),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n31 [13]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux8_b14  (
    .i0(\PWM6/n29 [14]),
    .i1(\PWM6/pnumr [14]),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n31 [14]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux8_b15  (
    .i0(\PWM6/n29 [15]),
    .i1(\PWM6/pnumr [15]),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n31 [15]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux8_b16  (
    .i0(\PWM6/n29 [16]),
    .i1(\PWM6/pnumr [16]),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n31 [16]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux8_b17  (
    .i0(\PWM6/n29 [17]),
    .i1(\PWM6/pnumr [17]),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n31 [17]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux8_b18  (
    .i0(\PWM6/n29 [18]),
    .i1(\PWM6/pnumr [18]),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n31 [18]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux8_b19  (
    .i0(\PWM6/n29 [19]),
    .i1(\PWM6/pnumr [19]),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n31 [19]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux8_b2  (
    .i0(\PWM6/n29 [2]),
    .i1(\PWM6/pnumr [2]),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n31 [2]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux8_b20  (
    .i0(\PWM6/n29 [20]),
    .i1(\PWM6/pnumr [20]),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n31 [20]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux8_b21  (
    .i0(\PWM6/n29 [21]),
    .i1(\PWM6/pnumr [21]),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n31 [21]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux8_b22  (
    .i0(\PWM6/n29 [22]),
    .i1(\PWM6/pnumr [22]),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n31 [22]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux8_b23  (
    .i0(\PWM6/n29 [23]),
    .i1(\PWM6/pnumr [23]),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n31 [23]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux8_b3  (
    .i0(\PWM6/n29 [3]),
    .i1(\PWM6/pnumr [3]),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n31 [3]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux8_b4  (
    .i0(\PWM6/n29 [4]),
    .i1(\PWM6/pnumr [4]),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n31 [4]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux8_b5  (
    .i0(\PWM6/n29 [5]),
    .i1(\PWM6/pnumr [5]),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n31 [5]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux8_b6  (
    .i0(\PWM6/n29 [6]),
    .i1(\PWM6/pnumr [6]),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n31 [6]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux8_b7  (
    .i0(\PWM6/n29 [7]),
    .i1(\PWM6/pnumr [7]),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n31 [7]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux8_b8  (
    .i0(\PWM6/n29 [8]),
    .i1(\PWM6/pnumr [8]),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n31 [8]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM6/mux8_b9  (
    .i0(\PWM6/n29 [9]),
    .i1(\PWM6/pnumr [9]),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n31 [9]));  // src/OnePWM.v(57)
  not \PWM6/n17_inv  (\PWM6/n17_neg , \PWM6/n17 );
  not \PWM6/n25_inv  (\PWM6/n25_neg , \PWM6/n25 );
  not \PWM6/n4_inv  (\PWM6/n4_neg , \PWM6/n4 );
  not \PWM6/n6_inv  (\PWM6/n6_neg , \PWM6/n6 );
  ne_w24 \PWM6/neq0  (
    .i0(pnumcnt6),
    .i1(24'b000000000000000000000000),
    .o(\PWM6/n25 ));  // src/OnePWM.v(55)
  reg_sr_ss_w1 \PWM6/pwm_reg  (
    .clk(clk100m),
    .d(pwm[6]),
    .en(1'b1),
    .reset(~\PWM6/u14_sel_is_1_o ),
    .set(\PWM6/n18 ),
    .q(\PWM6/pwm_keep ));  // src/OnePWM.v(45)
  reg_sr_as_w1 \PWM6/reg0_b0  (
    .clk(clk100m),
    .d(\PWM6/n13 [0]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [0]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b1  (
    .clk(clk100m),
    .d(\PWM6/n13 [1]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [1]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b10  (
    .clk(clk100m),
    .d(\PWM6/n13 [10]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [10]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b11  (
    .clk(clk100m),
    .d(\PWM6/n13 [11]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [11]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b12  (
    .clk(clk100m),
    .d(\PWM6/n13 [12]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [12]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b13  (
    .clk(clk100m),
    .d(\PWM6/n13 [13]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [13]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b14  (
    .clk(clk100m),
    .d(\PWM6/n13 [14]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [14]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b15  (
    .clk(clk100m),
    .d(\PWM6/n13 [15]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [15]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b16  (
    .clk(clk100m),
    .d(\PWM6/n13 [16]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [16]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b17  (
    .clk(clk100m),
    .d(\PWM6/n13 [17]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [17]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b18  (
    .clk(clk100m),
    .d(\PWM6/n13 [18]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [18]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b19  (
    .clk(clk100m),
    .d(\PWM6/n13 [19]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [19]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b2  (
    .clk(clk100m),
    .d(\PWM6/n13 [2]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [2]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b20  (
    .clk(clk100m),
    .d(\PWM6/n13 [20]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [20]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b21  (
    .clk(clk100m),
    .d(\PWM6/n13 [21]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [21]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b22  (
    .clk(clk100m),
    .d(\PWM6/n13 [22]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [22]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b23  (
    .clk(clk100m),
    .d(\PWM6/n13 [23]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [23]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b24  (
    .clk(clk100m),
    .d(\PWM6/n13 [24]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [24]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b25  (
    .clk(clk100m),
    .d(\PWM6/n13 [25]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [25]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b26  (
    .clk(clk100m),
    .d(\PWM6/n13 [26]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [26]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b3  (
    .clk(clk100m),
    .d(\PWM6/n13 [3]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [3]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b4  (
    .clk(clk100m),
    .d(\PWM6/n13 [4]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [4]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b5  (
    .clk(clk100m),
    .d(\PWM6/n13 [5]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [5]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b6  (
    .clk(clk100m),
    .d(\PWM6/n13 [6]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [6]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b7  (
    .clk(clk100m),
    .d(\PWM6/n13 [7]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [7]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b8  (
    .clk(clk100m),
    .d(\PWM6/n13 [8]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [8]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM6/reg0_b9  (
    .clk(clk100m),
    .d(\PWM6/n13 [9]),
    .en(1'b1),
    .reset(~\PWM6/n11 ),
    .set(1'b0),
    .q(\PWM6/FreCnt [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b0  (
    .clk(clk100m),
    .d(freq6[0]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [0]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b1  (
    .clk(clk100m),
    .d(freq6[1]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [1]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b10  (
    .clk(clk100m),
    .d(freq6[10]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [10]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b11  (
    .clk(clk100m),
    .d(freq6[11]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [11]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b12  (
    .clk(clk100m),
    .d(freq6[12]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [12]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b13  (
    .clk(clk100m),
    .d(freq6[13]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [13]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b14  (
    .clk(clk100m),
    .d(freq6[14]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [14]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b15  (
    .clk(clk100m),
    .d(freq6[15]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [15]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b16  (
    .clk(clk100m),
    .d(freq6[16]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [16]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b17  (
    .clk(clk100m),
    .d(freq6[17]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [17]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b18  (
    .clk(clk100m),
    .d(freq6[18]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [18]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b19  (
    .clk(clk100m),
    .d(freq6[19]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [19]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b2  (
    .clk(clk100m),
    .d(freq6[2]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [2]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b20  (
    .clk(clk100m),
    .d(freq6[20]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [20]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b21  (
    .clk(clk100m),
    .d(freq6[21]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [21]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b22  (
    .clk(clk100m),
    .d(freq6[22]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [22]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b23  (
    .clk(clk100m),
    .d(freq6[23]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [23]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b24  (
    .clk(clk100m),
    .d(freq6[24]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [24]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b25  (
    .clk(clk100m),
    .d(freq6[25]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [25]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b26  (
    .clk(clk100m),
    .d(freq6[26]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [26]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b3  (
    .clk(clk100m),
    .d(freq6[3]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [3]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b4  (
    .clk(clk100m),
    .d(freq6[4]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [4]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b5  (
    .clk(clk100m),
    .d(freq6[5]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [5]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b6  (
    .clk(clk100m),
    .d(freq6[6]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [6]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b7  (
    .clk(clk100m),
    .d(freq6[7]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [7]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b8  (
    .clk(clk100m),
    .d(freq6[8]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [8]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg1_b9  (
    .clk(clk100m),
    .d(freq6[9]),
    .en(\PWM6/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/FreCntr [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM6/reg2_b0  (
    .clk(clk100m),
    .d(\PWM6/n23 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[0]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b1  (
    .clk(clk100m),
    .d(\PWM6/n23 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[1]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b10  (
    .clk(clk100m),
    .d(\PWM6/n23 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[10]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b11  (
    .clk(clk100m),
    .d(\PWM6/n23 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[11]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b12  (
    .clk(clk100m),
    .d(\PWM6/n23 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[12]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b13  (
    .clk(clk100m),
    .d(\PWM6/n23 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[13]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b14  (
    .clk(clk100m),
    .d(\PWM6/n23 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[14]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b15  (
    .clk(clk100m),
    .d(\PWM6/n23 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[15]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b16  (
    .clk(clk100m),
    .d(\PWM6/n23 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[16]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b17  (
    .clk(clk100m),
    .d(\PWM6/n23 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[17]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b18  (
    .clk(clk100m),
    .d(\PWM6/n23 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[18]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b19  (
    .clk(clk100m),
    .d(\PWM6/n23 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[19]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b2  (
    .clk(clk100m),
    .d(\PWM6/n23 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[2]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b20  (
    .clk(clk100m),
    .d(\PWM6/n23 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[20]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b21  (
    .clk(clk100m),
    .d(\PWM6/n23 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[21]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b22  (
    .clk(clk100m),
    .d(\PWM6/n23 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[22]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b23  (
    .clk(clk100m),
    .d(\PWM6/n23 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[23]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b24  (
    .clk(clk100m),
    .d(\PWM6/n23 [24]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[24]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b25  (
    .clk(clk100m),
    .d(\PWM6/n23 [25]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[25]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b26  (
    .clk(clk100m),
    .d(\PWM6/n23 [26]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[26]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b27  (
    .clk(clk100m),
    .d(\PWM6/n23 [27]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[27]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b28  (
    .clk(clk100m),
    .d(\PWM6/n23 [28]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[28]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b29  (
    .clk(clk100m),
    .d(\PWM6/n23 [29]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[29]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b3  (
    .clk(clk100m),
    .d(\PWM6/n23 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[3]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b30  (
    .clk(clk100m),
    .d(\PWM6/n23 [30]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[30]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b31  (
    .clk(clk100m),
    .d(\PWM6/n23 [31]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[31]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b4  (
    .clk(clk100m),
    .d(\PWM6/n23 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[4]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b5  (
    .clk(clk100m),
    .d(\PWM6/n23 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[5]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b6  (
    .clk(clk100m),
    .d(\PWM6/n23 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[6]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b7  (
    .clk(clk100m),
    .d(\PWM6/n23 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[7]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b8  (
    .clk(clk100m),
    .d(\PWM6/n23 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[8]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg2_b9  (
    .clk(clk100m),
    .d(\PWM6/n23 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/pnumr[9]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM6/reg3_b0  (
    .clk(clk100m),
    .d(\PWM6/n31 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[0]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b1  (
    .clk(clk100m),
    .d(\PWM6/n31 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[1]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b10  (
    .clk(clk100m),
    .d(\PWM6/n31 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[10]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b11  (
    .clk(clk100m),
    .d(\PWM6/n31 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[11]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b12  (
    .clk(clk100m),
    .d(\PWM6/n31 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[12]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b13  (
    .clk(clk100m),
    .d(\PWM6/n31 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[13]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b14  (
    .clk(clk100m),
    .d(\PWM6/n31 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[14]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b15  (
    .clk(clk100m),
    .d(\PWM6/n31 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[15]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b16  (
    .clk(clk100m),
    .d(\PWM6/n31 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[16]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b17  (
    .clk(clk100m),
    .d(\PWM6/n31 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[17]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b18  (
    .clk(clk100m),
    .d(\PWM6/n31 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[18]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b19  (
    .clk(clk100m),
    .d(\PWM6/n31 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[19]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b2  (
    .clk(clk100m),
    .d(\PWM6/n31 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[2]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b20  (
    .clk(clk100m),
    .d(\PWM6/n31 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[20]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b21  (
    .clk(clk100m),
    .d(\PWM6/n31 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[21]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b22  (
    .clk(clk100m),
    .d(\PWM6/n31 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[22]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b23  (
    .clk(clk100m),
    .d(\PWM6/n31 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[23]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b3  (
    .clk(clk100m),
    .d(\PWM6/n31 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[3]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b4  (
    .clk(clk100m),
    .d(\PWM6/n31 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[4]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b5  (
    .clk(clk100m),
    .d(\PWM6/n31 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[5]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b6  (
    .clk(clk100m),
    .d(\PWM6/n31 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[6]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b7  (
    .clk(clk100m),
    .d(\PWM6/n31 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[7]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b8  (
    .clk(clk100m),
    .d(\PWM6/n31 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[8]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM6/reg3_b9  (
    .clk(clk100m),
    .d(\PWM6/n31 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM6/RemaTxNum[9]_keep ));  // src/OnePWM.v(58)
  reg_ar_ss_w1 \PWM6/stopreq_reg  (
    .clk(clk100m),
    .d(\PWM6/n1 ),
    .en(1'b1),
    .reset(1'b0),
    .set(pwm_start_stop[6]),
    .q(\PWM6/stopreq_keep ));  // src/OnePWM.v(15)
  add_pu27_mu27_o27 \PWM6/sub0  (
    .i0(\PWM6/FreCnt ),
    .i1(27'b000000000000000000000000001),
    .o(\PWM6/n12 [26:0]));  // src/OnePWM.v(32)
  add_pu24_mu24_o24 \PWM6/sub1  (
    .i0(pnumcnt6),
    .i1(24'b000000000000000000000001),
    .o(\PWM6/n26 [23:0]));  // src/OnePWM.v(55)
  AL_MUX \PWM6/u10  (
    .i0(1'b0),
    .i1(\PWM6/n9 ),
    .sel(n17),
    .o(\PWM6/n10 ));  // src/OnePWM.v(26)
  or \PWM6/u11  (\PWM6/n11 , pwm_state_read[6], pwm_start_stop[22]);  // src/OnePWM.v(30)
  and \PWM6/u14_sel_is_1  (\PWM6/u14_sel_is_1_o , pwm_state_read[6], \PWM6/n17_neg );
  and \PWM6/u15  (\PWM6/n24 , \PWM6/n0 , pwm_state_read[6]);  // src/OnePWM.v(54)
  and \PWM6/u17_sel_is_1  (\PWM6/u17_sel_is_1_o , \PWM6/n24 , \PWM6/n25_neg );
  not \PWM6/u17_sel_is_1_o_inv  (\PWM6/u17_sel_is_1_o_neg , \PWM6/u17_sel_is_1_o );
  AL_MUX \PWM6/u18  (
    .i0(\PWM6/pnumr [31]),
    .i1(dir[6]),
    .sel(\PWM6/u18_sel_is_0_o ),
    .o(\PWM6/n32 ));
  and \PWM6/u18_sel_is_0  (\PWM6/u18_sel_is_0_o , \pwm_start_stop[22]_neg , \PWM6/u17_sel_is_1_o_neg );
  AL_MUX \PWM6/u2  (
    .i0(\PWM6/stopreq ),
    .i1(1'b0),
    .sel(\PWM6/n0 ),
    .o(\PWM6/n1 ));  // src/OnePWM.v(15)
  and \PWM6/u5  (\PWM6/n4 , \PWM6/stopreq , \PWM6/n0 );  // src/OnePWM.v(23)
  and \PWM6/u6  (\PWM6/n6 , \PWM6/n5 , \PWM6/n0 );  // src/OnePWM.v(25)
  AL_MUX \PWM6/u8  (
    .i0(1'b0),
    .i1(pwm_state_read[6]),
    .sel(\PWM6/u8_sel_is_0_o ),
    .o(\PWM6/n8 ));
  and \PWM6/u8_sel_is_0  (\PWM6/u8_sel_is_0_o , \PWM6/n4_neg , \PWM6/n6_neg );
  AL_MUX \PWM6/u9  (
    .i0(\PWM6/n8 ),
    .i1(1'b1),
    .sel(pwm_start_stop[22]),
    .o(\PWM6/n9 ));  // src/OnePWM.v(26)
  reg_ar_as_w1 \PWM7/State_reg  (
    .clk(clk100m),
    .d(\PWM7/n10 ),
    .en(1'b1),
    .reset(~rstn),
    .set(1'b0),
    .q(pwm_state_read[7]));  // src/OnePWM.v(26)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[0]  (
    .i(\PWM7/RemaTxNum[0]_keep ),
    .o(pnumcnt7[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[10]  (
    .i(\PWM7/RemaTxNum[10]_keep ),
    .o(pnumcnt7[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[11]  (
    .i(\PWM7/RemaTxNum[11]_keep ),
    .o(pnumcnt7[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[12]  (
    .i(\PWM7/RemaTxNum[12]_keep ),
    .o(pnumcnt7[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[13]  (
    .i(\PWM7/RemaTxNum[13]_keep ),
    .o(pnumcnt7[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[14]  (
    .i(\PWM7/RemaTxNum[14]_keep ),
    .o(pnumcnt7[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[15]  (
    .i(\PWM7/RemaTxNum[15]_keep ),
    .o(pnumcnt7[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[16]  (
    .i(\PWM7/RemaTxNum[16]_keep ),
    .o(pnumcnt7[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[17]  (
    .i(\PWM7/RemaTxNum[17]_keep ),
    .o(pnumcnt7[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[18]  (
    .i(\PWM7/RemaTxNum[18]_keep ),
    .o(pnumcnt7[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[19]  (
    .i(\PWM7/RemaTxNum[19]_keep ),
    .o(pnumcnt7[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[1]  (
    .i(\PWM7/RemaTxNum[1]_keep ),
    .o(pnumcnt7[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[20]  (
    .i(\PWM7/RemaTxNum[20]_keep ),
    .o(pnumcnt7[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[21]  (
    .i(\PWM7/RemaTxNum[21]_keep ),
    .o(pnumcnt7[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[22]  (
    .i(\PWM7/RemaTxNum[22]_keep ),
    .o(pnumcnt7[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[23]  (
    .i(\PWM7/RemaTxNum[23]_keep ),
    .o(pnumcnt7[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[2]  (
    .i(\PWM7/RemaTxNum[2]_keep ),
    .o(pnumcnt7[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[3]  (
    .i(\PWM7/RemaTxNum[3]_keep ),
    .o(pnumcnt7[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[4]  (
    .i(\PWM7/RemaTxNum[4]_keep ),
    .o(pnumcnt7[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[5]  (
    .i(\PWM7/RemaTxNum[5]_keep ),
    .o(pnumcnt7[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[6]  (
    .i(\PWM7/RemaTxNum[6]_keep ),
    .o(pnumcnt7[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[7]  (
    .i(\PWM7/RemaTxNum[7]_keep ),
    .o(pnumcnt7[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[8]  (
    .i(\PWM7/RemaTxNum[8]_keep ),
    .o(pnumcnt7[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_RemaTxNum[9]  (
    .i(\PWM7/RemaTxNum[9]_keep ),
    .o(pnumcnt7[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_dir  (
    .i(\PWM7/dir_keep ),
    .o(dir[7]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[0]  (
    .i(\PWM7/pnumr[0]_keep ),
    .o(\PWM7/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[10]  (
    .i(\PWM7/pnumr[10]_keep ),
    .o(\PWM7/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[11]  (
    .i(\PWM7/pnumr[11]_keep ),
    .o(\PWM7/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[12]  (
    .i(\PWM7/pnumr[12]_keep ),
    .o(\PWM7/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[13]  (
    .i(\PWM7/pnumr[13]_keep ),
    .o(\PWM7/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[14]  (
    .i(\PWM7/pnumr[14]_keep ),
    .o(\PWM7/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[15]  (
    .i(\PWM7/pnumr[15]_keep ),
    .o(\PWM7/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[16]  (
    .i(\PWM7/pnumr[16]_keep ),
    .o(\PWM7/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[17]  (
    .i(\PWM7/pnumr[17]_keep ),
    .o(\PWM7/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[18]  (
    .i(\PWM7/pnumr[18]_keep ),
    .o(\PWM7/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[19]  (
    .i(\PWM7/pnumr[19]_keep ),
    .o(\PWM7/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[1]  (
    .i(\PWM7/pnumr[1]_keep ),
    .o(\PWM7/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[20]  (
    .i(\PWM7/pnumr[20]_keep ),
    .o(\PWM7/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[21]  (
    .i(\PWM7/pnumr[21]_keep ),
    .o(\PWM7/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[22]  (
    .i(\PWM7/pnumr[22]_keep ),
    .o(\PWM7/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[23]  (
    .i(\PWM7/pnumr[23]_keep ),
    .o(\PWM7/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[24]  (
    .i(\PWM7/pnumr[24]_keep ),
    .o(\PWM7/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[25]  (
    .i(\PWM7/pnumr[25]_keep ),
    .o(\PWM7/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[26]  (
    .i(\PWM7/pnumr[26]_keep ),
    .o(\PWM7/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[27]  (
    .i(\PWM7/pnumr[27]_keep ),
    .o(\PWM7/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[28]  (
    .i(\PWM7/pnumr[28]_keep ),
    .o(\PWM7/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[29]  (
    .i(\PWM7/pnumr[29]_keep ),
    .o(\PWM7/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[2]  (
    .i(\PWM7/pnumr[2]_keep ),
    .o(\PWM7/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[30]  (
    .i(\PWM7/pnumr[30]_keep ),
    .o(\PWM7/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[31]  (
    .i(\PWM7/pnumr[31]_keep ),
    .o(\PWM7/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[3]  (
    .i(\PWM7/pnumr[3]_keep ),
    .o(\PWM7/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[4]  (
    .i(\PWM7/pnumr[4]_keep ),
    .o(\PWM7/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[5]  (
    .i(\PWM7/pnumr[5]_keep ),
    .o(\PWM7/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[6]  (
    .i(\PWM7/pnumr[6]_keep ),
    .o(\PWM7/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[7]  (
    .i(\PWM7/pnumr[7]_keep ),
    .o(\PWM7/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[8]  (
    .i(\PWM7/pnumr[8]_keep ),
    .o(\PWM7/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pnumr[9]  (
    .i(\PWM7/pnumr[9]_keep ),
    .o(\PWM7/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_pwm  (
    .i(\PWM7/pwm_keep ),
    .o(pwm[7]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM7/_bufkeep_stopreq  (
    .i(\PWM7/stopreq_keep ),
    .o(\PWM7/stopreq ));  // src/OnePWM.v(14)
  reg_ar_as_w1 \PWM7/dir_reg  (
    .clk(clk100m),
    .d(\PWM7/n32 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/dir_keep ));  // src/OnePWM.v(58)
  eq_w27 \PWM7/eq0  (
    .i0(\PWM7/FreCnt ),
    .i1(27'b000000000000000000000000000),
    .o(\PWM7/n0 ));  // src/OnePWM.v(15)
  eq_w24 \PWM7/eq1  (
    .i0(pnumcnt7),
    .i1(24'b000000000000000000000001),
    .o(\PWM7/n5 ));  // src/OnePWM.v(25)
  eq_w27 \PWM7/eq2  (
    .i0(\PWM7/FreCnt ),
    .i1({1'b0,\PWM7/FreCntr [26:1]}),
    .o(\PWM7/n17 ));  // src/OnePWM.v(41)
  eq_w27 \PWM7/eq3  (
    .i0(\PWM7/FreCnt ),
    .i1(\PWM7/FreCntr ),
    .o(\PWM7/n18 ));  // src/OnePWM.v(43)
  binary_mux_s1_w1 \PWM7/mux0_b0  (
    .i0(\PWM7/n12 [0]),
    .i1(freq7[0]),
    .sel(\PWM7/n0 ),
    .o(\PWM7/n13 [0]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM7/mux0_b1  (
    .i0(\PWM7/n12 [1]),
    .i1(freq7[1]),
    .sel(\PWM7/n0 ),
    .o(\PWM7/n13 [1]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM7/mux0_b10  (
    .i0(\PWM7/n12 [10]),
    .i1(freq7[10]),
    .sel(\PWM7/n0 ),
    .o(\PWM7/n13 [10]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM7/mux0_b11  (
    .i0(\PWM7/n12 [11]),
    .i1(freq7[11]),
    .sel(\PWM7/n0 ),
    .o(\PWM7/n13 [11]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM7/mux0_b12  (
    .i0(\PWM7/n12 [12]),
    .i1(freq7[12]),
    .sel(\PWM7/n0 ),
    .o(\PWM7/n13 [12]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM7/mux0_b13  (
    .i0(\PWM7/n12 [13]),
    .i1(freq7[13]),
    .sel(\PWM7/n0 ),
    .o(\PWM7/n13 [13]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM7/mux0_b14  (
    .i0(\PWM7/n12 [14]),
    .i1(freq7[14]),
    .sel(\PWM7/n0 ),
    .o(\PWM7/n13 [14]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM7/mux0_b15  (
    .i0(\PWM7/n12 [15]),
    .i1(freq7[15]),
    .sel(\PWM7/n0 ),
    .o(\PWM7/n13 [15]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM7/mux0_b16  (
    .i0(\PWM7/n12 [16]),
    .i1(freq7[16]),
    .sel(\PWM7/n0 ),
    .o(\PWM7/n13 [16]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM7/mux0_b17  (
    .i0(\PWM7/n12 [17]),
    .i1(freq7[17]),
    .sel(\PWM7/n0 ),
    .o(\PWM7/n13 [17]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM7/mux0_b18  (
    .i0(\PWM7/n12 [18]),
    .i1(freq7[18]),
    .sel(\PWM7/n0 ),
    .o(\PWM7/n13 [18]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM7/mux0_b19  (
    .i0(\PWM7/n12 [19]),
    .i1(freq7[19]),
    .sel(\PWM7/n0 ),
    .o(\PWM7/n13 [19]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM7/mux0_b2  (
    .i0(\PWM7/n12 [2]),
    .i1(freq7[2]),
    .sel(\PWM7/n0 ),
    .o(\PWM7/n13 [2]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM7/mux0_b20  (
    .i0(\PWM7/n12 [20]),
    .i1(freq7[20]),
    .sel(\PWM7/n0 ),
    .o(\PWM7/n13 [20]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM7/mux0_b21  (
    .i0(\PWM7/n12 [21]),
    .i1(freq7[21]),
    .sel(\PWM7/n0 ),
    .o(\PWM7/n13 [21]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM7/mux0_b22  (
    .i0(\PWM7/n12 [22]),
    .i1(freq7[22]),
    .sel(\PWM7/n0 ),
    .o(\PWM7/n13 [22]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM7/mux0_b23  (
    .i0(\PWM7/n12 [23]),
    .i1(freq7[23]),
    .sel(\PWM7/n0 ),
    .o(\PWM7/n13 [23]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM7/mux0_b24  (
    .i0(\PWM7/n12 [24]),
    .i1(freq7[24]),
    .sel(\PWM7/n0 ),
    .o(\PWM7/n13 [24]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM7/mux0_b25  (
    .i0(\PWM7/n12 [25]),
    .i1(freq7[25]),
    .sel(\PWM7/n0 ),
    .o(\PWM7/n13 [25]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM7/mux0_b26  (
    .i0(\PWM7/n12 [26]),
    .i1(freq7[26]),
    .sel(\PWM7/n0 ),
    .o(\PWM7/n13 [26]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM7/mux0_b3  (
    .i0(\PWM7/n12 [3]),
    .i1(freq7[3]),
    .sel(\PWM7/n0 ),
    .o(\PWM7/n13 [3]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM7/mux0_b4  (
    .i0(\PWM7/n12 [4]),
    .i1(freq7[4]),
    .sel(\PWM7/n0 ),
    .o(\PWM7/n13 [4]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM7/mux0_b5  (
    .i0(\PWM7/n12 [5]),
    .i1(freq7[5]),
    .sel(\PWM7/n0 ),
    .o(\PWM7/n13 [5]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM7/mux0_b6  (
    .i0(\PWM7/n12 [6]),
    .i1(freq7[6]),
    .sel(\PWM7/n0 ),
    .o(\PWM7/n13 [6]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM7/mux0_b7  (
    .i0(\PWM7/n12 [7]),
    .i1(freq7[7]),
    .sel(\PWM7/n0 ),
    .o(\PWM7/n13 [7]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM7/mux0_b8  (
    .i0(\PWM7/n12 [8]),
    .i1(freq7[8]),
    .sel(\PWM7/n0 ),
    .o(\PWM7/n13 [8]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM7/mux0_b9  (
    .i0(\PWM7/n12 [9]),
    .i1(freq7[9]),
    .sel(\PWM7/n0 ),
    .o(\PWM7/n13 [9]));  // src/OnePWM.v(32)
  and \PWM7/mux3_b0_sel_is_3  (\PWM7/mux3_b0_sel_is_3_o , \PWM7/n11 , \PWM7/n0 );
  binary_mux_s1_w1 \PWM7/mux4_b0  (
    .i0(\PWM7/pnumr [0]),
    .i1(1'b0),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n22 [0]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux4_b1  (
    .i0(\PWM7/pnumr [1]),
    .i1(1'b0),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n22 [1]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux4_b10  (
    .i0(\PWM7/pnumr [10]),
    .i1(1'b0),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n22 [10]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux4_b11  (
    .i0(\PWM7/pnumr [11]),
    .i1(1'b0),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n22 [11]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux4_b12  (
    .i0(\PWM7/pnumr [12]),
    .i1(1'b0),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n22 [12]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux4_b13  (
    .i0(\PWM7/pnumr [13]),
    .i1(1'b0),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n22 [13]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux4_b14  (
    .i0(\PWM7/pnumr [14]),
    .i1(1'b0),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n22 [14]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux4_b15  (
    .i0(\PWM7/pnumr [15]),
    .i1(1'b0),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n22 [15]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux4_b16  (
    .i0(\PWM7/pnumr [16]),
    .i1(1'b0),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n22 [16]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux4_b17  (
    .i0(\PWM7/pnumr [17]),
    .i1(1'b0),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n22 [17]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux4_b18  (
    .i0(\PWM7/pnumr [18]),
    .i1(1'b0),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n22 [18]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux4_b19  (
    .i0(\PWM7/pnumr [19]),
    .i1(1'b0),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n22 [19]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux4_b2  (
    .i0(\PWM7/pnumr [2]),
    .i1(1'b0),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n22 [2]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux4_b20  (
    .i0(\PWM7/pnumr [20]),
    .i1(1'b0),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n22 [20]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux4_b21  (
    .i0(\PWM7/pnumr [21]),
    .i1(1'b0),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n22 [21]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux4_b22  (
    .i0(\PWM7/pnumr [22]),
    .i1(1'b0),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n22 [22]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux4_b23  (
    .i0(\PWM7/pnumr [23]),
    .i1(1'b0),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n22 [23]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux4_b24  (
    .i0(\PWM7/pnumr [24]),
    .i1(1'b0),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n22 [24]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux4_b25  (
    .i0(\PWM7/pnumr [25]),
    .i1(1'b0),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n22 [25]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux4_b26  (
    .i0(\PWM7/pnumr [26]),
    .i1(1'b0),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n22 [26]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux4_b27  (
    .i0(\PWM7/pnumr [27]),
    .i1(1'b0),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n22 [27]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux4_b28  (
    .i0(\PWM7/pnumr [28]),
    .i1(1'b0),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n22 [28]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux4_b29  (
    .i0(\PWM7/pnumr [29]),
    .i1(1'b0),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n22 [29]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux4_b3  (
    .i0(\PWM7/pnumr [3]),
    .i1(1'b0),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n22 [3]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux4_b30  (
    .i0(\PWM7/pnumr [30]),
    .i1(1'b0),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n22 [30]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux4_b31  (
    .i0(\PWM7/pnumr [31]),
    .i1(1'b0),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n22 [31]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux4_b4  (
    .i0(\PWM7/pnumr [4]),
    .i1(1'b0),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n22 [4]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux4_b5  (
    .i0(\PWM7/pnumr [5]),
    .i1(1'b0),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n22 [5]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux4_b6  (
    .i0(\PWM7/pnumr [6]),
    .i1(1'b0),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n22 [6]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux4_b7  (
    .i0(\PWM7/pnumr [7]),
    .i1(1'b0),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n22 [7]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux4_b8  (
    .i0(\PWM7/pnumr [8]),
    .i1(1'b0),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n22 [8]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux4_b9  (
    .i0(\PWM7/pnumr [9]),
    .i1(1'b0),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n22 [9]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux5_b0  (
    .i0(\PWM7/n22 [0]),
    .i1(pnum7[0]),
    .sel(pnum7[32]),
    .o(\PWM7/n23 [0]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux5_b1  (
    .i0(\PWM7/n22 [1]),
    .i1(pnum7[1]),
    .sel(pnum7[32]),
    .o(\PWM7/n23 [1]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux5_b10  (
    .i0(\PWM7/n22 [10]),
    .i1(pnum7[10]),
    .sel(pnum7[32]),
    .o(\PWM7/n23 [10]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux5_b11  (
    .i0(\PWM7/n22 [11]),
    .i1(pnum7[11]),
    .sel(pnum7[32]),
    .o(\PWM7/n23 [11]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux5_b12  (
    .i0(\PWM7/n22 [12]),
    .i1(pnum7[12]),
    .sel(pnum7[32]),
    .o(\PWM7/n23 [12]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux5_b13  (
    .i0(\PWM7/n22 [13]),
    .i1(pnum7[13]),
    .sel(pnum7[32]),
    .o(\PWM7/n23 [13]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux5_b14  (
    .i0(\PWM7/n22 [14]),
    .i1(pnum7[14]),
    .sel(pnum7[32]),
    .o(\PWM7/n23 [14]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux5_b15  (
    .i0(\PWM7/n22 [15]),
    .i1(pnum7[15]),
    .sel(pnum7[32]),
    .o(\PWM7/n23 [15]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux5_b16  (
    .i0(\PWM7/n22 [16]),
    .i1(pnum7[16]),
    .sel(pnum7[32]),
    .o(\PWM7/n23 [16]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux5_b17  (
    .i0(\PWM7/n22 [17]),
    .i1(pnum7[17]),
    .sel(pnum7[32]),
    .o(\PWM7/n23 [17]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux5_b18  (
    .i0(\PWM7/n22 [18]),
    .i1(pnum7[18]),
    .sel(pnum7[32]),
    .o(\PWM7/n23 [18]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux5_b19  (
    .i0(\PWM7/n22 [19]),
    .i1(pnum7[19]),
    .sel(pnum7[32]),
    .o(\PWM7/n23 [19]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux5_b2  (
    .i0(\PWM7/n22 [2]),
    .i1(pnum7[2]),
    .sel(pnum7[32]),
    .o(\PWM7/n23 [2]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux5_b20  (
    .i0(\PWM7/n22 [20]),
    .i1(pnum7[20]),
    .sel(pnum7[32]),
    .o(\PWM7/n23 [20]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux5_b21  (
    .i0(\PWM7/n22 [21]),
    .i1(pnum7[21]),
    .sel(pnum7[32]),
    .o(\PWM7/n23 [21]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux5_b22  (
    .i0(\PWM7/n22 [22]),
    .i1(pnum7[22]),
    .sel(pnum7[32]),
    .o(\PWM7/n23 [22]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux5_b23  (
    .i0(\PWM7/n22 [23]),
    .i1(pnum7[23]),
    .sel(pnum7[32]),
    .o(\PWM7/n23 [23]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux5_b24  (
    .i0(\PWM7/n22 [24]),
    .i1(pnum7[24]),
    .sel(pnum7[32]),
    .o(\PWM7/n23 [24]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux5_b25  (
    .i0(\PWM7/n22 [25]),
    .i1(pnum7[25]),
    .sel(pnum7[32]),
    .o(\PWM7/n23 [25]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux5_b26  (
    .i0(\PWM7/n22 [26]),
    .i1(pnum7[26]),
    .sel(pnum7[32]),
    .o(\PWM7/n23 [26]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux5_b27  (
    .i0(\PWM7/n22 [27]),
    .i1(pnum7[27]),
    .sel(pnum7[32]),
    .o(\PWM7/n23 [27]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux5_b28  (
    .i0(\PWM7/n22 [28]),
    .i1(pnum7[28]),
    .sel(pnum7[32]),
    .o(\PWM7/n23 [28]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux5_b29  (
    .i0(\PWM7/n22 [29]),
    .i1(pnum7[29]),
    .sel(pnum7[32]),
    .o(\PWM7/n23 [29]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux5_b3  (
    .i0(\PWM7/n22 [3]),
    .i1(pnum7[3]),
    .sel(pnum7[32]),
    .o(\PWM7/n23 [3]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux5_b30  (
    .i0(\PWM7/n22 [30]),
    .i1(pnum7[30]),
    .sel(pnum7[32]),
    .o(\PWM7/n23 [30]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux5_b31  (
    .i0(\PWM7/n22 [31]),
    .i1(pnum7[31]),
    .sel(pnum7[32]),
    .o(\PWM7/n23 [31]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux5_b4  (
    .i0(\PWM7/n22 [4]),
    .i1(pnum7[4]),
    .sel(pnum7[32]),
    .o(\PWM7/n23 [4]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux5_b5  (
    .i0(\PWM7/n22 [5]),
    .i1(pnum7[5]),
    .sel(pnum7[32]),
    .o(\PWM7/n23 [5]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux5_b6  (
    .i0(\PWM7/n22 [6]),
    .i1(pnum7[6]),
    .sel(pnum7[32]),
    .o(\PWM7/n23 [6]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux5_b7  (
    .i0(\PWM7/n22 [7]),
    .i1(pnum7[7]),
    .sel(pnum7[32]),
    .o(\PWM7/n23 [7]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux5_b8  (
    .i0(\PWM7/n22 [8]),
    .i1(pnum7[8]),
    .sel(pnum7[32]),
    .o(\PWM7/n23 [8]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux5_b9  (
    .i0(\PWM7/n22 [9]),
    .i1(pnum7[9]),
    .sel(pnum7[32]),
    .o(\PWM7/n23 [9]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM7/mux6_b0  (
    .i0(\PWM7/pnumr [0]),
    .i1(\PWM7/n26 [0]),
    .sel(\PWM7/n25 ),
    .o(\PWM7/n27 [0]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM7/mux6_b1  (
    .i0(\PWM7/pnumr [1]),
    .i1(\PWM7/n26 [1]),
    .sel(\PWM7/n25 ),
    .o(\PWM7/n27 [1]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM7/mux6_b10  (
    .i0(\PWM7/pnumr [10]),
    .i1(\PWM7/n26 [10]),
    .sel(\PWM7/n25 ),
    .o(\PWM7/n27 [10]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM7/mux6_b11  (
    .i0(\PWM7/pnumr [11]),
    .i1(\PWM7/n26 [11]),
    .sel(\PWM7/n25 ),
    .o(\PWM7/n27 [11]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM7/mux6_b12  (
    .i0(\PWM7/pnumr [12]),
    .i1(\PWM7/n26 [12]),
    .sel(\PWM7/n25 ),
    .o(\PWM7/n27 [12]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM7/mux6_b13  (
    .i0(\PWM7/pnumr [13]),
    .i1(\PWM7/n26 [13]),
    .sel(\PWM7/n25 ),
    .o(\PWM7/n27 [13]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM7/mux6_b14  (
    .i0(\PWM7/pnumr [14]),
    .i1(\PWM7/n26 [14]),
    .sel(\PWM7/n25 ),
    .o(\PWM7/n27 [14]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM7/mux6_b15  (
    .i0(\PWM7/pnumr [15]),
    .i1(\PWM7/n26 [15]),
    .sel(\PWM7/n25 ),
    .o(\PWM7/n27 [15]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM7/mux6_b16  (
    .i0(\PWM7/pnumr [16]),
    .i1(\PWM7/n26 [16]),
    .sel(\PWM7/n25 ),
    .o(\PWM7/n27 [16]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM7/mux6_b17  (
    .i0(\PWM7/pnumr [17]),
    .i1(\PWM7/n26 [17]),
    .sel(\PWM7/n25 ),
    .o(\PWM7/n27 [17]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM7/mux6_b18  (
    .i0(\PWM7/pnumr [18]),
    .i1(\PWM7/n26 [18]),
    .sel(\PWM7/n25 ),
    .o(\PWM7/n27 [18]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM7/mux6_b19  (
    .i0(\PWM7/pnumr [19]),
    .i1(\PWM7/n26 [19]),
    .sel(\PWM7/n25 ),
    .o(\PWM7/n27 [19]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM7/mux6_b2  (
    .i0(\PWM7/pnumr [2]),
    .i1(\PWM7/n26 [2]),
    .sel(\PWM7/n25 ),
    .o(\PWM7/n27 [2]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM7/mux6_b20  (
    .i0(\PWM7/pnumr [20]),
    .i1(\PWM7/n26 [20]),
    .sel(\PWM7/n25 ),
    .o(\PWM7/n27 [20]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM7/mux6_b21  (
    .i0(\PWM7/pnumr [21]),
    .i1(\PWM7/n26 [21]),
    .sel(\PWM7/n25 ),
    .o(\PWM7/n27 [21]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM7/mux6_b22  (
    .i0(\PWM7/pnumr [22]),
    .i1(\PWM7/n26 [22]),
    .sel(\PWM7/n25 ),
    .o(\PWM7/n27 [22]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM7/mux6_b23  (
    .i0(\PWM7/pnumr [23]),
    .i1(\PWM7/n26 [23]),
    .sel(\PWM7/n25 ),
    .o(\PWM7/n27 [23]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM7/mux6_b3  (
    .i0(\PWM7/pnumr [3]),
    .i1(\PWM7/n26 [3]),
    .sel(\PWM7/n25 ),
    .o(\PWM7/n27 [3]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM7/mux6_b4  (
    .i0(\PWM7/pnumr [4]),
    .i1(\PWM7/n26 [4]),
    .sel(\PWM7/n25 ),
    .o(\PWM7/n27 [4]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM7/mux6_b5  (
    .i0(\PWM7/pnumr [5]),
    .i1(\PWM7/n26 [5]),
    .sel(\PWM7/n25 ),
    .o(\PWM7/n27 [5]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM7/mux6_b6  (
    .i0(\PWM7/pnumr [6]),
    .i1(\PWM7/n26 [6]),
    .sel(\PWM7/n25 ),
    .o(\PWM7/n27 [6]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM7/mux6_b7  (
    .i0(\PWM7/pnumr [7]),
    .i1(\PWM7/n26 [7]),
    .sel(\PWM7/n25 ),
    .o(\PWM7/n27 [7]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM7/mux6_b8  (
    .i0(\PWM7/pnumr [8]),
    .i1(\PWM7/n26 [8]),
    .sel(\PWM7/n25 ),
    .o(\PWM7/n27 [8]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM7/mux6_b9  (
    .i0(\PWM7/pnumr [9]),
    .i1(\PWM7/n26 [9]),
    .sel(\PWM7/n25 ),
    .o(\PWM7/n27 [9]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM7/mux7_b0  (
    .i0(pnumcnt7[0]),
    .i1(\PWM7/n27 [0]),
    .sel(\PWM7/n24 ),
    .o(\PWM7/n29 [0]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux7_b1  (
    .i0(pnumcnt7[1]),
    .i1(\PWM7/n27 [1]),
    .sel(\PWM7/n24 ),
    .o(\PWM7/n29 [1]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux7_b10  (
    .i0(pnumcnt7[10]),
    .i1(\PWM7/n27 [10]),
    .sel(\PWM7/n24 ),
    .o(\PWM7/n29 [10]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux7_b11  (
    .i0(pnumcnt7[11]),
    .i1(\PWM7/n27 [11]),
    .sel(\PWM7/n24 ),
    .o(\PWM7/n29 [11]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux7_b12  (
    .i0(pnumcnt7[12]),
    .i1(\PWM7/n27 [12]),
    .sel(\PWM7/n24 ),
    .o(\PWM7/n29 [12]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux7_b13  (
    .i0(pnumcnt7[13]),
    .i1(\PWM7/n27 [13]),
    .sel(\PWM7/n24 ),
    .o(\PWM7/n29 [13]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux7_b14  (
    .i0(pnumcnt7[14]),
    .i1(\PWM7/n27 [14]),
    .sel(\PWM7/n24 ),
    .o(\PWM7/n29 [14]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux7_b15  (
    .i0(pnumcnt7[15]),
    .i1(\PWM7/n27 [15]),
    .sel(\PWM7/n24 ),
    .o(\PWM7/n29 [15]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux7_b16  (
    .i0(pnumcnt7[16]),
    .i1(\PWM7/n27 [16]),
    .sel(\PWM7/n24 ),
    .o(\PWM7/n29 [16]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux7_b17  (
    .i0(pnumcnt7[17]),
    .i1(\PWM7/n27 [17]),
    .sel(\PWM7/n24 ),
    .o(\PWM7/n29 [17]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux7_b18  (
    .i0(pnumcnt7[18]),
    .i1(\PWM7/n27 [18]),
    .sel(\PWM7/n24 ),
    .o(\PWM7/n29 [18]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux7_b19  (
    .i0(pnumcnt7[19]),
    .i1(\PWM7/n27 [19]),
    .sel(\PWM7/n24 ),
    .o(\PWM7/n29 [19]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux7_b2  (
    .i0(pnumcnt7[2]),
    .i1(\PWM7/n27 [2]),
    .sel(\PWM7/n24 ),
    .o(\PWM7/n29 [2]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux7_b20  (
    .i0(pnumcnt7[20]),
    .i1(\PWM7/n27 [20]),
    .sel(\PWM7/n24 ),
    .o(\PWM7/n29 [20]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux7_b21  (
    .i0(pnumcnt7[21]),
    .i1(\PWM7/n27 [21]),
    .sel(\PWM7/n24 ),
    .o(\PWM7/n29 [21]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux7_b22  (
    .i0(pnumcnt7[22]),
    .i1(\PWM7/n27 [22]),
    .sel(\PWM7/n24 ),
    .o(\PWM7/n29 [22]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux7_b23  (
    .i0(pnumcnt7[23]),
    .i1(\PWM7/n27 [23]),
    .sel(\PWM7/n24 ),
    .o(\PWM7/n29 [23]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux7_b3  (
    .i0(pnumcnt7[3]),
    .i1(\PWM7/n27 [3]),
    .sel(\PWM7/n24 ),
    .o(\PWM7/n29 [3]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux7_b4  (
    .i0(pnumcnt7[4]),
    .i1(\PWM7/n27 [4]),
    .sel(\PWM7/n24 ),
    .o(\PWM7/n29 [4]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux7_b5  (
    .i0(pnumcnt7[5]),
    .i1(\PWM7/n27 [5]),
    .sel(\PWM7/n24 ),
    .o(\PWM7/n29 [5]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux7_b6  (
    .i0(pnumcnt7[6]),
    .i1(\PWM7/n27 [6]),
    .sel(\PWM7/n24 ),
    .o(\PWM7/n29 [6]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux7_b7  (
    .i0(pnumcnt7[7]),
    .i1(\PWM7/n27 [7]),
    .sel(\PWM7/n24 ),
    .o(\PWM7/n29 [7]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux7_b8  (
    .i0(pnumcnt7[8]),
    .i1(\PWM7/n27 [8]),
    .sel(\PWM7/n24 ),
    .o(\PWM7/n29 [8]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux7_b9  (
    .i0(pnumcnt7[9]),
    .i1(\PWM7/n27 [9]),
    .sel(\PWM7/n24 ),
    .o(\PWM7/n29 [9]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux8_b0  (
    .i0(\PWM7/n29 [0]),
    .i1(\PWM7/pnumr [0]),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n31 [0]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux8_b1  (
    .i0(\PWM7/n29 [1]),
    .i1(\PWM7/pnumr [1]),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n31 [1]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux8_b10  (
    .i0(\PWM7/n29 [10]),
    .i1(\PWM7/pnumr [10]),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n31 [10]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux8_b11  (
    .i0(\PWM7/n29 [11]),
    .i1(\PWM7/pnumr [11]),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n31 [11]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux8_b12  (
    .i0(\PWM7/n29 [12]),
    .i1(\PWM7/pnumr [12]),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n31 [12]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux8_b13  (
    .i0(\PWM7/n29 [13]),
    .i1(\PWM7/pnumr [13]),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n31 [13]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux8_b14  (
    .i0(\PWM7/n29 [14]),
    .i1(\PWM7/pnumr [14]),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n31 [14]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux8_b15  (
    .i0(\PWM7/n29 [15]),
    .i1(\PWM7/pnumr [15]),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n31 [15]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux8_b16  (
    .i0(\PWM7/n29 [16]),
    .i1(\PWM7/pnumr [16]),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n31 [16]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux8_b17  (
    .i0(\PWM7/n29 [17]),
    .i1(\PWM7/pnumr [17]),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n31 [17]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux8_b18  (
    .i0(\PWM7/n29 [18]),
    .i1(\PWM7/pnumr [18]),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n31 [18]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux8_b19  (
    .i0(\PWM7/n29 [19]),
    .i1(\PWM7/pnumr [19]),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n31 [19]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux8_b2  (
    .i0(\PWM7/n29 [2]),
    .i1(\PWM7/pnumr [2]),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n31 [2]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux8_b20  (
    .i0(\PWM7/n29 [20]),
    .i1(\PWM7/pnumr [20]),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n31 [20]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux8_b21  (
    .i0(\PWM7/n29 [21]),
    .i1(\PWM7/pnumr [21]),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n31 [21]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux8_b22  (
    .i0(\PWM7/n29 [22]),
    .i1(\PWM7/pnumr [22]),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n31 [22]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux8_b23  (
    .i0(\PWM7/n29 [23]),
    .i1(\PWM7/pnumr [23]),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n31 [23]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux8_b3  (
    .i0(\PWM7/n29 [3]),
    .i1(\PWM7/pnumr [3]),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n31 [3]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux8_b4  (
    .i0(\PWM7/n29 [4]),
    .i1(\PWM7/pnumr [4]),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n31 [4]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux8_b5  (
    .i0(\PWM7/n29 [5]),
    .i1(\PWM7/pnumr [5]),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n31 [5]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux8_b6  (
    .i0(\PWM7/n29 [6]),
    .i1(\PWM7/pnumr [6]),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n31 [6]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux8_b7  (
    .i0(\PWM7/n29 [7]),
    .i1(\PWM7/pnumr [7]),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n31 [7]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux8_b8  (
    .i0(\PWM7/n29 [8]),
    .i1(\PWM7/pnumr [8]),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n31 [8]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM7/mux8_b9  (
    .i0(\PWM7/n29 [9]),
    .i1(\PWM7/pnumr [9]),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n31 [9]));  // src/OnePWM.v(57)
  not \PWM7/n17_inv  (\PWM7/n17_neg , \PWM7/n17 );
  not \PWM7/n25_inv  (\PWM7/n25_neg , \PWM7/n25 );
  not \PWM7/n4_inv  (\PWM7/n4_neg , \PWM7/n4 );
  not \PWM7/n6_inv  (\PWM7/n6_neg , \PWM7/n6 );
  ne_w24 \PWM7/neq0  (
    .i0(pnumcnt7),
    .i1(24'b000000000000000000000000),
    .o(\PWM7/n25 ));  // src/OnePWM.v(55)
  reg_sr_ss_w1 \PWM7/pwm_reg  (
    .clk(clk100m),
    .d(pwm[7]),
    .en(1'b1),
    .reset(~\PWM7/u14_sel_is_1_o ),
    .set(\PWM7/n18 ),
    .q(\PWM7/pwm_keep ));  // src/OnePWM.v(45)
  reg_sr_as_w1 \PWM7/reg0_b0  (
    .clk(clk100m),
    .d(\PWM7/n13 [0]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [0]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b1  (
    .clk(clk100m),
    .d(\PWM7/n13 [1]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [1]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b10  (
    .clk(clk100m),
    .d(\PWM7/n13 [10]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [10]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b11  (
    .clk(clk100m),
    .d(\PWM7/n13 [11]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [11]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b12  (
    .clk(clk100m),
    .d(\PWM7/n13 [12]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [12]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b13  (
    .clk(clk100m),
    .d(\PWM7/n13 [13]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [13]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b14  (
    .clk(clk100m),
    .d(\PWM7/n13 [14]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [14]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b15  (
    .clk(clk100m),
    .d(\PWM7/n13 [15]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [15]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b16  (
    .clk(clk100m),
    .d(\PWM7/n13 [16]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [16]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b17  (
    .clk(clk100m),
    .d(\PWM7/n13 [17]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [17]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b18  (
    .clk(clk100m),
    .d(\PWM7/n13 [18]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [18]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b19  (
    .clk(clk100m),
    .d(\PWM7/n13 [19]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [19]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b2  (
    .clk(clk100m),
    .d(\PWM7/n13 [2]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [2]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b20  (
    .clk(clk100m),
    .d(\PWM7/n13 [20]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [20]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b21  (
    .clk(clk100m),
    .d(\PWM7/n13 [21]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [21]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b22  (
    .clk(clk100m),
    .d(\PWM7/n13 [22]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [22]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b23  (
    .clk(clk100m),
    .d(\PWM7/n13 [23]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [23]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b24  (
    .clk(clk100m),
    .d(\PWM7/n13 [24]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [24]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b25  (
    .clk(clk100m),
    .d(\PWM7/n13 [25]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [25]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b26  (
    .clk(clk100m),
    .d(\PWM7/n13 [26]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [26]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b3  (
    .clk(clk100m),
    .d(\PWM7/n13 [3]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [3]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b4  (
    .clk(clk100m),
    .d(\PWM7/n13 [4]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [4]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b5  (
    .clk(clk100m),
    .d(\PWM7/n13 [5]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [5]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b6  (
    .clk(clk100m),
    .d(\PWM7/n13 [6]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [6]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b7  (
    .clk(clk100m),
    .d(\PWM7/n13 [7]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [7]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b8  (
    .clk(clk100m),
    .d(\PWM7/n13 [8]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [8]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM7/reg0_b9  (
    .clk(clk100m),
    .d(\PWM7/n13 [9]),
    .en(1'b1),
    .reset(~\PWM7/n11 ),
    .set(1'b0),
    .q(\PWM7/FreCnt [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b0  (
    .clk(clk100m),
    .d(freq7[0]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [0]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b1  (
    .clk(clk100m),
    .d(freq7[1]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [1]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b10  (
    .clk(clk100m),
    .d(freq7[10]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [10]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b11  (
    .clk(clk100m),
    .d(freq7[11]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [11]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b12  (
    .clk(clk100m),
    .d(freq7[12]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [12]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b13  (
    .clk(clk100m),
    .d(freq7[13]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [13]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b14  (
    .clk(clk100m),
    .d(freq7[14]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [14]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b15  (
    .clk(clk100m),
    .d(freq7[15]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [15]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b16  (
    .clk(clk100m),
    .d(freq7[16]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [16]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b17  (
    .clk(clk100m),
    .d(freq7[17]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [17]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b18  (
    .clk(clk100m),
    .d(freq7[18]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [18]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b19  (
    .clk(clk100m),
    .d(freq7[19]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [19]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b2  (
    .clk(clk100m),
    .d(freq7[2]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [2]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b20  (
    .clk(clk100m),
    .d(freq7[20]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [20]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b21  (
    .clk(clk100m),
    .d(freq7[21]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [21]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b22  (
    .clk(clk100m),
    .d(freq7[22]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [22]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b23  (
    .clk(clk100m),
    .d(freq7[23]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [23]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b24  (
    .clk(clk100m),
    .d(freq7[24]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [24]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b25  (
    .clk(clk100m),
    .d(freq7[25]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [25]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b26  (
    .clk(clk100m),
    .d(freq7[26]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [26]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b3  (
    .clk(clk100m),
    .d(freq7[3]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [3]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b4  (
    .clk(clk100m),
    .d(freq7[4]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [4]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b5  (
    .clk(clk100m),
    .d(freq7[5]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [5]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b6  (
    .clk(clk100m),
    .d(freq7[6]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [6]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b7  (
    .clk(clk100m),
    .d(freq7[7]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [7]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b8  (
    .clk(clk100m),
    .d(freq7[8]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [8]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg1_b9  (
    .clk(clk100m),
    .d(freq7[9]),
    .en(\PWM7/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/FreCntr [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM7/reg2_b0  (
    .clk(clk100m),
    .d(\PWM7/n23 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[0]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b1  (
    .clk(clk100m),
    .d(\PWM7/n23 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[1]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b10  (
    .clk(clk100m),
    .d(\PWM7/n23 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[10]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b11  (
    .clk(clk100m),
    .d(\PWM7/n23 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[11]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b12  (
    .clk(clk100m),
    .d(\PWM7/n23 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[12]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b13  (
    .clk(clk100m),
    .d(\PWM7/n23 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[13]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b14  (
    .clk(clk100m),
    .d(\PWM7/n23 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[14]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b15  (
    .clk(clk100m),
    .d(\PWM7/n23 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[15]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b16  (
    .clk(clk100m),
    .d(\PWM7/n23 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[16]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b17  (
    .clk(clk100m),
    .d(\PWM7/n23 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[17]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b18  (
    .clk(clk100m),
    .d(\PWM7/n23 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[18]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b19  (
    .clk(clk100m),
    .d(\PWM7/n23 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[19]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b2  (
    .clk(clk100m),
    .d(\PWM7/n23 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[2]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b20  (
    .clk(clk100m),
    .d(\PWM7/n23 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[20]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b21  (
    .clk(clk100m),
    .d(\PWM7/n23 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[21]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b22  (
    .clk(clk100m),
    .d(\PWM7/n23 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[22]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b23  (
    .clk(clk100m),
    .d(\PWM7/n23 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[23]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b24  (
    .clk(clk100m),
    .d(\PWM7/n23 [24]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[24]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b25  (
    .clk(clk100m),
    .d(\PWM7/n23 [25]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[25]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b26  (
    .clk(clk100m),
    .d(\PWM7/n23 [26]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[26]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b27  (
    .clk(clk100m),
    .d(\PWM7/n23 [27]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[27]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b28  (
    .clk(clk100m),
    .d(\PWM7/n23 [28]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[28]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b29  (
    .clk(clk100m),
    .d(\PWM7/n23 [29]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[29]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b3  (
    .clk(clk100m),
    .d(\PWM7/n23 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[3]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b30  (
    .clk(clk100m),
    .d(\PWM7/n23 [30]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[30]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b31  (
    .clk(clk100m),
    .d(\PWM7/n23 [31]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[31]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b4  (
    .clk(clk100m),
    .d(\PWM7/n23 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[4]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b5  (
    .clk(clk100m),
    .d(\PWM7/n23 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[5]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b6  (
    .clk(clk100m),
    .d(\PWM7/n23 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[6]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b7  (
    .clk(clk100m),
    .d(\PWM7/n23 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[7]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b8  (
    .clk(clk100m),
    .d(\PWM7/n23 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[8]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg2_b9  (
    .clk(clk100m),
    .d(\PWM7/n23 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/pnumr[9]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM7/reg3_b0  (
    .clk(clk100m),
    .d(\PWM7/n31 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[0]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b1  (
    .clk(clk100m),
    .d(\PWM7/n31 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[1]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b10  (
    .clk(clk100m),
    .d(\PWM7/n31 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[10]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b11  (
    .clk(clk100m),
    .d(\PWM7/n31 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[11]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b12  (
    .clk(clk100m),
    .d(\PWM7/n31 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[12]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b13  (
    .clk(clk100m),
    .d(\PWM7/n31 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[13]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b14  (
    .clk(clk100m),
    .d(\PWM7/n31 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[14]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b15  (
    .clk(clk100m),
    .d(\PWM7/n31 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[15]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b16  (
    .clk(clk100m),
    .d(\PWM7/n31 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[16]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b17  (
    .clk(clk100m),
    .d(\PWM7/n31 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[17]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b18  (
    .clk(clk100m),
    .d(\PWM7/n31 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[18]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b19  (
    .clk(clk100m),
    .d(\PWM7/n31 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[19]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b2  (
    .clk(clk100m),
    .d(\PWM7/n31 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[2]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b20  (
    .clk(clk100m),
    .d(\PWM7/n31 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[20]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b21  (
    .clk(clk100m),
    .d(\PWM7/n31 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[21]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b22  (
    .clk(clk100m),
    .d(\PWM7/n31 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[22]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b23  (
    .clk(clk100m),
    .d(\PWM7/n31 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[23]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b3  (
    .clk(clk100m),
    .d(\PWM7/n31 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[3]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b4  (
    .clk(clk100m),
    .d(\PWM7/n31 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[4]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b5  (
    .clk(clk100m),
    .d(\PWM7/n31 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[5]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b6  (
    .clk(clk100m),
    .d(\PWM7/n31 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[6]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b7  (
    .clk(clk100m),
    .d(\PWM7/n31 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[7]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b8  (
    .clk(clk100m),
    .d(\PWM7/n31 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[8]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM7/reg3_b9  (
    .clk(clk100m),
    .d(\PWM7/n31 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM7/RemaTxNum[9]_keep ));  // src/OnePWM.v(58)
  reg_ar_ss_w1 \PWM7/stopreq_reg  (
    .clk(clk100m),
    .d(\PWM7/n1 ),
    .en(1'b1),
    .reset(1'b0),
    .set(pwm_start_stop[7]),
    .q(\PWM7/stopreq_keep ));  // src/OnePWM.v(15)
  add_pu27_mu27_o27 \PWM7/sub0  (
    .i0(\PWM7/FreCnt ),
    .i1(27'b000000000000000000000000001),
    .o(\PWM7/n12 [26:0]));  // src/OnePWM.v(32)
  add_pu24_mu24_o24 \PWM7/sub1  (
    .i0(pnumcnt7),
    .i1(24'b000000000000000000000001),
    .o(\PWM7/n26 [23:0]));  // src/OnePWM.v(55)
  AL_MUX \PWM7/u10  (
    .i0(1'b0),
    .i1(\PWM7/n9 ),
    .sel(n18),
    .o(\PWM7/n10 ));  // src/OnePWM.v(26)
  or \PWM7/u11  (\PWM7/n11 , pwm_state_read[7], pwm_start_stop[23]);  // src/OnePWM.v(30)
  and \PWM7/u14_sel_is_1  (\PWM7/u14_sel_is_1_o , pwm_state_read[7], \PWM7/n17_neg );
  and \PWM7/u15  (\PWM7/n24 , \PWM7/n0 , pwm_state_read[7]);  // src/OnePWM.v(54)
  and \PWM7/u17_sel_is_1  (\PWM7/u17_sel_is_1_o , \PWM7/n24 , \PWM7/n25_neg );
  not \PWM7/u17_sel_is_1_o_inv  (\PWM7/u17_sel_is_1_o_neg , \PWM7/u17_sel_is_1_o );
  AL_MUX \PWM7/u18  (
    .i0(\PWM7/pnumr [31]),
    .i1(dir[7]),
    .sel(\PWM7/u18_sel_is_0_o ),
    .o(\PWM7/n32 ));
  and \PWM7/u18_sel_is_0  (\PWM7/u18_sel_is_0_o , \pwm_start_stop[23]_neg , \PWM7/u17_sel_is_1_o_neg );
  AL_MUX \PWM7/u2  (
    .i0(\PWM7/stopreq ),
    .i1(1'b0),
    .sel(\PWM7/n0 ),
    .o(\PWM7/n1 ));  // src/OnePWM.v(15)
  and \PWM7/u5  (\PWM7/n4 , \PWM7/stopreq , \PWM7/n0 );  // src/OnePWM.v(23)
  and \PWM7/u6  (\PWM7/n6 , \PWM7/n5 , \PWM7/n0 );  // src/OnePWM.v(25)
  AL_MUX \PWM7/u8  (
    .i0(1'b0),
    .i1(pwm_state_read[7]),
    .sel(\PWM7/u8_sel_is_0_o ),
    .o(\PWM7/n8 ));
  and \PWM7/u8_sel_is_0  (\PWM7/u8_sel_is_0_o , \PWM7/n4_neg , \PWM7/n6_neg );
  AL_MUX \PWM7/u9  (
    .i0(\PWM7/n8 ),
    .i1(1'b1),
    .sel(pwm_start_stop[23]),
    .o(\PWM7/n9 ));  // src/OnePWM.v(26)
  reg_ar_as_w1 \PWM8/State_reg  (
    .clk(clk100m),
    .d(\PWM8/n10 ),
    .en(1'b1),
    .reset(~rstn),
    .set(1'b0),
    .q(pwm_state_read[8]));  // src/OnePWM.v(26)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[0]  (
    .i(\PWM8/RemaTxNum[0]_keep ),
    .o(pnumcnt8[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[10]  (
    .i(\PWM8/RemaTxNum[10]_keep ),
    .o(pnumcnt8[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[11]  (
    .i(\PWM8/RemaTxNum[11]_keep ),
    .o(pnumcnt8[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[12]  (
    .i(\PWM8/RemaTxNum[12]_keep ),
    .o(pnumcnt8[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[13]  (
    .i(\PWM8/RemaTxNum[13]_keep ),
    .o(pnumcnt8[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[14]  (
    .i(\PWM8/RemaTxNum[14]_keep ),
    .o(pnumcnt8[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[15]  (
    .i(\PWM8/RemaTxNum[15]_keep ),
    .o(pnumcnt8[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[16]  (
    .i(\PWM8/RemaTxNum[16]_keep ),
    .o(pnumcnt8[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[17]  (
    .i(\PWM8/RemaTxNum[17]_keep ),
    .o(pnumcnt8[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[18]  (
    .i(\PWM8/RemaTxNum[18]_keep ),
    .o(pnumcnt8[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[19]  (
    .i(\PWM8/RemaTxNum[19]_keep ),
    .o(pnumcnt8[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[1]  (
    .i(\PWM8/RemaTxNum[1]_keep ),
    .o(pnumcnt8[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[20]  (
    .i(\PWM8/RemaTxNum[20]_keep ),
    .o(pnumcnt8[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[21]  (
    .i(\PWM8/RemaTxNum[21]_keep ),
    .o(pnumcnt8[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[22]  (
    .i(\PWM8/RemaTxNum[22]_keep ),
    .o(pnumcnt8[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[23]  (
    .i(\PWM8/RemaTxNum[23]_keep ),
    .o(pnumcnt8[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[2]  (
    .i(\PWM8/RemaTxNum[2]_keep ),
    .o(pnumcnt8[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[3]  (
    .i(\PWM8/RemaTxNum[3]_keep ),
    .o(pnumcnt8[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[4]  (
    .i(\PWM8/RemaTxNum[4]_keep ),
    .o(pnumcnt8[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[5]  (
    .i(\PWM8/RemaTxNum[5]_keep ),
    .o(pnumcnt8[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[6]  (
    .i(\PWM8/RemaTxNum[6]_keep ),
    .o(pnumcnt8[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[7]  (
    .i(\PWM8/RemaTxNum[7]_keep ),
    .o(pnumcnt8[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[8]  (
    .i(\PWM8/RemaTxNum[8]_keep ),
    .o(pnumcnt8[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_RemaTxNum[9]  (
    .i(\PWM8/RemaTxNum[9]_keep ),
    .o(pnumcnt8[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_dir  (
    .i(\PWM8/dir_keep ),
    .o(dir[8]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[0]  (
    .i(\PWM8/pnumr[0]_keep ),
    .o(\PWM8/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[10]  (
    .i(\PWM8/pnumr[10]_keep ),
    .o(\PWM8/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[11]  (
    .i(\PWM8/pnumr[11]_keep ),
    .o(\PWM8/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[12]  (
    .i(\PWM8/pnumr[12]_keep ),
    .o(\PWM8/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[13]  (
    .i(\PWM8/pnumr[13]_keep ),
    .o(\PWM8/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[14]  (
    .i(\PWM8/pnumr[14]_keep ),
    .o(\PWM8/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[15]  (
    .i(\PWM8/pnumr[15]_keep ),
    .o(\PWM8/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[16]  (
    .i(\PWM8/pnumr[16]_keep ),
    .o(\PWM8/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[17]  (
    .i(\PWM8/pnumr[17]_keep ),
    .o(\PWM8/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[18]  (
    .i(\PWM8/pnumr[18]_keep ),
    .o(\PWM8/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[19]  (
    .i(\PWM8/pnumr[19]_keep ),
    .o(\PWM8/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[1]  (
    .i(\PWM8/pnumr[1]_keep ),
    .o(\PWM8/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[20]  (
    .i(\PWM8/pnumr[20]_keep ),
    .o(\PWM8/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[21]  (
    .i(\PWM8/pnumr[21]_keep ),
    .o(\PWM8/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[22]  (
    .i(\PWM8/pnumr[22]_keep ),
    .o(\PWM8/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[23]  (
    .i(\PWM8/pnumr[23]_keep ),
    .o(\PWM8/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[24]  (
    .i(\PWM8/pnumr[24]_keep ),
    .o(\PWM8/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[25]  (
    .i(\PWM8/pnumr[25]_keep ),
    .o(\PWM8/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[26]  (
    .i(\PWM8/pnumr[26]_keep ),
    .o(\PWM8/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[27]  (
    .i(\PWM8/pnumr[27]_keep ),
    .o(\PWM8/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[28]  (
    .i(\PWM8/pnumr[28]_keep ),
    .o(\PWM8/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[29]  (
    .i(\PWM8/pnumr[29]_keep ),
    .o(\PWM8/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[2]  (
    .i(\PWM8/pnumr[2]_keep ),
    .o(\PWM8/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[30]  (
    .i(\PWM8/pnumr[30]_keep ),
    .o(\PWM8/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[31]  (
    .i(\PWM8/pnumr[31]_keep ),
    .o(\PWM8/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[3]  (
    .i(\PWM8/pnumr[3]_keep ),
    .o(\PWM8/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[4]  (
    .i(\PWM8/pnumr[4]_keep ),
    .o(\PWM8/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[5]  (
    .i(\PWM8/pnumr[5]_keep ),
    .o(\PWM8/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[6]  (
    .i(\PWM8/pnumr[6]_keep ),
    .o(\PWM8/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[7]  (
    .i(\PWM8/pnumr[7]_keep ),
    .o(\PWM8/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[8]  (
    .i(\PWM8/pnumr[8]_keep ),
    .o(\PWM8/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pnumr[9]  (
    .i(\PWM8/pnumr[9]_keep ),
    .o(\PWM8/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_pwm  (
    .i(\PWM8/pwm_keep ),
    .o(pwm[8]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM8/_bufkeep_stopreq  (
    .i(\PWM8/stopreq_keep ),
    .o(\PWM8/stopreq ));  // src/OnePWM.v(14)
  reg_ar_as_w1 \PWM8/dir_reg  (
    .clk(clk100m),
    .d(\PWM8/n32 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/dir_keep ));  // src/OnePWM.v(58)
  eq_w27 \PWM8/eq0  (
    .i0(\PWM8/FreCnt ),
    .i1(27'b000000000000000000000000000),
    .o(\PWM8/n0 ));  // src/OnePWM.v(15)
  eq_w24 \PWM8/eq1  (
    .i0(pnumcnt8),
    .i1(24'b000000000000000000000001),
    .o(\PWM8/n5 ));  // src/OnePWM.v(25)
  eq_w27 \PWM8/eq2  (
    .i0(\PWM8/FreCnt ),
    .i1({1'b0,\PWM8/FreCntr [26:1]}),
    .o(\PWM8/n17 ));  // src/OnePWM.v(41)
  eq_w27 \PWM8/eq3  (
    .i0(\PWM8/FreCnt ),
    .i1(\PWM8/FreCntr ),
    .o(\PWM8/n18 ));  // src/OnePWM.v(43)
  binary_mux_s1_w1 \PWM8/mux0_b0  (
    .i0(\PWM8/n12 [0]),
    .i1(freq8[0]),
    .sel(\PWM8/n0 ),
    .o(\PWM8/n13 [0]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM8/mux0_b1  (
    .i0(\PWM8/n12 [1]),
    .i1(freq8[1]),
    .sel(\PWM8/n0 ),
    .o(\PWM8/n13 [1]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM8/mux0_b10  (
    .i0(\PWM8/n12 [10]),
    .i1(freq8[10]),
    .sel(\PWM8/n0 ),
    .o(\PWM8/n13 [10]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM8/mux0_b11  (
    .i0(\PWM8/n12 [11]),
    .i1(freq8[11]),
    .sel(\PWM8/n0 ),
    .o(\PWM8/n13 [11]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM8/mux0_b12  (
    .i0(\PWM8/n12 [12]),
    .i1(freq8[12]),
    .sel(\PWM8/n0 ),
    .o(\PWM8/n13 [12]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM8/mux0_b13  (
    .i0(\PWM8/n12 [13]),
    .i1(freq8[13]),
    .sel(\PWM8/n0 ),
    .o(\PWM8/n13 [13]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM8/mux0_b14  (
    .i0(\PWM8/n12 [14]),
    .i1(freq8[14]),
    .sel(\PWM8/n0 ),
    .o(\PWM8/n13 [14]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM8/mux0_b15  (
    .i0(\PWM8/n12 [15]),
    .i1(freq8[15]),
    .sel(\PWM8/n0 ),
    .o(\PWM8/n13 [15]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM8/mux0_b16  (
    .i0(\PWM8/n12 [16]),
    .i1(freq8[16]),
    .sel(\PWM8/n0 ),
    .o(\PWM8/n13 [16]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM8/mux0_b17  (
    .i0(\PWM8/n12 [17]),
    .i1(freq8[17]),
    .sel(\PWM8/n0 ),
    .o(\PWM8/n13 [17]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM8/mux0_b18  (
    .i0(\PWM8/n12 [18]),
    .i1(freq8[18]),
    .sel(\PWM8/n0 ),
    .o(\PWM8/n13 [18]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM8/mux0_b19  (
    .i0(\PWM8/n12 [19]),
    .i1(freq8[19]),
    .sel(\PWM8/n0 ),
    .o(\PWM8/n13 [19]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM8/mux0_b2  (
    .i0(\PWM8/n12 [2]),
    .i1(freq8[2]),
    .sel(\PWM8/n0 ),
    .o(\PWM8/n13 [2]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM8/mux0_b20  (
    .i0(\PWM8/n12 [20]),
    .i1(freq8[20]),
    .sel(\PWM8/n0 ),
    .o(\PWM8/n13 [20]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM8/mux0_b21  (
    .i0(\PWM8/n12 [21]),
    .i1(freq8[21]),
    .sel(\PWM8/n0 ),
    .o(\PWM8/n13 [21]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM8/mux0_b22  (
    .i0(\PWM8/n12 [22]),
    .i1(freq8[22]),
    .sel(\PWM8/n0 ),
    .o(\PWM8/n13 [22]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM8/mux0_b23  (
    .i0(\PWM8/n12 [23]),
    .i1(freq8[23]),
    .sel(\PWM8/n0 ),
    .o(\PWM8/n13 [23]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM8/mux0_b24  (
    .i0(\PWM8/n12 [24]),
    .i1(freq8[24]),
    .sel(\PWM8/n0 ),
    .o(\PWM8/n13 [24]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM8/mux0_b25  (
    .i0(\PWM8/n12 [25]),
    .i1(freq8[25]),
    .sel(\PWM8/n0 ),
    .o(\PWM8/n13 [25]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM8/mux0_b26  (
    .i0(\PWM8/n12 [26]),
    .i1(freq8[26]),
    .sel(\PWM8/n0 ),
    .o(\PWM8/n13 [26]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM8/mux0_b3  (
    .i0(\PWM8/n12 [3]),
    .i1(freq8[3]),
    .sel(\PWM8/n0 ),
    .o(\PWM8/n13 [3]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM8/mux0_b4  (
    .i0(\PWM8/n12 [4]),
    .i1(freq8[4]),
    .sel(\PWM8/n0 ),
    .o(\PWM8/n13 [4]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM8/mux0_b5  (
    .i0(\PWM8/n12 [5]),
    .i1(freq8[5]),
    .sel(\PWM8/n0 ),
    .o(\PWM8/n13 [5]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM8/mux0_b6  (
    .i0(\PWM8/n12 [6]),
    .i1(freq8[6]),
    .sel(\PWM8/n0 ),
    .o(\PWM8/n13 [6]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM8/mux0_b7  (
    .i0(\PWM8/n12 [7]),
    .i1(freq8[7]),
    .sel(\PWM8/n0 ),
    .o(\PWM8/n13 [7]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM8/mux0_b8  (
    .i0(\PWM8/n12 [8]),
    .i1(freq8[8]),
    .sel(\PWM8/n0 ),
    .o(\PWM8/n13 [8]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM8/mux0_b9  (
    .i0(\PWM8/n12 [9]),
    .i1(freq8[9]),
    .sel(\PWM8/n0 ),
    .o(\PWM8/n13 [9]));  // src/OnePWM.v(32)
  and \PWM8/mux3_b0_sel_is_3  (\PWM8/mux3_b0_sel_is_3_o , \PWM8/n11 , \PWM8/n0 );
  binary_mux_s1_w1 \PWM8/mux4_b0  (
    .i0(\PWM8/pnumr [0]),
    .i1(1'b0),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n22 [0]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux4_b1  (
    .i0(\PWM8/pnumr [1]),
    .i1(1'b0),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n22 [1]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux4_b10  (
    .i0(\PWM8/pnumr [10]),
    .i1(1'b0),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n22 [10]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux4_b11  (
    .i0(\PWM8/pnumr [11]),
    .i1(1'b0),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n22 [11]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux4_b12  (
    .i0(\PWM8/pnumr [12]),
    .i1(1'b0),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n22 [12]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux4_b13  (
    .i0(\PWM8/pnumr [13]),
    .i1(1'b0),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n22 [13]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux4_b14  (
    .i0(\PWM8/pnumr [14]),
    .i1(1'b0),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n22 [14]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux4_b15  (
    .i0(\PWM8/pnumr [15]),
    .i1(1'b0),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n22 [15]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux4_b16  (
    .i0(\PWM8/pnumr [16]),
    .i1(1'b0),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n22 [16]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux4_b17  (
    .i0(\PWM8/pnumr [17]),
    .i1(1'b0),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n22 [17]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux4_b18  (
    .i0(\PWM8/pnumr [18]),
    .i1(1'b0),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n22 [18]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux4_b19  (
    .i0(\PWM8/pnumr [19]),
    .i1(1'b0),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n22 [19]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux4_b2  (
    .i0(\PWM8/pnumr [2]),
    .i1(1'b0),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n22 [2]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux4_b20  (
    .i0(\PWM8/pnumr [20]),
    .i1(1'b0),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n22 [20]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux4_b21  (
    .i0(\PWM8/pnumr [21]),
    .i1(1'b0),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n22 [21]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux4_b22  (
    .i0(\PWM8/pnumr [22]),
    .i1(1'b0),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n22 [22]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux4_b23  (
    .i0(\PWM8/pnumr [23]),
    .i1(1'b0),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n22 [23]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux4_b24  (
    .i0(\PWM8/pnumr [24]),
    .i1(1'b0),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n22 [24]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux4_b25  (
    .i0(\PWM8/pnumr [25]),
    .i1(1'b0),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n22 [25]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux4_b26  (
    .i0(\PWM8/pnumr [26]),
    .i1(1'b0),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n22 [26]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux4_b27  (
    .i0(\PWM8/pnumr [27]),
    .i1(1'b0),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n22 [27]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux4_b28  (
    .i0(\PWM8/pnumr [28]),
    .i1(1'b0),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n22 [28]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux4_b29  (
    .i0(\PWM8/pnumr [29]),
    .i1(1'b0),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n22 [29]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux4_b3  (
    .i0(\PWM8/pnumr [3]),
    .i1(1'b0),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n22 [3]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux4_b30  (
    .i0(\PWM8/pnumr [30]),
    .i1(1'b0),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n22 [30]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux4_b31  (
    .i0(\PWM8/pnumr [31]),
    .i1(1'b0),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n22 [31]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux4_b4  (
    .i0(\PWM8/pnumr [4]),
    .i1(1'b0),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n22 [4]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux4_b5  (
    .i0(\PWM8/pnumr [5]),
    .i1(1'b0),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n22 [5]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux4_b6  (
    .i0(\PWM8/pnumr [6]),
    .i1(1'b0),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n22 [6]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux4_b7  (
    .i0(\PWM8/pnumr [7]),
    .i1(1'b0),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n22 [7]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux4_b8  (
    .i0(\PWM8/pnumr [8]),
    .i1(1'b0),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n22 [8]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux4_b9  (
    .i0(\PWM8/pnumr [9]),
    .i1(1'b0),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n22 [9]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux5_b0  (
    .i0(\PWM8/n22 [0]),
    .i1(pnum8[0]),
    .sel(pnum8[32]),
    .o(\PWM8/n23 [0]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux5_b1  (
    .i0(\PWM8/n22 [1]),
    .i1(pnum8[1]),
    .sel(pnum8[32]),
    .o(\PWM8/n23 [1]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux5_b10  (
    .i0(\PWM8/n22 [10]),
    .i1(pnum8[10]),
    .sel(pnum8[32]),
    .o(\PWM8/n23 [10]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux5_b11  (
    .i0(\PWM8/n22 [11]),
    .i1(pnum8[11]),
    .sel(pnum8[32]),
    .o(\PWM8/n23 [11]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux5_b12  (
    .i0(\PWM8/n22 [12]),
    .i1(pnum8[12]),
    .sel(pnum8[32]),
    .o(\PWM8/n23 [12]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux5_b13  (
    .i0(\PWM8/n22 [13]),
    .i1(pnum8[13]),
    .sel(pnum8[32]),
    .o(\PWM8/n23 [13]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux5_b14  (
    .i0(\PWM8/n22 [14]),
    .i1(pnum8[14]),
    .sel(pnum8[32]),
    .o(\PWM8/n23 [14]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux5_b15  (
    .i0(\PWM8/n22 [15]),
    .i1(pnum8[15]),
    .sel(pnum8[32]),
    .o(\PWM8/n23 [15]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux5_b16  (
    .i0(\PWM8/n22 [16]),
    .i1(pnum8[16]),
    .sel(pnum8[32]),
    .o(\PWM8/n23 [16]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux5_b17  (
    .i0(\PWM8/n22 [17]),
    .i1(pnum8[17]),
    .sel(pnum8[32]),
    .o(\PWM8/n23 [17]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux5_b18  (
    .i0(\PWM8/n22 [18]),
    .i1(pnum8[18]),
    .sel(pnum8[32]),
    .o(\PWM8/n23 [18]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux5_b19  (
    .i0(\PWM8/n22 [19]),
    .i1(pnum8[19]),
    .sel(pnum8[32]),
    .o(\PWM8/n23 [19]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux5_b2  (
    .i0(\PWM8/n22 [2]),
    .i1(pnum8[2]),
    .sel(pnum8[32]),
    .o(\PWM8/n23 [2]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux5_b20  (
    .i0(\PWM8/n22 [20]),
    .i1(pnum8[20]),
    .sel(pnum8[32]),
    .o(\PWM8/n23 [20]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux5_b21  (
    .i0(\PWM8/n22 [21]),
    .i1(pnum8[21]),
    .sel(pnum8[32]),
    .o(\PWM8/n23 [21]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux5_b22  (
    .i0(\PWM8/n22 [22]),
    .i1(pnum8[22]),
    .sel(pnum8[32]),
    .o(\PWM8/n23 [22]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux5_b23  (
    .i0(\PWM8/n22 [23]),
    .i1(pnum8[23]),
    .sel(pnum8[32]),
    .o(\PWM8/n23 [23]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux5_b24  (
    .i0(\PWM8/n22 [24]),
    .i1(pnum8[24]),
    .sel(pnum8[32]),
    .o(\PWM8/n23 [24]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux5_b25  (
    .i0(\PWM8/n22 [25]),
    .i1(pnum8[25]),
    .sel(pnum8[32]),
    .o(\PWM8/n23 [25]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux5_b26  (
    .i0(\PWM8/n22 [26]),
    .i1(pnum8[26]),
    .sel(pnum8[32]),
    .o(\PWM8/n23 [26]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux5_b27  (
    .i0(\PWM8/n22 [27]),
    .i1(pnum8[27]),
    .sel(pnum8[32]),
    .o(\PWM8/n23 [27]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux5_b28  (
    .i0(\PWM8/n22 [28]),
    .i1(pnum8[28]),
    .sel(pnum8[32]),
    .o(\PWM8/n23 [28]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux5_b29  (
    .i0(\PWM8/n22 [29]),
    .i1(pnum8[29]),
    .sel(pnum8[32]),
    .o(\PWM8/n23 [29]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux5_b3  (
    .i0(\PWM8/n22 [3]),
    .i1(pnum8[3]),
    .sel(pnum8[32]),
    .o(\PWM8/n23 [3]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux5_b30  (
    .i0(\PWM8/n22 [30]),
    .i1(pnum8[30]),
    .sel(pnum8[32]),
    .o(\PWM8/n23 [30]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux5_b31  (
    .i0(\PWM8/n22 [31]),
    .i1(pnum8[31]),
    .sel(pnum8[32]),
    .o(\PWM8/n23 [31]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux5_b4  (
    .i0(\PWM8/n22 [4]),
    .i1(pnum8[4]),
    .sel(pnum8[32]),
    .o(\PWM8/n23 [4]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux5_b5  (
    .i0(\PWM8/n22 [5]),
    .i1(pnum8[5]),
    .sel(pnum8[32]),
    .o(\PWM8/n23 [5]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux5_b6  (
    .i0(\PWM8/n22 [6]),
    .i1(pnum8[6]),
    .sel(pnum8[32]),
    .o(\PWM8/n23 [6]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux5_b7  (
    .i0(\PWM8/n22 [7]),
    .i1(pnum8[7]),
    .sel(pnum8[32]),
    .o(\PWM8/n23 [7]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux5_b8  (
    .i0(\PWM8/n22 [8]),
    .i1(pnum8[8]),
    .sel(pnum8[32]),
    .o(\PWM8/n23 [8]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux5_b9  (
    .i0(\PWM8/n22 [9]),
    .i1(pnum8[9]),
    .sel(pnum8[32]),
    .o(\PWM8/n23 [9]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM8/mux6_b0  (
    .i0(\PWM8/pnumr [0]),
    .i1(\PWM8/n26 [0]),
    .sel(\PWM8/n25 ),
    .o(\PWM8/n27 [0]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM8/mux6_b1  (
    .i0(\PWM8/pnumr [1]),
    .i1(\PWM8/n26 [1]),
    .sel(\PWM8/n25 ),
    .o(\PWM8/n27 [1]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM8/mux6_b10  (
    .i0(\PWM8/pnumr [10]),
    .i1(\PWM8/n26 [10]),
    .sel(\PWM8/n25 ),
    .o(\PWM8/n27 [10]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM8/mux6_b11  (
    .i0(\PWM8/pnumr [11]),
    .i1(\PWM8/n26 [11]),
    .sel(\PWM8/n25 ),
    .o(\PWM8/n27 [11]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM8/mux6_b12  (
    .i0(\PWM8/pnumr [12]),
    .i1(\PWM8/n26 [12]),
    .sel(\PWM8/n25 ),
    .o(\PWM8/n27 [12]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM8/mux6_b13  (
    .i0(\PWM8/pnumr [13]),
    .i1(\PWM8/n26 [13]),
    .sel(\PWM8/n25 ),
    .o(\PWM8/n27 [13]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM8/mux6_b14  (
    .i0(\PWM8/pnumr [14]),
    .i1(\PWM8/n26 [14]),
    .sel(\PWM8/n25 ),
    .o(\PWM8/n27 [14]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM8/mux6_b15  (
    .i0(\PWM8/pnumr [15]),
    .i1(\PWM8/n26 [15]),
    .sel(\PWM8/n25 ),
    .o(\PWM8/n27 [15]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM8/mux6_b16  (
    .i0(\PWM8/pnumr [16]),
    .i1(\PWM8/n26 [16]),
    .sel(\PWM8/n25 ),
    .o(\PWM8/n27 [16]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM8/mux6_b17  (
    .i0(\PWM8/pnumr [17]),
    .i1(\PWM8/n26 [17]),
    .sel(\PWM8/n25 ),
    .o(\PWM8/n27 [17]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM8/mux6_b18  (
    .i0(\PWM8/pnumr [18]),
    .i1(\PWM8/n26 [18]),
    .sel(\PWM8/n25 ),
    .o(\PWM8/n27 [18]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM8/mux6_b19  (
    .i0(\PWM8/pnumr [19]),
    .i1(\PWM8/n26 [19]),
    .sel(\PWM8/n25 ),
    .o(\PWM8/n27 [19]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM8/mux6_b2  (
    .i0(\PWM8/pnumr [2]),
    .i1(\PWM8/n26 [2]),
    .sel(\PWM8/n25 ),
    .o(\PWM8/n27 [2]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM8/mux6_b20  (
    .i0(\PWM8/pnumr [20]),
    .i1(\PWM8/n26 [20]),
    .sel(\PWM8/n25 ),
    .o(\PWM8/n27 [20]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM8/mux6_b21  (
    .i0(\PWM8/pnumr [21]),
    .i1(\PWM8/n26 [21]),
    .sel(\PWM8/n25 ),
    .o(\PWM8/n27 [21]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM8/mux6_b22  (
    .i0(\PWM8/pnumr [22]),
    .i1(\PWM8/n26 [22]),
    .sel(\PWM8/n25 ),
    .o(\PWM8/n27 [22]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM8/mux6_b23  (
    .i0(\PWM8/pnumr [23]),
    .i1(\PWM8/n26 [23]),
    .sel(\PWM8/n25 ),
    .o(\PWM8/n27 [23]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM8/mux6_b3  (
    .i0(\PWM8/pnumr [3]),
    .i1(\PWM8/n26 [3]),
    .sel(\PWM8/n25 ),
    .o(\PWM8/n27 [3]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM8/mux6_b4  (
    .i0(\PWM8/pnumr [4]),
    .i1(\PWM8/n26 [4]),
    .sel(\PWM8/n25 ),
    .o(\PWM8/n27 [4]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM8/mux6_b5  (
    .i0(\PWM8/pnumr [5]),
    .i1(\PWM8/n26 [5]),
    .sel(\PWM8/n25 ),
    .o(\PWM8/n27 [5]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM8/mux6_b6  (
    .i0(\PWM8/pnumr [6]),
    .i1(\PWM8/n26 [6]),
    .sel(\PWM8/n25 ),
    .o(\PWM8/n27 [6]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM8/mux6_b7  (
    .i0(\PWM8/pnumr [7]),
    .i1(\PWM8/n26 [7]),
    .sel(\PWM8/n25 ),
    .o(\PWM8/n27 [7]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM8/mux6_b8  (
    .i0(\PWM8/pnumr [8]),
    .i1(\PWM8/n26 [8]),
    .sel(\PWM8/n25 ),
    .o(\PWM8/n27 [8]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM8/mux6_b9  (
    .i0(\PWM8/pnumr [9]),
    .i1(\PWM8/n26 [9]),
    .sel(\PWM8/n25 ),
    .o(\PWM8/n27 [9]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM8/mux7_b0  (
    .i0(pnumcnt8[0]),
    .i1(\PWM8/n27 [0]),
    .sel(\PWM8/n24 ),
    .o(\PWM8/n29 [0]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux7_b1  (
    .i0(pnumcnt8[1]),
    .i1(\PWM8/n27 [1]),
    .sel(\PWM8/n24 ),
    .o(\PWM8/n29 [1]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux7_b10  (
    .i0(pnumcnt8[10]),
    .i1(\PWM8/n27 [10]),
    .sel(\PWM8/n24 ),
    .o(\PWM8/n29 [10]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux7_b11  (
    .i0(pnumcnt8[11]),
    .i1(\PWM8/n27 [11]),
    .sel(\PWM8/n24 ),
    .o(\PWM8/n29 [11]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux7_b12  (
    .i0(pnumcnt8[12]),
    .i1(\PWM8/n27 [12]),
    .sel(\PWM8/n24 ),
    .o(\PWM8/n29 [12]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux7_b13  (
    .i0(pnumcnt8[13]),
    .i1(\PWM8/n27 [13]),
    .sel(\PWM8/n24 ),
    .o(\PWM8/n29 [13]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux7_b14  (
    .i0(pnumcnt8[14]),
    .i1(\PWM8/n27 [14]),
    .sel(\PWM8/n24 ),
    .o(\PWM8/n29 [14]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux7_b15  (
    .i0(pnumcnt8[15]),
    .i1(\PWM8/n27 [15]),
    .sel(\PWM8/n24 ),
    .o(\PWM8/n29 [15]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux7_b16  (
    .i0(pnumcnt8[16]),
    .i1(\PWM8/n27 [16]),
    .sel(\PWM8/n24 ),
    .o(\PWM8/n29 [16]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux7_b17  (
    .i0(pnumcnt8[17]),
    .i1(\PWM8/n27 [17]),
    .sel(\PWM8/n24 ),
    .o(\PWM8/n29 [17]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux7_b18  (
    .i0(pnumcnt8[18]),
    .i1(\PWM8/n27 [18]),
    .sel(\PWM8/n24 ),
    .o(\PWM8/n29 [18]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux7_b19  (
    .i0(pnumcnt8[19]),
    .i1(\PWM8/n27 [19]),
    .sel(\PWM8/n24 ),
    .o(\PWM8/n29 [19]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux7_b2  (
    .i0(pnumcnt8[2]),
    .i1(\PWM8/n27 [2]),
    .sel(\PWM8/n24 ),
    .o(\PWM8/n29 [2]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux7_b20  (
    .i0(pnumcnt8[20]),
    .i1(\PWM8/n27 [20]),
    .sel(\PWM8/n24 ),
    .o(\PWM8/n29 [20]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux7_b21  (
    .i0(pnumcnt8[21]),
    .i1(\PWM8/n27 [21]),
    .sel(\PWM8/n24 ),
    .o(\PWM8/n29 [21]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux7_b22  (
    .i0(pnumcnt8[22]),
    .i1(\PWM8/n27 [22]),
    .sel(\PWM8/n24 ),
    .o(\PWM8/n29 [22]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux7_b23  (
    .i0(pnumcnt8[23]),
    .i1(\PWM8/n27 [23]),
    .sel(\PWM8/n24 ),
    .o(\PWM8/n29 [23]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux7_b3  (
    .i0(pnumcnt8[3]),
    .i1(\PWM8/n27 [3]),
    .sel(\PWM8/n24 ),
    .o(\PWM8/n29 [3]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux7_b4  (
    .i0(pnumcnt8[4]),
    .i1(\PWM8/n27 [4]),
    .sel(\PWM8/n24 ),
    .o(\PWM8/n29 [4]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux7_b5  (
    .i0(pnumcnt8[5]),
    .i1(\PWM8/n27 [5]),
    .sel(\PWM8/n24 ),
    .o(\PWM8/n29 [5]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux7_b6  (
    .i0(pnumcnt8[6]),
    .i1(\PWM8/n27 [6]),
    .sel(\PWM8/n24 ),
    .o(\PWM8/n29 [6]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux7_b7  (
    .i0(pnumcnt8[7]),
    .i1(\PWM8/n27 [7]),
    .sel(\PWM8/n24 ),
    .o(\PWM8/n29 [7]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux7_b8  (
    .i0(pnumcnt8[8]),
    .i1(\PWM8/n27 [8]),
    .sel(\PWM8/n24 ),
    .o(\PWM8/n29 [8]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux7_b9  (
    .i0(pnumcnt8[9]),
    .i1(\PWM8/n27 [9]),
    .sel(\PWM8/n24 ),
    .o(\PWM8/n29 [9]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux8_b0  (
    .i0(\PWM8/n29 [0]),
    .i1(\PWM8/pnumr [0]),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n31 [0]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux8_b1  (
    .i0(\PWM8/n29 [1]),
    .i1(\PWM8/pnumr [1]),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n31 [1]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux8_b10  (
    .i0(\PWM8/n29 [10]),
    .i1(\PWM8/pnumr [10]),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n31 [10]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux8_b11  (
    .i0(\PWM8/n29 [11]),
    .i1(\PWM8/pnumr [11]),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n31 [11]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux8_b12  (
    .i0(\PWM8/n29 [12]),
    .i1(\PWM8/pnumr [12]),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n31 [12]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux8_b13  (
    .i0(\PWM8/n29 [13]),
    .i1(\PWM8/pnumr [13]),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n31 [13]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux8_b14  (
    .i0(\PWM8/n29 [14]),
    .i1(\PWM8/pnumr [14]),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n31 [14]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux8_b15  (
    .i0(\PWM8/n29 [15]),
    .i1(\PWM8/pnumr [15]),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n31 [15]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux8_b16  (
    .i0(\PWM8/n29 [16]),
    .i1(\PWM8/pnumr [16]),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n31 [16]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux8_b17  (
    .i0(\PWM8/n29 [17]),
    .i1(\PWM8/pnumr [17]),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n31 [17]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux8_b18  (
    .i0(\PWM8/n29 [18]),
    .i1(\PWM8/pnumr [18]),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n31 [18]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux8_b19  (
    .i0(\PWM8/n29 [19]),
    .i1(\PWM8/pnumr [19]),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n31 [19]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux8_b2  (
    .i0(\PWM8/n29 [2]),
    .i1(\PWM8/pnumr [2]),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n31 [2]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux8_b20  (
    .i0(\PWM8/n29 [20]),
    .i1(\PWM8/pnumr [20]),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n31 [20]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux8_b21  (
    .i0(\PWM8/n29 [21]),
    .i1(\PWM8/pnumr [21]),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n31 [21]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux8_b22  (
    .i0(\PWM8/n29 [22]),
    .i1(\PWM8/pnumr [22]),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n31 [22]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux8_b23  (
    .i0(\PWM8/n29 [23]),
    .i1(\PWM8/pnumr [23]),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n31 [23]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux8_b3  (
    .i0(\PWM8/n29 [3]),
    .i1(\PWM8/pnumr [3]),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n31 [3]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux8_b4  (
    .i0(\PWM8/n29 [4]),
    .i1(\PWM8/pnumr [4]),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n31 [4]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux8_b5  (
    .i0(\PWM8/n29 [5]),
    .i1(\PWM8/pnumr [5]),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n31 [5]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux8_b6  (
    .i0(\PWM8/n29 [6]),
    .i1(\PWM8/pnumr [6]),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n31 [6]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux8_b7  (
    .i0(\PWM8/n29 [7]),
    .i1(\PWM8/pnumr [7]),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n31 [7]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux8_b8  (
    .i0(\PWM8/n29 [8]),
    .i1(\PWM8/pnumr [8]),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n31 [8]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM8/mux8_b9  (
    .i0(\PWM8/n29 [9]),
    .i1(\PWM8/pnumr [9]),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n31 [9]));  // src/OnePWM.v(57)
  not \PWM8/n17_inv  (\PWM8/n17_neg , \PWM8/n17 );
  not \PWM8/n25_inv  (\PWM8/n25_neg , \PWM8/n25 );
  not \PWM8/n4_inv  (\PWM8/n4_neg , \PWM8/n4 );
  not \PWM8/n6_inv  (\PWM8/n6_neg , \PWM8/n6 );
  ne_w24 \PWM8/neq0  (
    .i0(pnumcnt8),
    .i1(24'b000000000000000000000000),
    .o(\PWM8/n25 ));  // src/OnePWM.v(55)
  reg_sr_ss_w1 \PWM8/pwm_reg  (
    .clk(clk100m),
    .d(pwm[8]),
    .en(1'b1),
    .reset(~\PWM8/u14_sel_is_1_o ),
    .set(\PWM8/n18 ),
    .q(\PWM8/pwm_keep ));  // src/OnePWM.v(45)
  reg_sr_as_w1 \PWM8/reg0_b0  (
    .clk(clk100m),
    .d(\PWM8/n13 [0]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [0]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b1  (
    .clk(clk100m),
    .d(\PWM8/n13 [1]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [1]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b10  (
    .clk(clk100m),
    .d(\PWM8/n13 [10]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [10]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b11  (
    .clk(clk100m),
    .d(\PWM8/n13 [11]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [11]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b12  (
    .clk(clk100m),
    .d(\PWM8/n13 [12]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [12]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b13  (
    .clk(clk100m),
    .d(\PWM8/n13 [13]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [13]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b14  (
    .clk(clk100m),
    .d(\PWM8/n13 [14]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [14]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b15  (
    .clk(clk100m),
    .d(\PWM8/n13 [15]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [15]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b16  (
    .clk(clk100m),
    .d(\PWM8/n13 [16]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [16]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b17  (
    .clk(clk100m),
    .d(\PWM8/n13 [17]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [17]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b18  (
    .clk(clk100m),
    .d(\PWM8/n13 [18]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [18]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b19  (
    .clk(clk100m),
    .d(\PWM8/n13 [19]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [19]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b2  (
    .clk(clk100m),
    .d(\PWM8/n13 [2]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [2]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b20  (
    .clk(clk100m),
    .d(\PWM8/n13 [20]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [20]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b21  (
    .clk(clk100m),
    .d(\PWM8/n13 [21]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [21]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b22  (
    .clk(clk100m),
    .d(\PWM8/n13 [22]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [22]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b23  (
    .clk(clk100m),
    .d(\PWM8/n13 [23]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [23]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b24  (
    .clk(clk100m),
    .d(\PWM8/n13 [24]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [24]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b25  (
    .clk(clk100m),
    .d(\PWM8/n13 [25]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [25]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b26  (
    .clk(clk100m),
    .d(\PWM8/n13 [26]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [26]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b3  (
    .clk(clk100m),
    .d(\PWM8/n13 [3]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [3]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b4  (
    .clk(clk100m),
    .d(\PWM8/n13 [4]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [4]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b5  (
    .clk(clk100m),
    .d(\PWM8/n13 [5]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [5]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b6  (
    .clk(clk100m),
    .d(\PWM8/n13 [6]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [6]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b7  (
    .clk(clk100m),
    .d(\PWM8/n13 [7]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [7]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b8  (
    .clk(clk100m),
    .d(\PWM8/n13 [8]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [8]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM8/reg0_b9  (
    .clk(clk100m),
    .d(\PWM8/n13 [9]),
    .en(1'b1),
    .reset(~\PWM8/n11 ),
    .set(1'b0),
    .q(\PWM8/FreCnt [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b0  (
    .clk(clk100m),
    .d(freq8[0]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [0]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b1  (
    .clk(clk100m),
    .d(freq8[1]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [1]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b10  (
    .clk(clk100m),
    .d(freq8[10]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [10]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b11  (
    .clk(clk100m),
    .d(freq8[11]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [11]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b12  (
    .clk(clk100m),
    .d(freq8[12]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [12]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b13  (
    .clk(clk100m),
    .d(freq8[13]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [13]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b14  (
    .clk(clk100m),
    .d(freq8[14]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [14]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b15  (
    .clk(clk100m),
    .d(freq8[15]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [15]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b16  (
    .clk(clk100m),
    .d(freq8[16]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [16]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b17  (
    .clk(clk100m),
    .d(freq8[17]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [17]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b18  (
    .clk(clk100m),
    .d(freq8[18]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [18]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b19  (
    .clk(clk100m),
    .d(freq8[19]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [19]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b2  (
    .clk(clk100m),
    .d(freq8[2]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [2]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b20  (
    .clk(clk100m),
    .d(freq8[20]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [20]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b21  (
    .clk(clk100m),
    .d(freq8[21]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [21]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b22  (
    .clk(clk100m),
    .d(freq8[22]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [22]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b23  (
    .clk(clk100m),
    .d(freq8[23]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [23]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b24  (
    .clk(clk100m),
    .d(freq8[24]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [24]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b25  (
    .clk(clk100m),
    .d(freq8[25]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [25]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b26  (
    .clk(clk100m),
    .d(freq8[26]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [26]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b3  (
    .clk(clk100m),
    .d(freq8[3]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [3]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b4  (
    .clk(clk100m),
    .d(freq8[4]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [4]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b5  (
    .clk(clk100m),
    .d(freq8[5]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [5]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b6  (
    .clk(clk100m),
    .d(freq8[6]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [6]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b7  (
    .clk(clk100m),
    .d(freq8[7]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [7]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b8  (
    .clk(clk100m),
    .d(freq8[8]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [8]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg1_b9  (
    .clk(clk100m),
    .d(freq8[9]),
    .en(\PWM8/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/FreCntr [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM8/reg2_b0  (
    .clk(clk100m),
    .d(\PWM8/n23 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[0]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b1  (
    .clk(clk100m),
    .d(\PWM8/n23 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[1]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b10  (
    .clk(clk100m),
    .d(\PWM8/n23 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[10]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b11  (
    .clk(clk100m),
    .d(\PWM8/n23 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[11]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b12  (
    .clk(clk100m),
    .d(\PWM8/n23 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[12]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b13  (
    .clk(clk100m),
    .d(\PWM8/n23 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[13]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b14  (
    .clk(clk100m),
    .d(\PWM8/n23 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[14]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b15  (
    .clk(clk100m),
    .d(\PWM8/n23 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[15]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b16  (
    .clk(clk100m),
    .d(\PWM8/n23 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[16]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b17  (
    .clk(clk100m),
    .d(\PWM8/n23 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[17]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b18  (
    .clk(clk100m),
    .d(\PWM8/n23 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[18]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b19  (
    .clk(clk100m),
    .d(\PWM8/n23 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[19]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b2  (
    .clk(clk100m),
    .d(\PWM8/n23 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[2]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b20  (
    .clk(clk100m),
    .d(\PWM8/n23 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[20]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b21  (
    .clk(clk100m),
    .d(\PWM8/n23 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[21]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b22  (
    .clk(clk100m),
    .d(\PWM8/n23 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[22]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b23  (
    .clk(clk100m),
    .d(\PWM8/n23 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[23]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b24  (
    .clk(clk100m),
    .d(\PWM8/n23 [24]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[24]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b25  (
    .clk(clk100m),
    .d(\PWM8/n23 [25]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[25]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b26  (
    .clk(clk100m),
    .d(\PWM8/n23 [26]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[26]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b27  (
    .clk(clk100m),
    .d(\PWM8/n23 [27]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[27]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b28  (
    .clk(clk100m),
    .d(\PWM8/n23 [28]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[28]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b29  (
    .clk(clk100m),
    .d(\PWM8/n23 [29]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[29]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b3  (
    .clk(clk100m),
    .d(\PWM8/n23 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[3]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b30  (
    .clk(clk100m),
    .d(\PWM8/n23 [30]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[30]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b31  (
    .clk(clk100m),
    .d(\PWM8/n23 [31]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[31]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b4  (
    .clk(clk100m),
    .d(\PWM8/n23 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[4]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b5  (
    .clk(clk100m),
    .d(\PWM8/n23 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[5]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b6  (
    .clk(clk100m),
    .d(\PWM8/n23 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[6]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b7  (
    .clk(clk100m),
    .d(\PWM8/n23 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[7]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b8  (
    .clk(clk100m),
    .d(\PWM8/n23 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[8]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg2_b9  (
    .clk(clk100m),
    .d(\PWM8/n23 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/pnumr[9]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM8/reg3_b0  (
    .clk(clk100m),
    .d(\PWM8/n31 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[0]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b1  (
    .clk(clk100m),
    .d(\PWM8/n31 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[1]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b10  (
    .clk(clk100m),
    .d(\PWM8/n31 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[10]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b11  (
    .clk(clk100m),
    .d(\PWM8/n31 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[11]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b12  (
    .clk(clk100m),
    .d(\PWM8/n31 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[12]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b13  (
    .clk(clk100m),
    .d(\PWM8/n31 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[13]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b14  (
    .clk(clk100m),
    .d(\PWM8/n31 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[14]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b15  (
    .clk(clk100m),
    .d(\PWM8/n31 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[15]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b16  (
    .clk(clk100m),
    .d(\PWM8/n31 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[16]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b17  (
    .clk(clk100m),
    .d(\PWM8/n31 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[17]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b18  (
    .clk(clk100m),
    .d(\PWM8/n31 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[18]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b19  (
    .clk(clk100m),
    .d(\PWM8/n31 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[19]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b2  (
    .clk(clk100m),
    .d(\PWM8/n31 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[2]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b20  (
    .clk(clk100m),
    .d(\PWM8/n31 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[20]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b21  (
    .clk(clk100m),
    .d(\PWM8/n31 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[21]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b22  (
    .clk(clk100m),
    .d(\PWM8/n31 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[22]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b23  (
    .clk(clk100m),
    .d(\PWM8/n31 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[23]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b3  (
    .clk(clk100m),
    .d(\PWM8/n31 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[3]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b4  (
    .clk(clk100m),
    .d(\PWM8/n31 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[4]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b5  (
    .clk(clk100m),
    .d(\PWM8/n31 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[5]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b6  (
    .clk(clk100m),
    .d(\PWM8/n31 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[6]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b7  (
    .clk(clk100m),
    .d(\PWM8/n31 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[7]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b8  (
    .clk(clk100m),
    .d(\PWM8/n31 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[8]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM8/reg3_b9  (
    .clk(clk100m),
    .d(\PWM8/n31 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM8/RemaTxNum[9]_keep ));  // src/OnePWM.v(58)
  reg_ar_ss_w1 \PWM8/stopreq_reg  (
    .clk(clk100m),
    .d(\PWM8/n1 ),
    .en(1'b1),
    .reset(1'b0),
    .set(pwm_start_stop[8]),
    .q(\PWM8/stopreq_keep ));  // src/OnePWM.v(15)
  add_pu27_mu27_o27 \PWM8/sub0  (
    .i0(\PWM8/FreCnt ),
    .i1(27'b000000000000000000000000001),
    .o(\PWM8/n12 [26:0]));  // src/OnePWM.v(32)
  add_pu24_mu24_o24 \PWM8/sub1  (
    .i0(pnumcnt8),
    .i1(24'b000000000000000000000001),
    .o(\PWM8/n26 [23:0]));  // src/OnePWM.v(55)
  AL_MUX \PWM8/u10  (
    .i0(1'b0),
    .i1(\PWM8/n9 ),
    .sel(n19),
    .o(\PWM8/n10 ));  // src/OnePWM.v(26)
  or \PWM8/u11  (\PWM8/n11 , pwm_state_read[8], pwm_start_stop[24]);  // src/OnePWM.v(30)
  and \PWM8/u14_sel_is_1  (\PWM8/u14_sel_is_1_o , pwm_state_read[8], \PWM8/n17_neg );
  and \PWM8/u15  (\PWM8/n24 , \PWM8/n0 , pwm_state_read[8]);  // src/OnePWM.v(54)
  and \PWM8/u17_sel_is_1  (\PWM8/u17_sel_is_1_o , \PWM8/n24 , \PWM8/n25_neg );
  not \PWM8/u17_sel_is_1_o_inv  (\PWM8/u17_sel_is_1_o_neg , \PWM8/u17_sel_is_1_o );
  AL_MUX \PWM8/u18  (
    .i0(\PWM8/pnumr [31]),
    .i1(dir[8]),
    .sel(\PWM8/u18_sel_is_0_o ),
    .o(\PWM8/n32 ));
  and \PWM8/u18_sel_is_0  (\PWM8/u18_sel_is_0_o , \pwm_start_stop[24]_neg , \PWM8/u17_sel_is_1_o_neg );
  AL_MUX \PWM8/u2  (
    .i0(\PWM8/stopreq ),
    .i1(1'b0),
    .sel(\PWM8/n0 ),
    .o(\PWM8/n1 ));  // src/OnePWM.v(15)
  and \PWM8/u5  (\PWM8/n4 , \PWM8/stopreq , \PWM8/n0 );  // src/OnePWM.v(23)
  and \PWM8/u6  (\PWM8/n6 , \PWM8/n5 , \PWM8/n0 );  // src/OnePWM.v(25)
  AL_MUX \PWM8/u8  (
    .i0(1'b0),
    .i1(pwm_state_read[8]),
    .sel(\PWM8/u8_sel_is_0_o ),
    .o(\PWM8/n8 ));
  and \PWM8/u8_sel_is_0  (\PWM8/u8_sel_is_0_o , \PWM8/n4_neg , \PWM8/n6_neg );
  AL_MUX \PWM8/u9  (
    .i0(\PWM8/n8 ),
    .i1(1'b1),
    .sel(pwm_start_stop[24]),
    .o(\PWM8/n9 ));  // src/OnePWM.v(26)
  reg_ar_as_w1 \PWM9/State_reg  (
    .clk(clk100m),
    .d(\PWM9/n10 ),
    .en(1'b1),
    .reset(~rstn),
    .set(1'b0),
    .q(pwm_state_read[9]));  // src/OnePWM.v(26)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[0]  (
    .i(\PWM9/RemaTxNum[0]_keep ),
    .o(pnumcnt9[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[10]  (
    .i(\PWM9/RemaTxNum[10]_keep ),
    .o(pnumcnt9[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[11]  (
    .i(\PWM9/RemaTxNum[11]_keep ),
    .o(pnumcnt9[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[12]  (
    .i(\PWM9/RemaTxNum[12]_keep ),
    .o(pnumcnt9[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[13]  (
    .i(\PWM9/RemaTxNum[13]_keep ),
    .o(pnumcnt9[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[14]  (
    .i(\PWM9/RemaTxNum[14]_keep ),
    .o(pnumcnt9[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[15]  (
    .i(\PWM9/RemaTxNum[15]_keep ),
    .o(pnumcnt9[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[16]  (
    .i(\PWM9/RemaTxNum[16]_keep ),
    .o(pnumcnt9[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[17]  (
    .i(\PWM9/RemaTxNum[17]_keep ),
    .o(pnumcnt9[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[18]  (
    .i(\PWM9/RemaTxNum[18]_keep ),
    .o(pnumcnt9[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[19]  (
    .i(\PWM9/RemaTxNum[19]_keep ),
    .o(pnumcnt9[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[1]  (
    .i(\PWM9/RemaTxNum[1]_keep ),
    .o(pnumcnt9[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[20]  (
    .i(\PWM9/RemaTxNum[20]_keep ),
    .o(pnumcnt9[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[21]  (
    .i(\PWM9/RemaTxNum[21]_keep ),
    .o(pnumcnt9[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[22]  (
    .i(\PWM9/RemaTxNum[22]_keep ),
    .o(pnumcnt9[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[23]  (
    .i(\PWM9/RemaTxNum[23]_keep ),
    .o(pnumcnt9[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[2]  (
    .i(\PWM9/RemaTxNum[2]_keep ),
    .o(pnumcnt9[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[3]  (
    .i(\PWM9/RemaTxNum[3]_keep ),
    .o(pnumcnt9[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[4]  (
    .i(\PWM9/RemaTxNum[4]_keep ),
    .o(pnumcnt9[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[5]  (
    .i(\PWM9/RemaTxNum[5]_keep ),
    .o(pnumcnt9[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[6]  (
    .i(\PWM9/RemaTxNum[6]_keep ),
    .o(pnumcnt9[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[7]  (
    .i(\PWM9/RemaTxNum[7]_keep ),
    .o(pnumcnt9[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[8]  (
    .i(\PWM9/RemaTxNum[8]_keep ),
    .o(pnumcnt9[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_RemaTxNum[9]  (
    .i(\PWM9/RemaTxNum[9]_keep ),
    .o(pnumcnt9[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_dir  (
    .i(\PWM9/dir_keep ),
    .o(dir[9]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[0]  (
    .i(\PWM9/pnumr[0]_keep ),
    .o(\PWM9/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[10]  (
    .i(\PWM9/pnumr[10]_keep ),
    .o(\PWM9/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[11]  (
    .i(\PWM9/pnumr[11]_keep ),
    .o(\PWM9/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[12]  (
    .i(\PWM9/pnumr[12]_keep ),
    .o(\PWM9/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[13]  (
    .i(\PWM9/pnumr[13]_keep ),
    .o(\PWM9/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[14]  (
    .i(\PWM9/pnumr[14]_keep ),
    .o(\PWM9/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[15]  (
    .i(\PWM9/pnumr[15]_keep ),
    .o(\PWM9/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[16]  (
    .i(\PWM9/pnumr[16]_keep ),
    .o(\PWM9/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[17]  (
    .i(\PWM9/pnumr[17]_keep ),
    .o(\PWM9/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[18]  (
    .i(\PWM9/pnumr[18]_keep ),
    .o(\PWM9/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[19]  (
    .i(\PWM9/pnumr[19]_keep ),
    .o(\PWM9/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[1]  (
    .i(\PWM9/pnumr[1]_keep ),
    .o(\PWM9/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[20]  (
    .i(\PWM9/pnumr[20]_keep ),
    .o(\PWM9/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[21]  (
    .i(\PWM9/pnumr[21]_keep ),
    .o(\PWM9/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[22]  (
    .i(\PWM9/pnumr[22]_keep ),
    .o(\PWM9/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[23]  (
    .i(\PWM9/pnumr[23]_keep ),
    .o(\PWM9/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[24]  (
    .i(\PWM9/pnumr[24]_keep ),
    .o(\PWM9/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[25]  (
    .i(\PWM9/pnumr[25]_keep ),
    .o(\PWM9/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[26]  (
    .i(\PWM9/pnumr[26]_keep ),
    .o(\PWM9/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[27]  (
    .i(\PWM9/pnumr[27]_keep ),
    .o(\PWM9/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[28]  (
    .i(\PWM9/pnumr[28]_keep ),
    .o(\PWM9/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[29]  (
    .i(\PWM9/pnumr[29]_keep ),
    .o(\PWM9/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[2]  (
    .i(\PWM9/pnumr[2]_keep ),
    .o(\PWM9/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[30]  (
    .i(\PWM9/pnumr[30]_keep ),
    .o(\PWM9/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[31]  (
    .i(\PWM9/pnumr[31]_keep ),
    .o(\PWM9/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[3]  (
    .i(\PWM9/pnumr[3]_keep ),
    .o(\PWM9/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[4]  (
    .i(\PWM9/pnumr[4]_keep ),
    .o(\PWM9/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[5]  (
    .i(\PWM9/pnumr[5]_keep ),
    .o(\PWM9/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[6]  (
    .i(\PWM9/pnumr[6]_keep ),
    .o(\PWM9/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[7]  (
    .i(\PWM9/pnumr[7]_keep ),
    .o(\PWM9/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[8]  (
    .i(\PWM9/pnumr[8]_keep ),
    .o(\PWM9/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pnumr[9]  (
    .i(\PWM9/pnumr[9]_keep ),
    .o(\PWM9/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_pwm  (
    .i(\PWM9/pwm_keep ),
    .o(pwm[9]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWM9/_bufkeep_stopreq  (
    .i(\PWM9/stopreq_keep ),
    .o(\PWM9/stopreq ));  // src/OnePWM.v(14)
  reg_ar_as_w1 \PWM9/dir_reg  (
    .clk(clk100m),
    .d(\PWM9/n32 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/dir_keep ));  // src/OnePWM.v(58)
  eq_w27 \PWM9/eq0  (
    .i0(\PWM9/FreCnt ),
    .i1(27'b000000000000000000000000000),
    .o(\PWM9/n0 ));  // src/OnePWM.v(15)
  eq_w24 \PWM9/eq1  (
    .i0(pnumcnt9),
    .i1(24'b000000000000000000000001),
    .o(\PWM9/n5 ));  // src/OnePWM.v(25)
  eq_w27 \PWM9/eq2  (
    .i0(\PWM9/FreCnt ),
    .i1({1'b0,\PWM9/FreCntr [26:1]}),
    .o(\PWM9/n17 ));  // src/OnePWM.v(41)
  eq_w27 \PWM9/eq3  (
    .i0(\PWM9/FreCnt ),
    .i1(\PWM9/FreCntr ),
    .o(\PWM9/n18 ));  // src/OnePWM.v(43)
  binary_mux_s1_w1 \PWM9/mux0_b0  (
    .i0(\PWM9/n12 [0]),
    .i1(freq9[0]),
    .sel(\PWM9/n0 ),
    .o(\PWM9/n13 [0]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM9/mux0_b1  (
    .i0(\PWM9/n12 [1]),
    .i1(freq9[1]),
    .sel(\PWM9/n0 ),
    .o(\PWM9/n13 [1]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM9/mux0_b10  (
    .i0(\PWM9/n12 [10]),
    .i1(freq9[10]),
    .sel(\PWM9/n0 ),
    .o(\PWM9/n13 [10]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM9/mux0_b11  (
    .i0(\PWM9/n12 [11]),
    .i1(freq9[11]),
    .sel(\PWM9/n0 ),
    .o(\PWM9/n13 [11]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM9/mux0_b12  (
    .i0(\PWM9/n12 [12]),
    .i1(freq9[12]),
    .sel(\PWM9/n0 ),
    .o(\PWM9/n13 [12]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM9/mux0_b13  (
    .i0(\PWM9/n12 [13]),
    .i1(freq9[13]),
    .sel(\PWM9/n0 ),
    .o(\PWM9/n13 [13]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM9/mux0_b14  (
    .i0(\PWM9/n12 [14]),
    .i1(freq9[14]),
    .sel(\PWM9/n0 ),
    .o(\PWM9/n13 [14]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM9/mux0_b15  (
    .i0(\PWM9/n12 [15]),
    .i1(freq9[15]),
    .sel(\PWM9/n0 ),
    .o(\PWM9/n13 [15]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM9/mux0_b16  (
    .i0(\PWM9/n12 [16]),
    .i1(freq9[16]),
    .sel(\PWM9/n0 ),
    .o(\PWM9/n13 [16]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM9/mux0_b17  (
    .i0(\PWM9/n12 [17]),
    .i1(freq9[17]),
    .sel(\PWM9/n0 ),
    .o(\PWM9/n13 [17]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM9/mux0_b18  (
    .i0(\PWM9/n12 [18]),
    .i1(freq9[18]),
    .sel(\PWM9/n0 ),
    .o(\PWM9/n13 [18]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM9/mux0_b19  (
    .i0(\PWM9/n12 [19]),
    .i1(freq9[19]),
    .sel(\PWM9/n0 ),
    .o(\PWM9/n13 [19]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM9/mux0_b2  (
    .i0(\PWM9/n12 [2]),
    .i1(freq9[2]),
    .sel(\PWM9/n0 ),
    .o(\PWM9/n13 [2]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM9/mux0_b20  (
    .i0(\PWM9/n12 [20]),
    .i1(freq9[20]),
    .sel(\PWM9/n0 ),
    .o(\PWM9/n13 [20]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM9/mux0_b21  (
    .i0(\PWM9/n12 [21]),
    .i1(freq9[21]),
    .sel(\PWM9/n0 ),
    .o(\PWM9/n13 [21]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM9/mux0_b22  (
    .i0(\PWM9/n12 [22]),
    .i1(freq9[22]),
    .sel(\PWM9/n0 ),
    .o(\PWM9/n13 [22]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM9/mux0_b23  (
    .i0(\PWM9/n12 [23]),
    .i1(freq9[23]),
    .sel(\PWM9/n0 ),
    .o(\PWM9/n13 [23]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM9/mux0_b24  (
    .i0(\PWM9/n12 [24]),
    .i1(freq9[24]),
    .sel(\PWM9/n0 ),
    .o(\PWM9/n13 [24]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM9/mux0_b25  (
    .i0(\PWM9/n12 [25]),
    .i1(freq9[25]),
    .sel(\PWM9/n0 ),
    .o(\PWM9/n13 [25]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM9/mux0_b26  (
    .i0(\PWM9/n12 [26]),
    .i1(freq9[26]),
    .sel(\PWM9/n0 ),
    .o(\PWM9/n13 [26]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM9/mux0_b3  (
    .i0(\PWM9/n12 [3]),
    .i1(freq9[3]),
    .sel(\PWM9/n0 ),
    .o(\PWM9/n13 [3]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM9/mux0_b4  (
    .i0(\PWM9/n12 [4]),
    .i1(freq9[4]),
    .sel(\PWM9/n0 ),
    .o(\PWM9/n13 [4]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM9/mux0_b5  (
    .i0(\PWM9/n12 [5]),
    .i1(freq9[5]),
    .sel(\PWM9/n0 ),
    .o(\PWM9/n13 [5]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM9/mux0_b6  (
    .i0(\PWM9/n12 [6]),
    .i1(freq9[6]),
    .sel(\PWM9/n0 ),
    .o(\PWM9/n13 [6]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM9/mux0_b7  (
    .i0(\PWM9/n12 [7]),
    .i1(freq9[7]),
    .sel(\PWM9/n0 ),
    .o(\PWM9/n13 [7]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM9/mux0_b8  (
    .i0(\PWM9/n12 [8]),
    .i1(freq9[8]),
    .sel(\PWM9/n0 ),
    .o(\PWM9/n13 [8]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWM9/mux0_b9  (
    .i0(\PWM9/n12 [9]),
    .i1(freq9[9]),
    .sel(\PWM9/n0 ),
    .o(\PWM9/n13 [9]));  // src/OnePWM.v(32)
  and \PWM9/mux3_b0_sel_is_3  (\PWM9/mux3_b0_sel_is_3_o , \PWM9/n11 , \PWM9/n0 );
  binary_mux_s1_w1 \PWM9/mux4_b0  (
    .i0(\PWM9/pnumr [0]),
    .i1(1'b0),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n22 [0]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux4_b1  (
    .i0(\PWM9/pnumr [1]),
    .i1(1'b0),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n22 [1]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux4_b10  (
    .i0(\PWM9/pnumr [10]),
    .i1(1'b0),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n22 [10]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux4_b11  (
    .i0(\PWM9/pnumr [11]),
    .i1(1'b0),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n22 [11]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux4_b12  (
    .i0(\PWM9/pnumr [12]),
    .i1(1'b0),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n22 [12]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux4_b13  (
    .i0(\PWM9/pnumr [13]),
    .i1(1'b0),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n22 [13]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux4_b14  (
    .i0(\PWM9/pnumr [14]),
    .i1(1'b0),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n22 [14]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux4_b15  (
    .i0(\PWM9/pnumr [15]),
    .i1(1'b0),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n22 [15]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux4_b16  (
    .i0(\PWM9/pnumr [16]),
    .i1(1'b0),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n22 [16]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux4_b17  (
    .i0(\PWM9/pnumr [17]),
    .i1(1'b0),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n22 [17]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux4_b18  (
    .i0(\PWM9/pnumr [18]),
    .i1(1'b0),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n22 [18]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux4_b19  (
    .i0(\PWM9/pnumr [19]),
    .i1(1'b0),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n22 [19]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux4_b2  (
    .i0(\PWM9/pnumr [2]),
    .i1(1'b0),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n22 [2]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux4_b20  (
    .i0(\PWM9/pnumr [20]),
    .i1(1'b0),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n22 [20]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux4_b21  (
    .i0(\PWM9/pnumr [21]),
    .i1(1'b0),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n22 [21]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux4_b22  (
    .i0(\PWM9/pnumr [22]),
    .i1(1'b0),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n22 [22]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux4_b23  (
    .i0(\PWM9/pnumr [23]),
    .i1(1'b0),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n22 [23]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux4_b24  (
    .i0(\PWM9/pnumr [24]),
    .i1(1'b0),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n22 [24]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux4_b25  (
    .i0(\PWM9/pnumr [25]),
    .i1(1'b0),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n22 [25]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux4_b26  (
    .i0(\PWM9/pnumr [26]),
    .i1(1'b0),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n22 [26]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux4_b27  (
    .i0(\PWM9/pnumr [27]),
    .i1(1'b0),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n22 [27]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux4_b28  (
    .i0(\PWM9/pnumr [28]),
    .i1(1'b0),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n22 [28]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux4_b29  (
    .i0(\PWM9/pnumr [29]),
    .i1(1'b0),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n22 [29]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux4_b3  (
    .i0(\PWM9/pnumr [3]),
    .i1(1'b0),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n22 [3]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux4_b30  (
    .i0(\PWM9/pnumr [30]),
    .i1(1'b0),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n22 [30]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux4_b31  (
    .i0(\PWM9/pnumr [31]),
    .i1(1'b0),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n22 [31]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux4_b4  (
    .i0(\PWM9/pnumr [4]),
    .i1(1'b0),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n22 [4]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux4_b5  (
    .i0(\PWM9/pnumr [5]),
    .i1(1'b0),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n22 [5]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux4_b6  (
    .i0(\PWM9/pnumr [6]),
    .i1(1'b0),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n22 [6]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux4_b7  (
    .i0(\PWM9/pnumr [7]),
    .i1(1'b0),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n22 [7]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux4_b8  (
    .i0(\PWM9/pnumr [8]),
    .i1(1'b0),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n22 [8]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux4_b9  (
    .i0(\PWM9/pnumr [9]),
    .i1(1'b0),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n22 [9]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux5_b0  (
    .i0(\PWM9/n22 [0]),
    .i1(pnum9[0]),
    .sel(pnum9[32]),
    .o(\PWM9/n23 [0]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux5_b1  (
    .i0(\PWM9/n22 [1]),
    .i1(pnum9[1]),
    .sel(pnum9[32]),
    .o(\PWM9/n23 [1]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux5_b10  (
    .i0(\PWM9/n22 [10]),
    .i1(pnum9[10]),
    .sel(pnum9[32]),
    .o(\PWM9/n23 [10]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux5_b11  (
    .i0(\PWM9/n22 [11]),
    .i1(pnum9[11]),
    .sel(pnum9[32]),
    .o(\PWM9/n23 [11]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux5_b12  (
    .i0(\PWM9/n22 [12]),
    .i1(pnum9[12]),
    .sel(pnum9[32]),
    .o(\PWM9/n23 [12]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux5_b13  (
    .i0(\PWM9/n22 [13]),
    .i1(pnum9[13]),
    .sel(pnum9[32]),
    .o(\PWM9/n23 [13]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux5_b14  (
    .i0(\PWM9/n22 [14]),
    .i1(pnum9[14]),
    .sel(pnum9[32]),
    .o(\PWM9/n23 [14]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux5_b15  (
    .i0(\PWM9/n22 [15]),
    .i1(pnum9[15]),
    .sel(pnum9[32]),
    .o(\PWM9/n23 [15]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux5_b16  (
    .i0(\PWM9/n22 [16]),
    .i1(pnum9[16]),
    .sel(pnum9[32]),
    .o(\PWM9/n23 [16]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux5_b17  (
    .i0(\PWM9/n22 [17]),
    .i1(pnum9[17]),
    .sel(pnum9[32]),
    .o(\PWM9/n23 [17]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux5_b18  (
    .i0(\PWM9/n22 [18]),
    .i1(pnum9[18]),
    .sel(pnum9[32]),
    .o(\PWM9/n23 [18]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux5_b19  (
    .i0(\PWM9/n22 [19]),
    .i1(pnum9[19]),
    .sel(pnum9[32]),
    .o(\PWM9/n23 [19]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux5_b2  (
    .i0(\PWM9/n22 [2]),
    .i1(pnum9[2]),
    .sel(pnum9[32]),
    .o(\PWM9/n23 [2]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux5_b20  (
    .i0(\PWM9/n22 [20]),
    .i1(pnum9[20]),
    .sel(pnum9[32]),
    .o(\PWM9/n23 [20]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux5_b21  (
    .i0(\PWM9/n22 [21]),
    .i1(pnum9[21]),
    .sel(pnum9[32]),
    .o(\PWM9/n23 [21]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux5_b22  (
    .i0(\PWM9/n22 [22]),
    .i1(pnum9[22]),
    .sel(pnum9[32]),
    .o(\PWM9/n23 [22]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux5_b23  (
    .i0(\PWM9/n22 [23]),
    .i1(pnum9[23]),
    .sel(pnum9[32]),
    .o(\PWM9/n23 [23]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux5_b24  (
    .i0(\PWM9/n22 [24]),
    .i1(pnum9[24]),
    .sel(pnum9[32]),
    .o(\PWM9/n23 [24]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux5_b25  (
    .i0(\PWM9/n22 [25]),
    .i1(pnum9[25]),
    .sel(pnum9[32]),
    .o(\PWM9/n23 [25]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux5_b26  (
    .i0(\PWM9/n22 [26]),
    .i1(pnum9[26]),
    .sel(pnum9[32]),
    .o(\PWM9/n23 [26]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux5_b27  (
    .i0(\PWM9/n22 [27]),
    .i1(pnum9[27]),
    .sel(pnum9[32]),
    .o(\PWM9/n23 [27]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux5_b28  (
    .i0(\PWM9/n22 [28]),
    .i1(pnum9[28]),
    .sel(pnum9[32]),
    .o(\PWM9/n23 [28]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux5_b29  (
    .i0(\PWM9/n22 [29]),
    .i1(pnum9[29]),
    .sel(pnum9[32]),
    .o(\PWM9/n23 [29]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux5_b3  (
    .i0(\PWM9/n22 [3]),
    .i1(pnum9[3]),
    .sel(pnum9[32]),
    .o(\PWM9/n23 [3]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux5_b30  (
    .i0(\PWM9/n22 [30]),
    .i1(pnum9[30]),
    .sel(pnum9[32]),
    .o(\PWM9/n23 [30]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux5_b31  (
    .i0(\PWM9/n22 [31]),
    .i1(pnum9[31]),
    .sel(pnum9[32]),
    .o(\PWM9/n23 [31]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux5_b4  (
    .i0(\PWM9/n22 [4]),
    .i1(pnum9[4]),
    .sel(pnum9[32]),
    .o(\PWM9/n23 [4]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux5_b5  (
    .i0(\PWM9/n22 [5]),
    .i1(pnum9[5]),
    .sel(pnum9[32]),
    .o(\PWM9/n23 [5]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux5_b6  (
    .i0(\PWM9/n22 [6]),
    .i1(pnum9[6]),
    .sel(pnum9[32]),
    .o(\PWM9/n23 [6]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux5_b7  (
    .i0(\PWM9/n22 [7]),
    .i1(pnum9[7]),
    .sel(pnum9[32]),
    .o(\PWM9/n23 [7]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux5_b8  (
    .i0(\PWM9/n22 [8]),
    .i1(pnum9[8]),
    .sel(pnum9[32]),
    .o(\PWM9/n23 [8]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux5_b9  (
    .i0(\PWM9/n22 [9]),
    .i1(pnum9[9]),
    .sel(pnum9[32]),
    .o(\PWM9/n23 [9]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWM9/mux6_b0  (
    .i0(\PWM9/pnumr [0]),
    .i1(\PWM9/n26 [0]),
    .sel(\PWM9/n25 ),
    .o(\PWM9/n27 [0]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM9/mux6_b1  (
    .i0(\PWM9/pnumr [1]),
    .i1(\PWM9/n26 [1]),
    .sel(\PWM9/n25 ),
    .o(\PWM9/n27 [1]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM9/mux6_b10  (
    .i0(\PWM9/pnumr [10]),
    .i1(\PWM9/n26 [10]),
    .sel(\PWM9/n25 ),
    .o(\PWM9/n27 [10]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM9/mux6_b11  (
    .i0(\PWM9/pnumr [11]),
    .i1(\PWM9/n26 [11]),
    .sel(\PWM9/n25 ),
    .o(\PWM9/n27 [11]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM9/mux6_b12  (
    .i0(\PWM9/pnumr [12]),
    .i1(\PWM9/n26 [12]),
    .sel(\PWM9/n25 ),
    .o(\PWM9/n27 [12]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM9/mux6_b13  (
    .i0(\PWM9/pnumr [13]),
    .i1(\PWM9/n26 [13]),
    .sel(\PWM9/n25 ),
    .o(\PWM9/n27 [13]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM9/mux6_b14  (
    .i0(\PWM9/pnumr [14]),
    .i1(\PWM9/n26 [14]),
    .sel(\PWM9/n25 ),
    .o(\PWM9/n27 [14]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM9/mux6_b15  (
    .i0(\PWM9/pnumr [15]),
    .i1(\PWM9/n26 [15]),
    .sel(\PWM9/n25 ),
    .o(\PWM9/n27 [15]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM9/mux6_b16  (
    .i0(\PWM9/pnumr [16]),
    .i1(\PWM9/n26 [16]),
    .sel(\PWM9/n25 ),
    .o(\PWM9/n27 [16]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM9/mux6_b17  (
    .i0(\PWM9/pnumr [17]),
    .i1(\PWM9/n26 [17]),
    .sel(\PWM9/n25 ),
    .o(\PWM9/n27 [17]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM9/mux6_b18  (
    .i0(\PWM9/pnumr [18]),
    .i1(\PWM9/n26 [18]),
    .sel(\PWM9/n25 ),
    .o(\PWM9/n27 [18]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM9/mux6_b19  (
    .i0(\PWM9/pnumr [19]),
    .i1(\PWM9/n26 [19]),
    .sel(\PWM9/n25 ),
    .o(\PWM9/n27 [19]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM9/mux6_b2  (
    .i0(\PWM9/pnumr [2]),
    .i1(\PWM9/n26 [2]),
    .sel(\PWM9/n25 ),
    .o(\PWM9/n27 [2]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM9/mux6_b20  (
    .i0(\PWM9/pnumr [20]),
    .i1(\PWM9/n26 [20]),
    .sel(\PWM9/n25 ),
    .o(\PWM9/n27 [20]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM9/mux6_b21  (
    .i0(\PWM9/pnumr [21]),
    .i1(\PWM9/n26 [21]),
    .sel(\PWM9/n25 ),
    .o(\PWM9/n27 [21]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM9/mux6_b22  (
    .i0(\PWM9/pnumr [22]),
    .i1(\PWM9/n26 [22]),
    .sel(\PWM9/n25 ),
    .o(\PWM9/n27 [22]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM9/mux6_b23  (
    .i0(\PWM9/pnumr [23]),
    .i1(\PWM9/n26 [23]),
    .sel(\PWM9/n25 ),
    .o(\PWM9/n27 [23]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM9/mux6_b3  (
    .i0(\PWM9/pnumr [3]),
    .i1(\PWM9/n26 [3]),
    .sel(\PWM9/n25 ),
    .o(\PWM9/n27 [3]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM9/mux6_b4  (
    .i0(\PWM9/pnumr [4]),
    .i1(\PWM9/n26 [4]),
    .sel(\PWM9/n25 ),
    .o(\PWM9/n27 [4]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM9/mux6_b5  (
    .i0(\PWM9/pnumr [5]),
    .i1(\PWM9/n26 [5]),
    .sel(\PWM9/n25 ),
    .o(\PWM9/n27 [5]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM9/mux6_b6  (
    .i0(\PWM9/pnumr [6]),
    .i1(\PWM9/n26 [6]),
    .sel(\PWM9/n25 ),
    .o(\PWM9/n27 [6]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM9/mux6_b7  (
    .i0(\PWM9/pnumr [7]),
    .i1(\PWM9/n26 [7]),
    .sel(\PWM9/n25 ),
    .o(\PWM9/n27 [7]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM9/mux6_b8  (
    .i0(\PWM9/pnumr [8]),
    .i1(\PWM9/n26 [8]),
    .sel(\PWM9/n25 ),
    .o(\PWM9/n27 [8]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM9/mux6_b9  (
    .i0(\PWM9/pnumr [9]),
    .i1(\PWM9/n26 [9]),
    .sel(\PWM9/n25 ),
    .o(\PWM9/n27 [9]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWM9/mux7_b0  (
    .i0(pnumcnt9[0]),
    .i1(\PWM9/n27 [0]),
    .sel(\PWM9/n24 ),
    .o(\PWM9/n29 [0]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux7_b1  (
    .i0(pnumcnt9[1]),
    .i1(\PWM9/n27 [1]),
    .sel(\PWM9/n24 ),
    .o(\PWM9/n29 [1]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux7_b10  (
    .i0(pnumcnt9[10]),
    .i1(\PWM9/n27 [10]),
    .sel(\PWM9/n24 ),
    .o(\PWM9/n29 [10]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux7_b11  (
    .i0(pnumcnt9[11]),
    .i1(\PWM9/n27 [11]),
    .sel(\PWM9/n24 ),
    .o(\PWM9/n29 [11]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux7_b12  (
    .i0(pnumcnt9[12]),
    .i1(\PWM9/n27 [12]),
    .sel(\PWM9/n24 ),
    .o(\PWM9/n29 [12]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux7_b13  (
    .i0(pnumcnt9[13]),
    .i1(\PWM9/n27 [13]),
    .sel(\PWM9/n24 ),
    .o(\PWM9/n29 [13]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux7_b14  (
    .i0(pnumcnt9[14]),
    .i1(\PWM9/n27 [14]),
    .sel(\PWM9/n24 ),
    .o(\PWM9/n29 [14]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux7_b15  (
    .i0(pnumcnt9[15]),
    .i1(\PWM9/n27 [15]),
    .sel(\PWM9/n24 ),
    .o(\PWM9/n29 [15]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux7_b16  (
    .i0(pnumcnt9[16]),
    .i1(\PWM9/n27 [16]),
    .sel(\PWM9/n24 ),
    .o(\PWM9/n29 [16]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux7_b17  (
    .i0(pnumcnt9[17]),
    .i1(\PWM9/n27 [17]),
    .sel(\PWM9/n24 ),
    .o(\PWM9/n29 [17]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux7_b18  (
    .i0(pnumcnt9[18]),
    .i1(\PWM9/n27 [18]),
    .sel(\PWM9/n24 ),
    .o(\PWM9/n29 [18]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux7_b19  (
    .i0(pnumcnt9[19]),
    .i1(\PWM9/n27 [19]),
    .sel(\PWM9/n24 ),
    .o(\PWM9/n29 [19]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux7_b2  (
    .i0(pnumcnt9[2]),
    .i1(\PWM9/n27 [2]),
    .sel(\PWM9/n24 ),
    .o(\PWM9/n29 [2]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux7_b20  (
    .i0(pnumcnt9[20]),
    .i1(\PWM9/n27 [20]),
    .sel(\PWM9/n24 ),
    .o(\PWM9/n29 [20]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux7_b21  (
    .i0(pnumcnt9[21]),
    .i1(\PWM9/n27 [21]),
    .sel(\PWM9/n24 ),
    .o(\PWM9/n29 [21]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux7_b22  (
    .i0(pnumcnt9[22]),
    .i1(\PWM9/n27 [22]),
    .sel(\PWM9/n24 ),
    .o(\PWM9/n29 [22]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux7_b23  (
    .i0(pnumcnt9[23]),
    .i1(\PWM9/n27 [23]),
    .sel(\PWM9/n24 ),
    .o(\PWM9/n29 [23]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux7_b3  (
    .i0(pnumcnt9[3]),
    .i1(\PWM9/n27 [3]),
    .sel(\PWM9/n24 ),
    .o(\PWM9/n29 [3]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux7_b4  (
    .i0(pnumcnt9[4]),
    .i1(\PWM9/n27 [4]),
    .sel(\PWM9/n24 ),
    .o(\PWM9/n29 [4]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux7_b5  (
    .i0(pnumcnt9[5]),
    .i1(\PWM9/n27 [5]),
    .sel(\PWM9/n24 ),
    .o(\PWM9/n29 [5]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux7_b6  (
    .i0(pnumcnt9[6]),
    .i1(\PWM9/n27 [6]),
    .sel(\PWM9/n24 ),
    .o(\PWM9/n29 [6]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux7_b7  (
    .i0(pnumcnt9[7]),
    .i1(\PWM9/n27 [7]),
    .sel(\PWM9/n24 ),
    .o(\PWM9/n29 [7]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux7_b8  (
    .i0(pnumcnt9[8]),
    .i1(\PWM9/n27 [8]),
    .sel(\PWM9/n24 ),
    .o(\PWM9/n29 [8]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux7_b9  (
    .i0(pnumcnt9[9]),
    .i1(\PWM9/n27 [9]),
    .sel(\PWM9/n24 ),
    .o(\PWM9/n29 [9]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux8_b0  (
    .i0(\PWM9/n29 [0]),
    .i1(\PWM9/pnumr [0]),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n31 [0]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux8_b1  (
    .i0(\PWM9/n29 [1]),
    .i1(\PWM9/pnumr [1]),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n31 [1]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux8_b10  (
    .i0(\PWM9/n29 [10]),
    .i1(\PWM9/pnumr [10]),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n31 [10]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux8_b11  (
    .i0(\PWM9/n29 [11]),
    .i1(\PWM9/pnumr [11]),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n31 [11]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux8_b12  (
    .i0(\PWM9/n29 [12]),
    .i1(\PWM9/pnumr [12]),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n31 [12]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux8_b13  (
    .i0(\PWM9/n29 [13]),
    .i1(\PWM9/pnumr [13]),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n31 [13]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux8_b14  (
    .i0(\PWM9/n29 [14]),
    .i1(\PWM9/pnumr [14]),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n31 [14]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux8_b15  (
    .i0(\PWM9/n29 [15]),
    .i1(\PWM9/pnumr [15]),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n31 [15]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux8_b16  (
    .i0(\PWM9/n29 [16]),
    .i1(\PWM9/pnumr [16]),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n31 [16]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux8_b17  (
    .i0(\PWM9/n29 [17]),
    .i1(\PWM9/pnumr [17]),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n31 [17]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux8_b18  (
    .i0(\PWM9/n29 [18]),
    .i1(\PWM9/pnumr [18]),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n31 [18]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux8_b19  (
    .i0(\PWM9/n29 [19]),
    .i1(\PWM9/pnumr [19]),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n31 [19]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux8_b2  (
    .i0(\PWM9/n29 [2]),
    .i1(\PWM9/pnumr [2]),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n31 [2]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux8_b20  (
    .i0(\PWM9/n29 [20]),
    .i1(\PWM9/pnumr [20]),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n31 [20]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux8_b21  (
    .i0(\PWM9/n29 [21]),
    .i1(\PWM9/pnumr [21]),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n31 [21]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux8_b22  (
    .i0(\PWM9/n29 [22]),
    .i1(\PWM9/pnumr [22]),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n31 [22]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux8_b23  (
    .i0(\PWM9/n29 [23]),
    .i1(\PWM9/pnumr [23]),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n31 [23]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux8_b3  (
    .i0(\PWM9/n29 [3]),
    .i1(\PWM9/pnumr [3]),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n31 [3]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux8_b4  (
    .i0(\PWM9/n29 [4]),
    .i1(\PWM9/pnumr [4]),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n31 [4]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux8_b5  (
    .i0(\PWM9/n29 [5]),
    .i1(\PWM9/pnumr [5]),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n31 [5]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux8_b6  (
    .i0(\PWM9/n29 [6]),
    .i1(\PWM9/pnumr [6]),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n31 [6]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux8_b7  (
    .i0(\PWM9/n29 [7]),
    .i1(\PWM9/pnumr [7]),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n31 [7]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux8_b8  (
    .i0(\PWM9/n29 [8]),
    .i1(\PWM9/pnumr [8]),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n31 [8]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWM9/mux8_b9  (
    .i0(\PWM9/n29 [9]),
    .i1(\PWM9/pnumr [9]),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n31 [9]));  // src/OnePWM.v(57)
  not \PWM9/n17_inv  (\PWM9/n17_neg , \PWM9/n17 );
  not \PWM9/n25_inv  (\PWM9/n25_neg , \PWM9/n25 );
  not \PWM9/n4_inv  (\PWM9/n4_neg , \PWM9/n4 );
  not \PWM9/n6_inv  (\PWM9/n6_neg , \PWM9/n6 );
  ne_w24 \PWM9/neq0  (
    .i0(pnumcnt9),
    .i1(24'b000000000000000000000000),
    .o(\PWM9/n25 ));  // src/OnePWM.v(55)
  reg_sr_ss_w1 \PWM9/pwm_reg  (
    .clk(clk100m),
    .d(pwm[9]),
    .en(1'b1),
    .reset(~\PWM9/u14_sel_is_1_o ),
    .set(\PWM9/n18 ),
    .q(\PWM9/pwm_keep ));  // src/OnePWM.v(45)
  reg_sr_as_w1 \PWM9/reg0_b0  (
    .clk(clk100m),
    .d(\PWM9/n13 [0]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [0]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b1  (
    .clk(clk100m),
    .d(\PWM9/n13 [1]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [1]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b10  (
    .clk(clk100m),
    .d(\PWM9/n13 [10]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [10]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b11  (
    .clk(clk100m),
    .d(\PWM9/n13 [11]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [11]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b12  (
    .clk(clk100m),
    .d(\PWM9/n13 [12]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [12]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b13  (
    .clk(clk100m),
    .d(\PWM9/n13 [13]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [13]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b14  (
    .clk(clk100m),
    .d(\PWM9/n13 [14]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [14]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b15  (
    .clk(clk100m),
    .d(\PWM9/n13 [15]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [15]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b16  (
    .clk(clk100m),
    .d(\PWM9/n13 [16]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [16]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b17  (
    .clk(clk100m),
    .d(\PWM9/n13 [17]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [17]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b18  (
    .clk(clk100m),
    .d(\PWM9/n13 [18]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [18]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b19  (
    .clk(clk100m),
    .d(\PWM9/n13 [19]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [19]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b2  (
    .clk(clk100m),
    .d(\PWM9/n13 [2]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [2]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b20  (
    .clk(clk100m),
    .d(\PWM9/n13 [20]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [20]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b21  (
    .clk(clk100m),
    .d(\PWM9/n13 [21]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [21]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b22  (
    .clk(clk100m),
    .d(\PWM9/n13 [22]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [22]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b23  (
    .clk(clk100m),
    .d(\PWM9/n13 [23]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [23]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b24  (
    .clk(clk100m),
    .d(\PWM9/n13 [24]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [24]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b25  (
    .clk(clk100m),
    .d(\PWM9/n13 [25]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [25]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b26  (
    .clk(clk100m),
    .d(\PWM9/n13 [26]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [26]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b3  (
    .clk(clk100m),
    .d(\PWM9/n13 [3]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [3]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b4  (
    .clk(clk100m),
    .d(\PWM9/n13 [4]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [4]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b5  (
    .clk(clk100m),
    .d(\PWM9/n13 [5]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [5]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b6  (
    .clk(clk100m),
    .d(\PWM9/n13 [6]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [6]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b7  (
    .clk(clk100m),
    .d(\PWM9/n13 [7]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [7]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b8  (
    .clk(clk100m),
    .d(\PWM9/n13 [8]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [8]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWM9/reg0_b9  (
    .clk(clk100m),
    .d(\PWM9/n13 [9]),
    .en(1'b1),
    .reset(~\PWM9/n11 ),
    .set(1'b0),
    .q(\PWM9/FreCnt [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b0  (
    .clk(clk100m),
    .d(freq9[0]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [0]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b1  (
    .clk(clk100m),
    .d(freq9[1]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [1]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b10  (
    .clk(clk100m),
    .d(freq9[10]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [10]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b11  (
    .clk(clk100m),
    .d(freq9[11]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [11]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b12  (
    .clk(clk100m),
    .d(freq9[12]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [12]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b13  (
    .clk(clk100m),
    .d(freq9[13]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [13]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b14  (
    .clk(clk100m),
    .d(freq9[14]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [14]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b15  (
    .clk(clk100m),
    .d(freq9[15]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [15]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b16  (
    .clk(clk100m),
    .d(freq9[16]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [16]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b17  (
    .clk(clk100m),
    .d(freq9[17]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [17]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b18  (
    .clk(clk100m),
    .d(freq9[18]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [18]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b19  (
    .clk(clk100m),
    .d(freq9[19]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [19]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b2  (
    .clk(clk100m),
    .d(freq9[2]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [2]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b20  (
    .clk(clk100m),
    .d(freq9[20]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [20]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b21  (
    .clk(clk100m),
    .d(freq9[21]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [21]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b22  (
    .clk(clk100m),
    .d(freq9[22]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [22]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b23  (
    .clk(clk100m),
    .d(freq9[23]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [23]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b24  (
    .clk(clk100m),
    .d(freq9[24]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [24]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b25  (
    .clk(clk100m),
    .d(freq9[25]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [25]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b26  (
    .clk(clk100m),
    .d(freq9[26]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [26]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b3  (
    .clk(clk100m),
    .d(freq9[3]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [3]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b4  (
    .clk(clk100m),
    .d(freq9[4]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [4]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b5  (
    .clk(clk100m),
    .d(freq9[5]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [5]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b6  (
    .clk(clk100m),
    .d(freq9[6]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [6]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b7  (
    .clk(clk100m),
    .d(freq9[7]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [7]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b8  (
    .clk(clk100m),
    .d(freq9[8]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [8]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg1_b9  (
    .clk(clk100m),
    .d(freq9[9]),
    .en(\PWM9/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/FreCntr [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWM9/reg2_b0  (
    .clk(clk100m),
    .d(\PWM9/n23 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[0]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b1  (
    .clk(clk100m),
    .d(\PWM9/n23 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[1]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b10  (
    .clk(clk100m),
    .d(\PWM9/n23 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[10]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b11  (
    .clk(clk100m),
    .d(\PWM9/n23 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[11]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b12  (
    .clk(clk100m),
    .d(\PWM9/n23 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[12]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b13  (
    .clk(clk100m),
    .d(\PWM9/n23 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[13]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b14  (
    .clk(clk100m),
    .d(\PWM9/n23 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[14]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b15  (
    .clk(clk100m),
    .d(\PWM9/n23 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[15]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b16  (
    .clk(clk100m),
    .d(\PWM9/n23 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[16]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b17  (
    .clk(clk100m),
    .d(\PWM9/n23 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[17]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b18  (
    .clk(clk100m),
    .d(\PWM9/n23 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[18]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b19  (
    .clk(clk100m),
    .d(\PWM9/n23 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[19]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b2  (
    .clk(clk100m),
    .d(\PWM9/n23 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[2]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b20  (
    .clk(clk100m),
    .d(\PWM9/n23 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[20]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b21  (
    .clk(clk100m),
    .d(\PWM9/n23 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[21]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b22  (
    .clk(clk100m),
    .d(\PWM9/n23 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[22]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b23  (
    .clk(clk100m),
    .d(\PWM9/n23 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[23]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b24  (
    .clk(clk100m),
    .d(\PWM9/n23 [24]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[24]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b25  (
    .clk(clk100m),
    .d(\PWM9/n23 [25]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[25]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b26  (
    .clk(clk100m),
    .d(\PWM9/n23 [26]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[26]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b27  (
    .clk(clk100m),
    .d(\PWM9/n23 [27]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[27]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b28  (
    .clk(clk100m),
    .d(\PWM9/n23 [28]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[28]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b29  (
    .clk(clk100m),
    .d(\PWM9/n23 [29]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[29]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b3  (
    .clk(clk100m),
    .d(\PWM9/n23 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[3]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b30  (
    .clk(clk100m),
    .d(\PWM9/n23 [30]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[30]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b31  (
    .clk(clk100m),
    .d(\PWM9/n23 [31]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[31]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b4  (
    .clk(clk100m),
    .d(\PWM9/n23 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[4]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b5  (
    .clk(clk100m),
    .d(\PWM9/n23 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[5]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b6  (
    .clk(clk100m),
    .d(\PWM9/n23 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[6]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b7  (
    .clk(clk100m),
    .d(\PWM9/n23 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[7]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b8  (
    .clk(clk100m),
    .d(\PWM9/n23 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[8]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg2_b9  (
    .clk(clk100m),
    .d(\PWM9/n23 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/pnumr[9]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWM9/reg3_b0  (
    .clk(clk100m),
    .d(\PWM9/n31 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[0]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b1  (
    .clk(clk100m),
    .d(\PWM9/n31 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[1]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b10  (
    .clk(clk100m),
    .d(\PWM9/n31 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[10]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b11  (
    .clk(clk100m),
    .d(\PWM9/n31 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[11]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b12  (
    .clk(clk100m),
    .d(\PWM9/n31 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[12]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b13  (
    .clk(clk100m),
    .d(\PWM9/n31 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[13]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b14  (
    .clk(clk100m),
    .d(\PWM9/n31 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[14]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b15  (
    .clk(clk100m),
    .d(\PWM9/n31 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[15]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b16  (
    .clk(clk100m),
    .d(\PWM9/n31 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[16]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b17  (
    .clk(clk100m),
    .d(\PWM9/n31 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[17]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b18  (
    .clk(clk100m),
    .d(\PWM9/n31 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[18]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b19  (
    .clk(clk100m),
    .d(\PWM9/n31 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[19]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b2  (
    .clk(clk100m),
    .d(\PWM9/n31 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[2]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b20  (
    .clk(clk100m),
    .d(\PWM9/n31 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[20]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b21  (
    .clk(clk100m),
    .d(\PWM9/n31 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[21]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b22  (
    .clk(clk100m),
    .d(\PWM9/n31 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[22]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b23  (
    .clk(clk100m),
    .d(\PWM9/n31 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[23]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b3  (
    .clk(clk100m),
    .d(\PWM9/n31 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[3]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b4  (
    .clk(clk100m),
    .d(\PWM9/n31 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[4]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b5  (
    .clk(clk100m),
    .d(\PWM9/n31 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[5]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b6  (
    .clk(clk100m),
    .d(\PWM9/n31 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[6]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b7  (
    .clk(clk100m),
    .d(\PWM9/n31 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[7]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b8  (
    .clk(clk100m),
    .d(\PWM9/n31 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[8]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWM9/reg3_b9  (
    .clk(clk100m),
    .d(\PWM9/n31 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWM9/RemaTxNum[9]_keep ));  // src/OnePWM.v(58)
  reg_ar_ss_w1 \PWM9/stopreq_reg  (
    .clk(clk100m),
    .d(\PWM9/n1 ),
    .en(1'b1),
    .reset(1'b0),
    .set(pwm_start_stop[9]),
    .q(\PWM9/stopreq_keep ));  // src/OnePWM.v(15)
  add_pu27_mu27_o27 \PWM9/sub0  (
    .i0(\PWM9/FreCnt ),
    .i1(27'b000000000000000000000000001),
    .o(\PWM9/n12 [26:0]));  // src/OnePWM.v(32)
  add_pu24_mu24_o24 \PWM9/sub1  (
    .i0(pnumcnt9),
    .i1(24'b000000000000000000000001),
    .o(\PWM9/n26 [23:0]));  // src/OnePWM.v(55)
  AL_MUX \PWM9/u10  (
    .i0(1'b0),
    .i1(\PWM9/n9 ),
    .sel(n20),
    .o(\PWM9/n10 ));  // src/OnePWM.v(26)
  or \PWM9/u11  (\PWM9/n11 , pwm_state_read[9], pwm_start_stop[25]);  // src/OnePWM.v(30)
  and \PWM9/u14_sel_is_1  (\PWM9/u14_sel_is_1_o , pwm_state_read[9], \PWM9/n17_neg );
  and \PWM9/u15  (\PWM9/n24 , \PWM9/n0 , pwm_state_read[9]);  // src/OnePWM.v(54)
  and \PWM9/u17_sel_is_1  (\PWM9/u17_sel_is_1_o , \PWM9/n24 , \PWM9/n25_neg );
  not \PWM9/u17_sel_is_1_o_inv  (\PWM9/u17_sel_is_1_o_neg , \PWM9/u17_sel_is_1_o );
  AL_MUX \PWM9/u18  (
    .i0(\PWM9/pnumr [31]),
    .i1(dir[9]),
    .sel(\PWM9/u18_sel_is_0_o ),
    .o(\PWM9/n32 ));
  and \PWM9/u18_sel_is_0  (\PWM9/u18_sel_is_0_o , \pwm_start_stop[25]_neg , \PWM9/u17_sel_is_1_o_neg );
  AL_MUX \PWM9/u2  (
    .i0(\PWM9/stopreq ),
    .i1(1'b0),
    .sel(\PWM9/n0 ),
    .o(\PWM9/n1 ));  // src/OnePWM.v(15)
  and \PWM9/u5  (\PWM9/n4 , \PWM9/stopreq , \PWM9/n0 );  // src/OnePWM.v(23)
  and \PWM9/u6  (\PWM9/n6 , \PWM9/n5 , \PWM9/n0 );  // src/OnePWM.v(25)
  AL_MUX \PWM9/u8  (
    .i0(1'b0),
    .i1(pwm_state_read[9]),
    .sel(\PWM9/u8_sel_is_0_o ),
    .o(\PWM9/n8 ));
  and \PWM9/u8_sel_is_0  (\PWM9/u8_sel_is_0_o , \PWM9/n4_neg , \PWM9/n6_neg );
  AL_MUX \PWM9/u9  (
    .i0(\PWM9/n8 ),
    .i1(1'b1),
    .sel(pwm_start_stop[25]),
    .o(\PWM9/n9 ));  // src/OnePWM.v(26)
  reg_ar_as_w1 \PWMA/State_reg  (
    .clk(clk100m),
    .d(\PWMA/n10 ),
    .en(1'b1),
    .reset(~rstn),
    .set(1'b0),
    .q(pwm_state_read[10]));  // src/OnePWM.v(26)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[0]  (
    .i(\PWMA/RemaTxNum[0]_keep ),
    .o(pnumcntA[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[10]  (
    .i(\PWMA/RemaTxNum[10]_keep ),
    .o(pnumcntA[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[11]  (
    .i(\PWMA/RemaTxNum[11]_keep ),
    .o(pnumcntA[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[12]  (
    .i(\PWMA/RemaTxNum[12]_keep ),
    .o(pnumcntA[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[13]  (
    .i(\PWMA/RemaTxNum[13]_keep ),
    .o(pnumcntA[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[14]  (
    .i(\PWMA/RemaTxNum[14]_keep ),
    .o(pnumcntA[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[15]  (
    .i(\PWMA/RemaTxNum[15]_keep ),
    .o(pnumcntA[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[16]  (
    .i(\PWMA/RemaTxNum[16]_keep ),
    .o(pnumcntA[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[17]  (
    .i(\PWMA/RemaTxNum[17]_keep ),
    .o(pnumcntA[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[18]  (
    .i(\PWMA/RemaTxNum[18]_keep ),
    .o(pnumcntA[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[19]  (
    .i(\PWMA/RemaTxNum[19]_keep ),
    .o(pnumcntA[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[1]  (
    .i(\PWMA/RemaTxNum[1]_keep ),
    .o(pnumcntA[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[20]  (
    .i(\PWMA/RemaTxNum[20]_keep ),
    .o(pnumcntA[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[21]  (
    .i(\PWMA/RemaTxNum[21]_keep ),
    .o(pnumcntA[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[22]  (
    .i(\PWMA/RemaTxNum[22]_keep ),
    .o(pnumcntA[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[23]  (
    .i(\PWMA/RemaTxNum[23]_keep ),
    .o(pnumcntA[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[2]  (
    .i(\PWMA/RemaTxNum[2]_keep ),
    .o(pnumcntA[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[3]  (
    .i(\PWMA/RemaTxNum[3]_keep ),
    .o(pnumcntA[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[4]  (
    .i(\PWMA/RemaTxNum[4]_keep ),
    .o(pnumcntA[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[5]  (
    .i(\PWMA/RemaTxNum[5]_keep ),
    .o(pnumcntA[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[6]  (
    .i(\PWMA/RemaTxNum[6]_keep ),
    .o(pnumcntA[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[7]  (
    .i(\PWMA/RemaTxNum[7]_keep ),
    .o(pnumcntA[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[8]  (
    .i(\PWMA/RemaTxNum[8]_keep ),
    .o(pnumcntA[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_RemaTxNum[9]  (
    .i(\PWMA/RemaTxNum[9]_keep ),
    .o(pnumcntA[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_dir  (
    .i(\PWMA/dir_keep ),
    .o(dir[10]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[0]  (
    .i(\PWMA/pnumr[0]_keep ),
    .o(\PWMA/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[10]  (
    .i(\PWMA/pnumr[10]_keep ),
    .o(\PWMA/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[11]  (
    .i(\PWMA/pnumr[11]_keep ),
    .o(\PWMA/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[12]  (
    .i(\PWMA/pnumr[12]_keep ),
    .o(\PWMA/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[13]  (
    .i(\PWMA/pnumr[13]_keep ),
    .o(\PWMA/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[14]  (
    .i(\PWMA/pnumr[14]_keep ),
    .o(\PWMA/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[15]  (
    .i(\PWMA/pnumr[15]_keep ),
    .o(\PWMA/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[16]  (
    .i(\PWMA/pnumr[16]_keep ),
    .o(\PWMA/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[17]  (
    .i(\PWMA/pnumr[17]_keep ),
    .o(\PWMA/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[18]  (
    .i(\PWMA/pnumr[18]_keep ),
    .o(\PWMA/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[19]  (
    .i(\PWMA/pnumr[19]_keep ),
    .o(\PWMA/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[1]  (
    .i(\PWMA/pnumr[1]_keep ),
    .o(\PWMA/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[20]  (
    .i(\PWMA/pnumr[20]_keep ),
    .o(\PWMA/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[21]  (
    .i(\PWMA/pnumr[21]_keep ),
    .o(\PWMA/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[22]  (
    .i(\PWMA/pnumr[22]_keep ),
    .o(\PWMA/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[23]  (
    .i(\PWMA/pnumr[23]_keep ),
    .o(\PWMA/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[24]  (
    .i(\PWMA/pnumr[24]_keep ),
    .o(\PWMA/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[25]  (
    .i(\PWMA/pnumr[25]_keep ),
    .o(\PWMA/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[26]  (
    .i(\PWMA/pnumr[26]_keep ),
    .o(\PWMA/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[27]  (
    .i(\PWMA/pnumr[27]_keep ),
    .o(\PWMA/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[28]  (
    .i(\PWMA/pnumr[28]_keep ),
    .o(\PWMA/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[29]  (
    .i(\PWMA/pnumr[29]_keep ),
    .o(\PWMA/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[2]  (
    .i(\PWMA/pnumr[2]_keep ),
    .o(\PWMA/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[30]  (
    .i(\PWMA/pnumr[30]_keep ),
    .o(\PWMA/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[31]  (
    .i(\PWMA/pnumr[31]_keep ),
    .o(\PWMA/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[3]  (
    .i(\PWMA/pnumr[3]_keep ),
    .o(\PWMA/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[4]  (
    .i(\PWMA/pnumr[4]_keep ),
    .o(\PWMA/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[5]  (
    .i(\PWMA/pnumr[5]_keep ),
    .o(\PWMA/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[6]  (
    .i(\PWMA/pnumr[6]_keep ),
    .o(\PWMA/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[7]  (
    .i(\PWMA/pnumr[7]_keep ),
    .o(\PWMA/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[8]  (
    .i(\PWMA/pnumr[8]_keep ),
    .o(\PWMA/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pnumr[9]  (
    .i(\PWMA/pnumr[9]_keep ),
    .o(\PWMA/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_pwm  (
    .i(\PWMA/pwm_keep ),
    .o(pwm[10]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMA/_bufkeep_stopreq  (
    .i(\PWMA/stopreq_keep ),
    .o(\PWMA/stopreq ));  // src/OnePWM.v(14)
  reg_ar_as_w1 \PWMA/dir_reg  (
    .clk(clk100m),
    .d(\PWMA/n32 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/dir_keep ));  // src/OnePWM.v(58)
  eq_w27 \PWMA/eq0  (
    .i0(\PWMA/FreCnt ),
    .i1(27'b000000000000000000000000000),
    .o(\PWMA/n0 ));  // src/OnePWM.v(15)
  eq_w24 \PWMA/eq1  (
    .i0(pnumcntA),
    .i1(24'b000000000000000000000001),
    .o(\PWMA/n5 ));  // src/OnePWM.v(25)
  eq_w27 \PWMA/eq2  (
    .i0(\PWMA/FreCnt ),
    .i1({1'b0,\PWMA/FreCntr [26:1]}),
    .o(\PWMA/n17 ));  // src/OnePWM.v(41)
  eq_w27 \PWMA/eq3  (
    .i0(\PWMA/FreCnt ),
    .i1(\PWMA/FreCntr ),
    .o(\PWMA/n18 ));  // src/OnePWM.v(43)
  binary_mux_s1_w1 \PWMA/mux0_b0  (
    .i0(\PWMA/n12 [0]),
    .i1(freqA[0]),
    .sel(\PWMA/n0 ),
    .o(\PWMA/n13 [0]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMA/mux0_b1  (
    .i0(\PWMA/n12 [1]),
    .i1(freqA[1]),
    .sel(\PWMA/n0 ),
    .o(\PWMA/n13 [1]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMA/mux0_b10  (
    .i0(\PWMA/n12 [10]),
    .i1(freqA[10]),
    .sel(\PWMA/n0 ),
    .o(\PWMA/n13 [10]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMA/mux0_b11  (
    .i0(\PWMA/n12 [11]),
    .i1(freqA[11]),
    .sel(\PWMA/n0 ),
    .o(\PWMA/n13 [11]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMA/mux0_b12  (
    .i0(\PWMA/n12 [12]),
    .i1(freqA[12]),
    .sel(\PWMA/n0 ),
    .o(\PWMA/n13 [12]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMA/mux0_b13  (
    .i0(\PWMA/n12 [13]),
    .i1(freqA[13]),
    .sel(\PWMA/n0 ),
    .o(\PWMA/n13 [13]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMA/mux0_b14  (
    .i0(\PWMA/n12 [14]),
    .i1(freqA[14]),
    .sel(\PWMA/n0 ),
    .o(\PWMA/n13 [14]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMA/mux0_b15  (
    .i0(\PWMA/n12 [15]),
    .i1(freqA[15]),
    .sel(\PWMA/n0 ),
    .o(\PWMA/n13 [15]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMA/mux0_b16  (
    .i0(\PWMA/n12 [16]),
    .i1(freqA[16]),
    .sel(\PWMA/n0 ),
    .o(\PWMA/n13 [16]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMA/mux0_b17  (
    .i0(\PWMA/n12 [17]),
    .i1(freqA[17]),
    .sel(\PWMA/n0 ),
    .o(\PWMA/n13 [17]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMA/mux0_b18  (
    .i0(\PWMA/n12 [18]),
    .i1(freqA[18]),
    .sel(\PWMA/n0 ),
    .o(\PWMA/n13 [18]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMA/mux0_b19  (
    .i0(\PWMA/n12 [19]),
    .i1(freqA[19]),
    .sel(\PWMA/n0 ),
    .o(\PWMA/n13 [19]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMA/mux0_b2  (
    .i0(\PWMA/n12 [2]),
    .i1(freqA[2]),
    .sel(\PWMA/n0 ),
    .o(\PWMA/n13 [2]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMA/mux0_b20  (
    .i0(\PWMA/n12 [20]),
    .i1(freqA[20]),
    .sel(\PWMA/n0 ),
    .o(\PWMA/n13 [20]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMA/mux0_b21  (
    .i0(\PWMA/n12 [21]),
    .i1(freqA[21]),
    .sel(\PWMA/n0 ),
    .o(\PWMA/n13 [21]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMA/mux0_b22  (
    .i0(\PWMA/n12 [22]),
    .i1(freqA[22]),
    .sel(\PWMA/n0 ),
    .o(\PWMA/n13 [22]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMA/mux0_b23  (
    .i0(\PWMA/n12 [23]),
    .i1(freqA[23]),
    .sel(\PWMA/n0 ),
    .o(\PWMA/n13 [23]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMA/mux0_b24  (
    .i0(\PWMA/n12 [24]),
    .i1(freqA[24]),
    .sel(\PWMA/n0 ),
    .o(\PWMA/n13 [24]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMA/mux0_b25  (
    .i0(\PWMA/n12 [25]),
    .i1(freqA[25]),
    .sel(\PWMA/n0 ),
    .o(\PWMA/n13 [25]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMA/mux0_b26  (
    .i0(\PWMA/n12 [26]),
    .i1(freqA[26]),
    .sel(\PWMA/n0 ),
    .o(\PWMA/n13 [26]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMA/mux0_b3  (
    .i0(\PWMA/n12 [3]),
    .i1(freqA[3]),
    .sel(\PWMA/n0 ),
    .o(\PWMA/n13 [3]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMA/mux0_b4  (
    .i0(\PWMA/n12 [4]),
    .i1(freqA[4]),
    .sel(\PWMA/n0 ),
    .o(\PWMA/n13 [4]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMA/mux0_b5  (
    .i0(\PWMA/n12 [5]),
    .i1(freqA[5]),
    .sel(\PWMA/n0 ),
    .o(\PWMA/n13 [5]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMA/mux0_b6  (
    .i0(\PWMA/n12 [6]),
    .i1(freqA[6]),
    .sel(\PWMA/n0 ),
    .o(\PWMA/n13 [6]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMA/mux0_b7  (
    .i0(\PWMA/n12 [7]),
    .i1(freqA[7]),
    .sel(\PWMA/n0 ),
    .o(\PWMA/n13 [7]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMA/mux0_b8  (
    .i0(\PWMA/n12 [8]),
    .i1(freqA[8]),
    .sel(\PWMA/n0 ),
    .o(\PWMA/n13 [8]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMA/mux0_b9  (
    .i0(\PWMA/n12 [9]),
    .i1(freqA[9]),
    .sel(\PWMA/n0 ),
    .o(\PWMA/n13 [9]));  // src/OnePWM.v(32)
  and \PWMA/mux3_b0_sel_is_3  (\PWMA/mux3_b0_sel_is_3_o , \PWMA/n11 , \PWMA/n0 );
  binary_mux_s1_w1 \PWMA/mux4_b0  (
    .i0(\PWMA/pnumr [0]),
    .i1(1'b0),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n22 [0]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux4_b1  (
    .i0(\PWMA/pnumr [1]),
    .i1(1'b0),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n22 [1]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux4_b10  (
    .i0(\PWMA/pnumr [10]),
    .i1(1'b0),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n22 [10]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux4_b11  (
    .i0(\PWMA/pnumr [11]),
    .i1(1'b0),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n22 [11]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux4_b12  (
    .i0(\PWMA/pnumr [12]),
    .i1(1'b0),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n22 [12]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux4_b13  (
    .i0(\PWMA/pnumr [13]),
    .i1(1'b0),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n22 [13]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux4_b14  (
    .i0(\PWMA/pnumr [14]),
    .i1(1'b0),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n22 [14]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux4_b15  (
    .i0(\PWMA/pnumr [15]),
    .i1(1'b0),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n22 [15]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux4_b16  (
    .i0(\PWMA/pnumr [16]),
    .i1(1'b0),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n22 [16]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux4_b17  (
    .i0(\PWMA/pnumr [17]),
    .i1(1'b0),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n22 [17]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux4_b18  (
    .i0(\PWMA/pnumr [18]),
    .i1(1'b0),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n22 [18]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux4_b19  (
    .i0(\PWMA/pnumr [19]),
    .i1(1'b0),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n22 [19]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux4_b2  (
    .i0(\PWMA/pnumr [2]),
    .i1(1'b0),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n22 [2]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux4_b20  (
    .i0(\PWMA/pnumr [20]),
    .i1(1'b0),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n22 [20]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux4_b21  (
    .i0(\PWMA/pnumr [21]),
    .i1(1'b0),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n22 [21]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux4_b22  (
    .i0(\PWMA/pnumr [22]),
    .i1(1'b0),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n22 [22]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux4_b23  (
    .i0(\PWMA/pnumr [23]),
    .i1(1'b0),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n22 [23]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux4_b24  (
    .i0(\PWMA/pnumr [24]),
    .i1(1'b0),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n22 [24]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux4_b25  (
    .i0(\PWMA/pnumr [25]),
    .i1(1'b0),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n22 [25]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux4_b26  (
    .i0(\PWMA/pnumr [26]),
    .i1(1'b0),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n22 [26]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux4_b27  (
    .i0(\PWMA/pnumr [27]),
    .i1(1'b0),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n22 [27]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux4_b28  (
    .i0(\PWMA/pnumr [28]),
    .i1(1'b0),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n22 [28]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux4_b29  (
    .i0(\PWMA/pnumr [29]),
    .i1(1'b0),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n22 [29]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux4_b3  (
    .i0(\PWMA/pnumr [3]),
    .i1(1'b0),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n22 [3]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux4_b30  (
    .i0(\PWMA/pnumr [30]),
    .i1(1'b0),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n22 [30]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux4_b31  (
    .i0(\PWMA/pnumr [31]),
    .i1(1'b0),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n22 [31]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux4_b4  (
    .i0(\PWMA/pnumr [4]),
    .i1(1'b0),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n22 [4]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux4_b5  (
    .i0(\PWMA/pnumr [5]),
    .i1(1'b0),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n22 [5]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux4_b6  (
    .i0(\PWMA/pnumr [6]),
    .i1(1'b0),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n22 [6]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux4_b7  (
    .i0(\PWMA/pnumr [7]),
    .i1(1'b0),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n22 [7]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux4_b8  (
    .i0(\PWMA/pnumr [8]),
    .i1(1'b0),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n22 [8]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux4_b9  (
    .i0(\PWMA/pnumr [9]),
    .i1(1'b0),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n22 [9]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux5_b0  (
    .i0(\PWMA/n22 [0]),
    .i1(pnumA[0]),
    .sel(pnumA[32]),
    .o(\PWMA/n23 [0]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux5_b1  (
    .i0(\PWMA/n22 [1]),
    .i1(pnumA[1]),
    .sel(pnumA[32]),
    .o(\PWMA/n23 [1]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux5_b10  (
    .i0(\PWMA/n22 [10]),
    .i1(pnumA[10]),
    .sel(pnumA[32]),
    .o(\PWMA/n23 [10]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux5_b11  (
    .i0(\PWMA/n22 [11]),
    .i1(pnumA[11]),
    .sel(pnumA[32]),
    .o(\PWMA/n23 [11]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux5_b12  (
    .i0(\PWMA/n22 [12]),
    .i1(pnumA[12]),
    .sel(pnumA[32]),
    .o(\PWMA/n23 [12]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux5_b13  (
    .i0(\PWMA/n22 [13]),
    .i1(pnumA[13]),
    .sel(pnumA[32]),
    .o(\PWMA/n23 [13]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux5_b14  (
    .i0(\PWMA/n22 [14]),
    .i1(pnumA[14]),
    .sel(pnumA[32]),
    .o(\PWMA/n23 [14]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux5_b15  (
    .i0(\PWMA/n22 [15]),
    .i1(pnumA[15]),
    .sel(pnumA[32]),
    .o(\PWMA/n23 [15]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux5_b16  (
    .i0(\PWMA/n22 [16]),
    .i1(pnumA[16]),
    .sel(pnumA[32]),
    .o(\PWMA/n23 [16]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux5_b17  (
    .i0(\PWMA/n22 [17]),
    .i1(pnumA[17]),
    .sel(pnumA[32]),
    .o(\PWMA/n23 [17]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux5_b18  (
    .i0(\PWMA/n22 [18]),
    .i1(pnumA[18]),
    .sel(pnumA[32]),
    .o(\PWMA/n23 [18]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux5_b19  (
    .i0(\PWMA/n22 [19]),
    .i1(pnumA[19]),
    .sel(pnumA[32]),
    .o(\PWMA/n23 [19]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux5_b2  (
    .i0(\PWMA/n22 [2]),
    .i1(pnumA[2]),
    .sel(pnumA[32]),
    .o(\PWMA/n23 [2]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux5_b20  (
    .i0(\PWMA/n22 [20]),
    .i1(pnumA[20]),
    .sel(pnumA[32]),
    .o(\PWMA/n23 [20]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux5_b21  (
    .i0(\PWMA/n22 [21]),
    .i1(pnumA[21]),
    .sel(pnumA[32]),
    .o(\PWMA/n23 [21]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux5_b22  (
    .i0(\PWMA/n22 [22]),
    .i1(pnumA[22]),
    .sel(pnumA[32]),
    .o(\PWMA/n23 [22]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux5_b23  (
    .i0(\PWMA/n22 [23]),
    .i1(pnumA[23]),
    .sel(pnumA[32]),
    .o(\PWMA/n23 [23]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux5_b24  (
    .i0(\PWMA/n22 [24]),
    .i1(pnumA[24]),
    .sel(pnumA[32]),
    .o(\PWMA/n23 [24]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux5_b25  (
    .i0(\PWMA/n22 [25]),
    .i1(pnumA[25]),
    .sel(pnumA[32]),
    .o(\PWMA/n23 [25]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux5_b26  (
    .i0(\PWMA/n22 [26]),
    .i1(pnumA[26]),
    .sel(pnumA[32]),
    .o(\PWMA/n23 [26]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux5_b27  (
    .i0(\PWMA/n22 [27]),
    .i1(pnumA[27]),
    .sel(pnumA[32]),
    .o(\PWMA/n23 [27]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux5_b28  (
    .i0(\PWMA/n22 [28]),
    .i1(pnumA[28]),
    .sel(pnumA[32]),
    .o(\PWMA/n23 [28]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux5_b29  (
    .i0(\PWMA/n22 [29]),
    .i1(pnumA[29]),
    .sel(pnumA[32]),
    .o(\PWMA/n23 [29]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux5_b3  (
    .i0(\PWMA/n22 [3]),
    .i1(pnumA[3]),
    .sel(pnumA[32]),
    .o(\PWMA/n23 [3]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux5_b30  (
    .i0(\PWMA/n22 [30]),
    .i1(pnumA[30]),
    .sel(pnumA[32]),
    .o(\PWMA/n23 [30]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux5_b31  (
    .i0(\PWMA/n22 [31]),
    .i1(pnumA[31]),
    .sel(pnumA[32]),
    .o(\PWMA/n23 [31]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux5_b4  (
    .i0(\PWMA/n22 [4]),
    .i1(pnumA[4]),
    .sel(pnumA[32]),
    .o(\PWMA/n23 [4]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux5_b5  (
    .i0(\PWMA/n22 [5]),
    .i1(pnumA[5]),
    .sel(pnumA[32]),
    .o(\PWMA/n23 [5]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux5_b6  (
    .i0(\PWMA/n22 [6]),
    .i1(pnumA[6]),
    .sel(pnumA[32]),
    .o(\PWMA/n23 [6]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux5_b7  (
    .i0(\PWMA/n22 [7]),
    .i1(pnumA[7]),
    .sel(pnumA[32]),
    .o(\PWMA/n23 [7]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux5_b8  (
    .i0(\PWMA/n22 [8]),
    .i1(pnumA[8]),
    .sel(pnumA[32]),
    .o(\PWMA/n23 [8]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux5_b9  (
    .i0(\PWMA/n22 [9]),
    .i1(pnumA[9]),
    .sel(pnumA[32]),
    .o(\PWMA/n23 [9]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMA/mux6_b0  (
    .i0(\PWMA/pnumr [0]),
    .i1(\PWMA/n26 [0]),
    .sel(\PWMA/n25 ),
    .o(\PWMA/n27 [0]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMA/mux6_b1  (
    .i0(\PWMA/pnumr [1]),
    .i1(\PWMA/n26 [1]),
    .sel(\PWMA/n25 ),
    .o(\PWMA/n27 [1]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMA/mux6_b10  (
    .i0(\PWMA/pnumr [10]),
    .i1(\PWMA/n26 [10]),
    .sel(\PWMA/n25 ),
    .o(\PWMA/n27 [10]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMA/mux6_b11  (
    .i0(\PWMA/pnumr [11]),
    .i1(\PWMA/n26 [11]),
    .sel(\PWMA/n25 ),
    .o(\PWMA/n27 [11]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMA/mux6_b12  (
    .i0(\PWMA/pnumr [12]),
    .i1(\PWMA/n26 [12]),
    .sel(\PWMA/n25 ),
    .o(\PWMA/n27 [12]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMA/mux6_b13  (
    .i0(\PWMA/pnumr [13]),
    .i1(\PWMA/n26 [13]),
    .sel(\PWMA/n25 ),
    .o(\PWMA/n27 [13]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMA/mux6_b14  (
    .i0(\PWMA/pnumr [14]),
    .i1(\PWMA/n26 [14]),
    .sel(\PWMA/n25 ),
    .o(\PWMA/n27 [14]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMA/mux6_b15  (
    .i0(\PWMA/pnumr [15]),
    .i1(\PWMA/n26 [15]),
    .sel(\PWMA/n25 ),
    .o(\PWMA/n27 [15]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMA/mux6_b16  (
    .i0(\PWMA/pnumr [16]),
    .i1(\PWMA/n26 [16]),
    .sel(\PWMA/n25 ),
    .o(\PWMA/n27 [16]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMA/mux6_b17  (
    .i0(\PWMA/pnumr [17]),
    .i1(\PWMA/n26 [17]),
    .sel(\PWMA/n25 ),
    .o(\PWMA/n27 [17]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMA/mux6_b18  (
    .i0(\PWMA/pnumr [18]),
    .i1(\PWMA/n26 [18]),
    .sel(\PWMA/n25 ),
    .o(\PWMA/n27 [18]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMA/mux6_b19  (
    .i0(\PWMA/pnumr [19]),
    .i1(\PWMA/n26 [19]),
    .sel(\PWMA/n25 ),
    .o(\PWMA/n27 [19]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMA/mux6_b2  (
    .i0(\PWMA/pnumr [2]),
    .i1(\PWMA/n26 [2]),
    .sel(\PWMA/n25 ),
    .o(\PWMA/n27 [2]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMA/mux6_b20  (
    .i0(\PWMA/pnumr [20]),
    .i1(\PWMA/n26 [20]),
    .sel(\PWMA/n25 ),
    .o(\PWMA/n27 [20]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMA/mux6_b21  (
    .i0(\PWMA/pnumr [21]),
    .i1(\PWMA/n26 [21]),
    .sel(\PWMA/n25 ),
    .o(\PWMA/n27 [21]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMA/mux6_b22  (
    .i0(\PWMA/pnumr [22]),
    .i1(\PWMA/n26 [22]),
    .sel(\PWMA/n25 ),
    .o(\PWMA/n27 [22]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMA/mux6_b23  (
    .i0(\PWMA/pnumr [23]),
    .i1(\PWMA/n26 [23]),
    .sel(\PWMA/n25 ),
    .o(\PWMA/n27 [23]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMA/mux6_b3  (
    .i0(\PWMA/pnumr [3]),
    .i1(\PWMA/n26 [3]),
    .sel(\PWMA/n25 ),
    .o(\PWMA/n27 [3]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMA/mux6_b4  (
    .i0(\PWMA/pnumr [4]),
    .i1(\PWMA/n26 [4]),
    .sel(\PWMA/n25 ),
    .o(\PWMA/n27 [4]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMA/mux6_b5  (
    .i0(\PWMA/pnumr [5]),
    .i1(\PWMA/n26 [5]),
    .sel(\PWMA/n25 ),
    .o(\PWMA/n27 [5]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMA/mux6_b6  (
    .i0(\PWMA/pnumr [6]),
    .i1(\PWMA/n26 [6]),
    .sel(\PWMA/n25 ),
    .o(\PWMA/n27 [6]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMA/mux6_b7  (
    .i0(\PWMA/pnumr [7]),
    .i1(\PWMA/n26 [7]),
    .sel(\PWMA/n25 ),
    .o(\PWMA/n27 [7]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMA/mux6_b8  (
    .i0(\PWMA/pnumr [8]),
    .i1(\PWMA/n26 [8]),
    .sel(\PWMA/n25 ),
    .o(\PWMA/n27 [8]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMA/mux6_b9  (
    .i0(\PWMA/pnumr [9]),
    .i1(\PWMA/n26 [9]),
    .sel(\PWMA/n25 ),
    .o(\PWMA/n27 [9]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMA/mux7_b0  (
    .i0(pnumcntA[0]),
    .i1(\PWMA/n27 [0]),
    .sel(\PWMA/n24 ),
    .o(\PWMA/n29 [0]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux7_b1  (
    .i0(pnumcntA[1]),
    .i1(\PWMA/n27 [1]),
    .sel(\PWMA/n24 ),
    .o(\PWMA/n29 [1]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux7_b10  (
    .i0(pnumcntA[10]),
    .i1(\PWMA/n27 [10]),
    .sel(\PWMA/n24 ),
    .o(\PWMA/n29 [10]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux7_b11  (
    .i0(pnumcntA[11]),
    .i1(\PWMA/n27 [11]),
    .sel(\PWMA/n24 ),
    .o(\PWMA/n29 [11]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux7_b12  (
    .i0(pnumcntA[12]),
    .i1(\PWMA/n27 [12]),
    .sel(\PWMA/n24 ),
    .o(\PWMA/n29 [12]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux7_b13  (
    .i0(pnumcntA[13]),
    .i1(\PWMA/n27 [13]),
    .sel(\PWMA/n24 ),
    .o(\PWMA/n29 [13]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux7_b14  (
    .i0(pnumcntA[14]),
    .i1(\PWMA/n27 [14]),
    .sel(\PWMA/n24 ),
    .o(\PWMA/n29 [14]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux7_b15  (
    .i0(pnumcntA[15]),
    .i1(\PWMA/n27 [15]),
    .sel(\PWMA/n24 ),
    .o(\PWMA/n29 [15]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux7_b16  (
    .i0(pnumcntA[16]),
    .i1(\PWMA/n27 [16]),
    .sel(\PWMA/n24 ),
    .o(\PWMA/n29 [16]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux7_b17  (
    .i0(pnumcntA[17]),
    .i1(\PWMA/n27 [17]),
    .sel(\PWMA/n24 ),
    .o(\PWMA/n29 [17]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux7_b18  (
    .i0(pnumcntA[18]),
    .i1(\PWMA/n27 [18]),
    .sel(\PWMA/n24 ),
    .o(\PWMA/n29 [18]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux7_b19  (
    .i0(pnumcntA[19]),
    .i1(\PWMA/n27 [19]),
    .sel(\PWMA/n24 ),
    .o(\PWMA/n29 [19]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux7_b2  (
    .i0(pnumcntA[2]),
    .i1(\PWMA/n27 [2]),
    .sel(\PWMA/n24 ),
    .o(\PWMA/n29 [2]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux7_b20  (
    .i0(pnumcntA[20]),
    .i1(\PWMA/n27 [20]),
    .sel(\PWMA/n24 ),
    .o(\PWMA/n29 [20]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux7_b21  (
    .i0(pnumcntA[21]),
    .i1(\PWMA/n27 [21]),
    .sel(\PWMA/n24 ),
    .o(\PWMA/n29 [21]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux7_b22  (
    .i0(pnumcntA[22]),
    .i1(\PWMA/n27 [22]),
    .sel(\PWMA/n24 ),
    .o(\PWMA/n29 [22]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux7_b23  (
    .i0(pnumcntA[23]),
    .i1(\PWMA/n27 [23]),
    .sel(\PWMA/n24 ),
    .o(\PWMA/n29 [23]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux7_b3  (
    .i0(pnumcntA[3]),
    .i1(\PWMA/n27 [3]),
    .sel(\PWMA/n24 ),
    .o(\PWMA/n29 [3]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux7_b4  (
    .i0(pnumcntA[4]),
    .i1(\PWMA/n27 [4]),
    .sel(\PWMA/n24 ),
    .o(\PWMA/n29 [4]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux7_b5  (
    .i0(pnumcntA[5]),
    .i1(\PWMA/n27 [5]),
    .sel(\PWMA/n24 ),
    .o(\PWMA/n29 [5]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux7_b6  (
    .i0(pnumcntA[6]),
    .i1(\PWMA/n27 [6]),
    .sel(\PWMA/n24 ),
    .o(\PWMA/n29 [6]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux7_b7  (
    .i0(pnumcntA[7]),
    .i1(\PWMA/n27 [7]),
    .sel(\PWMA/n24 ),
    .o(\PWMA/n29 [7]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux7_b8  (
    .i0(pnumcntA[8]),
    .i1(\PWMA/n27 [8]),
    .sel(\PWMA/n24 ),
    .o(\PWMA/n29 [8]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux7_b9  (
    .i0(pnumcntA[9]),
    .i1(\PWMA/n27 [9]),
    .sel(\PWMA/n24 ),
    .o(\PWMA/n29 [9]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux8_b0  (
    .i0(\PWMA/n29 [0]),
    .i1(\PWMA/pnumr [0]),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n31 [0]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux8_b1  (
    .i0(\PWMA/n29 [1]),
    .i1(\PWMA/pnumr [1]),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n31 [1]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux8_b10  (
    .i0(\PWMA/n29 [10]),
    .i1(\PWMA/pnumr [10]),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n31 [10]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux8_b11  (
    .i0(\PWMA/n29 [11]),
    .i1(\PWMA/pnumr [11]),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n31 [11]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux8_b12  (
    .i0(\PWMA/n29 [12]),
    .i1(\PWMA/pnumr [12]),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n31 [12]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux8_b13  (
    .i0(\PWMA/n29 [13]),
    .i1(\PWMA/pnumr [13]),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n31 [13]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux8_b14  (
    .i0(\PWMA/n29 [14]),
    .i1(\PWMA/pnumr [14]),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n31 [14]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux8_b15  (
    .i0(\PWMA/n29 [15]),
    .i1(\PWMA/pnumr [15]),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n31 [15]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux8_b16  (
    .i0(\PWMA/n29 [16]),
    .i1(\PWMA/pnumr [16]),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n31 [16]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux8_b17  (
    .i0(\PWMA/n29 [17]),
    .i1(\PWMA/pnumr [17]),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n31 [17]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux8_b18  (
    .i0(\PWMA/n29 [18]),
    .i1(\PWMA/pnumr [18]),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n31 [18]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux8_b19  (
    .i0(\PWMA/n29 [19]),
    .i1(\PWMA/pnumr [19]),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n31 [19]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux8_b2  (
    .i0(\PWMA/n29 [2]),
    .i1(\PWMA/pnumr [2]),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n31 [2]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux8_b20  (
    .i0(\PWMA/n29 [20]),
    .i1(\PWMA/pnumr [20]),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n31 [20]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux8_b21  (
    .i0(\PWMA/n29 [21]),
    .i1(\PWMA/pnumr [21]),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n31 [21]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux8_b22  (
    .i0(\PWMA/n29 [22]),
    .i1(\PWMA/pnumr [22]),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n31 [22]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux8_b23  (
    .i0(\PWMA/n29 [23]),
    .i1(\PWMA/pnumr [23]),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n31 [23]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux8_b3  (
    .i0(\PWMA/n29 [3]),
    .i1(\PWMA/pnumr [3]),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n31 [3]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux8_b4  (
    .i0(\PWMA/n29 [4]),
    .i1(\PWMA/pnumr [4]),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n31 [4]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux8_b5  (
    .i0(\PWMA/n29 [5]),
    .i1(\PWMA/pnumr [5]),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n31 [5]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux8_b6  (
    .i0(\PWMA/n29 [6]),
    .i1(\PWMA/pnumr [6]),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n31 [6]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux8_b7  (
    .i0(\PWMA/n29 [7]),
    .i1(\PWMA/pnumr [7]),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n31 [7]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux8_b8  (
    .i0(\PWMA/n29 [8]),
    .i1(\PWMA/pnumr [8]),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n31 [8]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMA/mux8_b9  (
    .i0(\PWMA/n29 [9]),
    .i1(\PWMA/pnumr [9]),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n31 [9]));  // src/OnePWM.v(57)
  not \PWMA/n17_inv  (\PWMA/n17_neg , \PWMA/n17 );
  not \PWMA/n25_inv  (\PWMA/n25_neg , \PWMA/n25 );
  not \PWMA/n4_inv  (\PWMA/n4_neg , \PWMA/n4 );
  not \PWMA/n6_inv  (\PWMA/n6_neg , \PWMA/n6 );
  ne_w24 \PWMA/neq0  (
    .i0(pnumcntA),
    .i1(24'b000000000000000000000000),
    .o(\PWMA/n25 ));  // src/OnePWM.v(55)
  reg_sr_ss_w1 \PWMA/pwm_reg  (
    .clk(clk100m),
    .d(pwm[10]),
    .en(1'b1),
    .reset(~\PWMA/u14_sel_is_1_o ),
    .set(\PWMA/n18 ),
    .q(\PWMA/pwm_keep ));  // src/OnePWM.v(45)
  reg_sr_as_w1 \PWMA/reg0_b0  (
    .clk(clk100m),
    .d(\PWMA/n13 [0]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [0]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b1  (
    .clk(clk100m),
    .d(\PWMA/n13 [1]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [1]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b10  (
    .clk(clk100m),
    .d(\PWMA/n13 [10]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [10]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b11  (
    .clk(clk100m),
    .d(\PWMA/n13 [11]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [11]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b12  (
    .clk(clk100m),
    .d(\PWMA/n13 [12]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [12]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b13  (
    .clk(clk100m),
    .d(\PWMA/n13 [13]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [13]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b14  (
    .clk(clk100m),
    .d(\PWMA/n13 [14]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [14]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b15  (
    .clk(clk100m),
    .d(\PWMA/n13 [15]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [15]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b16  (
    .clk(clk100m),
    .d(\PWMA/n13 [16]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [16]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b17  (
    .clk(clk100m),
    .d(\PWMA/n13 [17]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [17]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b18  (
    .clk(clk100m),
    .d(\PWMA/n13 [18]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [18]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b19  (
    .clk(clk100m),
    .d(\PWMA/n13 [19]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [19]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b2  (
    .clk(clk100m),
    .d(\PWMA/n13 [2]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [2]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b20  (
    .clk(clk100m),
    .d(\PWMA/n13 [20]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [20]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b21  (
    .clk(clk100m),
    .d(\PWMA/n13 [21]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [21]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b22  (
    .clk(clk100m),
    .d(\PWMA/n13 [22]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [22]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b23  (
    .clk(clk100m),
    .d(\PWMA/n13 [23]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [23]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b24  (
    .clk(clk100m),
    .d(\PWMA/n13 [24]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [24]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b25  (
    .clk(clk100m),
    .d(\PWMA/n13 [25]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [25]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b26  (
    .clk(clk100m),
    .d(\PWMA/n13 [26]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [26]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b3  (
    .clk(clk100m),
    .d(\PWMA/n13 [3]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [3]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b4  (
    .clk(clk100m),
    .d(\PWMA/n13 [4]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [4]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b5  (
    .clk(clk100m),
    .d(\PWMA/n13 [5]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [5]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b6  (
    .clk(clk100m),
    .d(\PWMA/n13 [6]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [6]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b7  (
    .clk(clk100m),
    .d(\PWMA/n13 [7]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [7]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b8  (
    .clk(clk100m),
    .d(\PWMA/n13 [8]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [8]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMA/reg0_b9  (
    .clk(clk100m),
    .d(\PWMA/n13 [9]),
    .en(1'b1),
    .reset(~\PWMA/n11 ),
    .set(1'b0),
    .q(\PWMA/FreCnt [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b0  (
    .clk(clk100m),
    .d(freqA[0]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [0]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b1  (
    .clk(clk100m),
    .d(freqA[1]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [1]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b10  (
    .clk(clk100m),
    .d(freqA[10]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [10]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b11  (
    .clk(clk100m),
    .d(freqA[11]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [11]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b12  (
    .clk(clk100m),
    .d(freqA[12]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [12]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b13  (
    .clk(clk100m),
    .d(freqA[13]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [13]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b14  (
    .clk(clk100m),
    .d(freqA[14]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [14]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b15  (
    .clk(clk100m),
    .d(freqA[15]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [15]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b16  (
    .clk(clk100m),
    .d(freqA[16]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [16]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b17  (
    .clk(clk100m),
    .d(freqA[17]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [17]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b18  (
    .clk(clk100m),
    .d(freqA[18]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [18]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b19  (
    .clk(clk100m),
    .d(freqA[19]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [19]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b2  (
    .clk(clk100m),
    .d(freqA[2]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [2]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b20  (
    .clk(clk100m),
    .d(freqA[20]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [20]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b21  (
    .clk(clk100m),
    .d(freqA[21]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [21]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b22  (
    .clk(clk100m),
    .d(freqA[22]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [22]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b23  (
    .clk(clk100m),
    .d(freqA[23]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [23]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b24  (
    .clk(clk100m),
    .d(freqA[24]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [24]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b25  (
    .clk(clk100m),
    .d(freqA[25]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [25]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b26  (
    .clk(clk100m),
    .d(freqA[26]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [26]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b3  (
    .clk(clk100m),
    .d(freqA[3]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [3]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b4  (
    .clk(clk100m),
    .d(freqA[4]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [4]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b5  (
    .clk(clk100m),
    .d(freqA[5]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [5]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b6  (
    .clk(clk100m),
    .d(freqA[6]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [6]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b7  (
    .clk(clk100m),
    .d(freqA[7]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [7]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b8  (
    .clk(clk100m),
    .d(freqA[8]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [8]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg1_b9  (
    .clk(clk100m),
    .d(freqA[9]),
    .en(\PWMA/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/FreCntr [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMA/reg2_b0  (
    .clk(clk100m),
    .d(\PWMA/n23 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[0]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b1  (
    .clk(clk100m),
    .d(\PWMA/n23 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[1]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b10  (
    .clk(clk100m),
    .d(\PWMA/n23 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[10]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b11  (
    .clk(clk100m),
    .d(\PWMA/n23 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[11]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b12  (
    .clk(clk100m),
    .d(\PWMA/n23 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[12]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b13  (
    .clk(clk100m),
    .d(\PWMA/n23 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[13]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b14  (
    .clk(clk100m),
    .d(\PWMA/n23 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[14]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b15  (
    .clk(clk100m),
    .d(\PWMA/n23 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[15]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b16  (
    .clk(clk100m),
    .d(\PWMA/n23 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[16]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b17  (
    .clk(clk100m),
    .d(\PWMA/n23 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[17]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b18  (
    .clk(clk100m),
    .d(\PWMA/n23 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[18]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b19  (
    .clk(clk100m),
    .d(\PWMA/n23 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[19]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b2  (
    .clk(clk100m),
    .d(\PWMA/n23 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[2]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b20  (
    .clk(clk100m),
    .d(\PWMA/n23 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[20]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b21  (
    .clk(clk100m),
    .d(\PWMA/n23 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[21]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b22  (
    .clk(clk100m),
    .d(\PWMA/n23 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[22]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b23  (
    .clk(clk100m),
    .d(\PWMA/n23 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[23]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b24  (
    .clk(clk100m),
    .d(\PWMA/n23 [24]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[24]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b25  (
    .clk(clk100m),
    .d(\PWMA/n23 [25]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[25]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b26  (
    .clk(clk100m),
    .d(\PWMA/n23 [26]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[26]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b27  (
    .clk(clk100m),
    .d(\PWMA/n23 [27]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[27]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b28  (
    .clk(clk100m),
    .d(\PWMA/n23 [28]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[28]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b29  (
    .clk(clk100m),
    .d(\PWMA/n23 [29]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[29]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b3  (
    .clk(clk100m),
    .d(\PWMA/n23 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[3]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b30  (
    .clk(clk100m),
    .d(\PWMA/n23 [30]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[30]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b31  (
    .clk(clk100m),
    .d(\PWMA/n23 [31]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[31]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b4  (
    .clk(clk100m),
    .d(\PWMA/n23 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[4]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b5  (
    .clk(clk100m),
    .d(\PWMA/n23 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[5]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b6  (
    .clk(clk100m),
    .d(\PWMA/n23 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[6]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b7  (
    .clk(clk100m),
    .d(\PWMA/n23 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[7]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b8  (
    .clk(clk100m),
    .d(\PWMA/n23 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[8]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg2_b9  (
    .clk(clk100m),
    .d(\PWMA/n23 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/pnumr[9]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMA/reg3_b0  (
    .clk(clk100m),
    .d(\PWMA/n31 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[0]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b1  (
    .clk(clk100m),
    .d(\PWMA/n31 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[1]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b10  (
    .clk(clk100m),
    .d(\PWMA/n31 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[10]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b11  (
    .clk(clk100m),
    .d(\PWMA/n31 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[11]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b12  (
    .clk(clk100m),
    .d(\PWMA/n31 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[12]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b13  (
    .clk(clk100m),
    .d(\PWMA/n31 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[13]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b14  (
    .clk(clk100m),
    .d(\PWMA/n31 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[14]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b15  (
    .clk(clk100m),
    .d(\PWMA/n31 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[15]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b16  (
    .clk(clk100m),
    .d(\PWMA/n31 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[16]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b17  (
    .clk(clk100m),
    .d(\PWMA/n31 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[17]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b18  (
    .clk(clk100m),
    .d(\PWMA/n31 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[18]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b19  (
    .clk(clk100m),
    .d(\PWMA/n31 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[19]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b2  (
    .clk(clk100m),
    .d(\PWMA/n31 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[2]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b20  (
    .clk(clk100m),
    .d(\PWMA/n31 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[20]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b21  (
    .clk(clk100m),
    .d(\PWMA/n31 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[21]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b22  (
    .clk(clk100m),
    .d(\PWMA/n31 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[22]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b23  (
    .clk(clk100m),
    .d(\PWMA/n31 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[23]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b3  (
    .clk(clk100m),
    .d(\PWMA/n31 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[3]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b4  (
    .clk(clk100m),
    .d(\PWMA/n31 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[4]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b5  (
    .clk(clk100m),
    .d(\PWMA/n31 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[5]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b6  (
    .clk(clk100m),
    .d(\PWMA/n31 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[6]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b7  (
    .clk(clk100m),
    .d(\PWMA/n31 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[7]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b8  (
    .clk(clk100m),
    .d(\PWMA/n31 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[8]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMA/reg3_b9  (
    .clk(clk100m),
    .d(\PWMA/n31 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMA/RemaTxNum[9]_keep ));  // src/OnePWM.v(58)
  reg_ar_ss_w1 \PWMA/stopreq_reg  (
    .clk(clk100m),
    .d(\PWMA/n1 ),
    .en(1'b1),
    .reset(1'b0),
    .set(pwm_start_stop[10]),
    .q(\PWMA/stopreq_keep ));  // src/OnePWM.v(15)
  add_pu27_mu27_o27 \PWMA/sub0  (
    .i0(\PWMA/FreCnt ),
    .i1(27'b000000000000000000000000001),
    .o(\PWMA/n12 [26:0]));  // src/OnePWM.v(32)
  add_pu24_mu24_o24 \PWMA/sub1  (
    .i0(pnumcntA),
    .i1(24'b000000000000000000000001),
    .o(\PWMA/n26 [23:0]));  // src/OnePWM.v(55)
  AL_MUX \PWMA/u10  (
    .i0(1'b0),
    .i1(\PWMA/n9 ),
    .sel(n21),
    .o(\PWMA/n10 ));  // src/OnePWM.v(26)
  or \PWMA/u11  (\PWMA/n11 , pwm_state_read[10], pwm_start_stop[26]);  // src/OnePWM.v(30)
  and \PWMA/u14_sel_is_1  (\PWMA/u14_sel_is_1_o , pwm_state_read[10], \PWMA/n17_neg );
  and \PWMA/u15  (\PWMA/n24 , \PWMA/n0 , pwm_state_read[10]);  // src/OnePWM.v(54)
  and \PWMA/u17_sel_is_1  (\PWMA/u17_sel_is_1_o , \PWMA/n24 , \PWMA/n25_neg );
  not \PWMA/u17_sel_is_1_o_inv  (\PWMA/u17_sel_is_1_o_neg , \PWMA/u17_sel_is_1_o );
  AL_MUX \PWMA/u18  (
    .i0(\PWMA/pnumr [31]),
    .i1(dir[10]),
    .sel(\PWMA/u18_sel_is_0_o ),
    .o(\PWMA/n32 ));
  and \PWMA/u18_sel_is_0  (\PWMA/u18_sel_is_0_o , \pwm_start_stop[26]_neg , \PWMA/u17_sel_is_1_o_neg );
  AL_MUX \PWMA/u2  (
    .i0(\PWMA/stopreq ),
    .i1(1'b0),
    .sel(\PWMA/n0 ),
    .o(\PWMA/n1 ));  // src/OnePWM.v(15)
  and \PWMA/u5  (\PWMA/n4 , \PWMA/stopreq , \PWMA/n0 );  // src/OnePWM.v(23)
  and \PWMA/u6  (\PWMA/n6 , \PWMA/n5 , \PWMA/n0 );  // src/OnePWM.v(25)
  AL_MUX \PWMA/u8  (
    .i0(1'b0),
    .i1(pwm_state_read[10]),
    .sel(\PWMA/u8_sel_is_0_o ),
    .o(\PWMA/n8 ));
  and \PWMA/u8_sel_is_0  (\PWMA/u8_sel_is_0_o , \PWMA/n4_neg , \PWMA/n6_neg );
  AL_MUX \PWMA/u9  (
    .i0(\PWMA/n8 ),
    .i1(1'b1),
    .sel(pwm_start_stop[26]),
    .o(\PWMA/n9 ));  // src/OnePWM.v(26)
  reg_ar_as_w1 \PWMB/State_reg  (
    .clk(clk100m),
    .d(\PWMB/n10 ),
    .en(1'b1),
    .reset(~rstn),
    .set(1'b0),
    .q(pwm_state_read[11]));  // src/OnePWM.v(26)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[0]  (
    .i(\PWMB/RemaTxNum[0]_keep ),
    .o(pnumcntB[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[10]  (
    .i(\PWMB/RemaTxNum[10]_keep ),
    .o(pnumcntB[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[11]  (
    .i(\PWMB/RemaTxNum[11]_keep ),
    .o(pnumcntB[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[12]  (
    .i(\PWMB/RemaTxNum[12]_keep ),
    .o(pnumcntB[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[13]  (
    .i(\PWMB/RemaTxNum[13]_keep ),
    .o(pnumcntB[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[14]  (
    .i(\PWMB/RemaTxNum[14]_keep ),
    .o(pnumcntB[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[15]  (
    .i(\PWMB/RemaTxNum[15]_keep ),
    .o(pnumcntB[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[16]  (
    .i(\PWMB/RemaTxNum[16]_keep ),
    .o(pnumcntB[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[17]  (
    .i(\PWMB/RemaTxNum[17]_keep ),
    .o(pnumcntB[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[18]  (
    .i(\PWMB/RemaTxNum[18]_keep ),
    .o(pnumcntB[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[19]  (
    .i(\PWMB/RemaTxNum[19]_keep ),
    .o(pnumcntB[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[1]  (
    .i(\PWMB/RemaTxNum[1]_keep ),
    .o(pnumcntB[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[20]  (
    .i(\PWMB/RemaTxNum[20]_keep ),
    .o(pnumcntB[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[21]  (
    .i(\PWMB/RemaTxNum[21]_keep ),
    .o(pnumcntB[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[22]  (
    .i(\PWMB/RemaTxNum[22]_keep ),
    .o(pnumcntB[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[23]  (
    .i(\PWMB/RemaTxNum[23]_keep ),
    .o(pnumcntB[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[2]  (
    .i(\PWMB/RemaTxNum[2]_keep ),
    .o(pnumcntB[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[3]  (
    .i(\PWMB/RemaTxNum[3]_keep ),
    .o(pnumcntB[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[4]  (
    .i(\PWMB/RemaTxNum[4]_keep ),
    .o(pnumcntB[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[5]  (
    .i(\PWMB/RemaTxNum[5]_keep ),
    .o(pnumcntB[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[6]  (
    .i(\PWMB/RemaTxNum[6]_keep ),
    .o(pnumcntB[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[7]  (
    .i(\PWMB/RemaTxNum[7]_keep ),
    .o(pnumcntB[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[8]  (
    .i(\PWMB/RemaTxNum[8]_keep ),
    .o(pnumcntB[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_RemaTxNum[9]  (
    .i(\PWMB/RemaTxNum[9]_keep ),
    .o(pnumcntB[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_dir  (
    .i(\PWMB/dir_keep ),
    .o(dir[11]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[0]  (
    .i(\PWMB/pnumr[0]_keep ),
    .o(\PWMB/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[10]  (
    .i(\PWMB/pnumr[10]_keep ),
    .o(\PWMB/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[11]  (
    .i(\PWMB/pnumr[11]_keep ),
    .o(\PWMB/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[12]  (
    .i(\PWMB/pnumr[12]_keep ),
    .o(\PWMB/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[13]  (
    .i(\PWMB/pnumr[13]_keep ),
    .o(\PWMB/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[14]  (
    .i(\PWMB/pnumr[14]_keep ),
    .o(\PWMB/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[15]  (
    .i(\PWMB/pnumr[15]_keep ),
    .o(\PWMB/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[16]  (
    .i(\PWMB/pnumr[16]_keep ),
    .o(\PWMB/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[17]  (
    .i(\PWMB/pnumr[17]_keep ),
    .o(\PWMB/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[18]  (
    .i(\PWMB/pnumr[18]_keep ),
    .o(\PWMB/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[19]  (
    .i(\PWMB/pnumr[19]_keep ),
    .o(\PWMB/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[1]  (
    .i(\PWMB/pnumr[1]_keep ),
    .o(\PWMB/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[20]  (
    .i(\PWMB/pnumr[20]_keep ),
    .o(\PWMB/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[21]  (
    .i(\PWMB/pnumr[21]_keep ),
    .o(\PWMB/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[22]  (
    .i(\PWMB/pnumr[22]_keep ),
    .o(\PWMB/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[23]  (
    .i(\PWMB/pnumr[23]_keep ),
    .o(\PWMB/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[24]  (
    .i(\PWMB/pnumr[24]_keep ),
    .o(\PWMB/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[25]  (
    .i(\PWMB/pnumr[25]_keep ),
    .o(\PWMB/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[26]  (
    .i(\PWMB/pnumr[26]_keep ),
    .o(\PWMB/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[27]  (
    .i(\PWMB/pnumr[27]_keep ),
    .o(\PWMB/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[28]  (
    .i(\PWMB/pnumr[28]_keep ),
    .o(\PWMB/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[29]  (
    .i(\PWMB/pnumr[29]_keep ),
    .o(\PWMB/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[2]  (
    .i(\PWMB/pnumr[2]_keep ),
    .o(\PWMB/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[30]  (
    .i(\PWMB/pnumr[30]_keep ),
    .o(\PWMB/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[31]  (
    .i(\PWMB/pnumr[31]_keep ),
    .o(\PWMB/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[3]  (
    .i(\PWMB/pnumr[3]_keep ),
    .o(\PWMB/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[4]  (
    .i(\PWMB/pnumr[4]_keep ),
    .o(\PWMB/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[5]  (
    .i(\PWMB/pnumr[5]_keep ),
    .o(\PWMB/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[6]  (
    .i(\PWMB/pnumr[6]_keep ),
    .o(\PWMB/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[7]  (
    .i(\PWMB/pnumr[7]_keep ),
    .o(\PWMB/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[8]  (
    .i(\PWMB/pnumr[8]_keep ),
    .o(\PWMB/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pnumr[9]  (
    .i(\PWMB/pnumr[9]_keep ),
    .o(\PWMB/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_pwm  (
    .i(\PWMB/pwm_keep ),
    .o(pwm[11]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMB/_bufkeep_stopreq  (
    .i(\PWMB/stopreq_keep ),
    .o(\PWMB/stopreq ));  // src/OnePWM.v(14)
  reg_ar_as_w1 \PWMB/dir_reg  (
    .clk(clk100m),
    .d(\PWMB/n32 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/dir_keep ));  // src/OnePWM.v(58)
  eq_w27 \PWMB/eq0  (
    .i0(\PWMB/FreCnt ),
    .i1(27'b000000000000000000000000000),
    .o(\PWMB/n0 ));  // src/OnePWM.v(15)
  eq_w24 \PWMB/eq1  (
    .i0(pnumcntB),
    .i1(24'b000000000000000000000001),
    .o(\PWMB/n5 ));  // src/OnePWM.v(25)
  eq_w27 \PWMB/eq2  (
    .i0(\PWMB/FreCnt ),
    .i1({1'b0,\PWMB/FreCntr [26:1]}),
    .o(\PWMB/n17 ));  // src/OnePWM.v(41)
  eq_w27 \PWMB/eq3  (
    .i0(\PWMB/FreCnt ),
    .i1(\PWMB/FreCntr ),
    .o(\PWMB/n18 ));  // src/OnePWM.v(43)
  binary_mux_s1_w1 \PWMB/mux0_b0  (
    .i0(\PWMB/n12 [0]),
    .i1(freqB[0]),
    .sel(\PWMB/n0 ),
    .o(\PWMB/n13 [0]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMB/mux0_b1  (
    .i0(\PWMB/n12 [1]),
    .i1(freqB[1]),
    .sel(\PWMB/n0 ),
    .o(\PWMB/n13 [1]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMB/mux0_b10  (
    .i0(\PWMB/n12 [10]),
    .i1(freqB[10]),
    .sel(\PWMB/n0 ),
    .o(\PWMB/n13 [10]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMB/mux0_b11  (
    .i0(\PWMB/n12 [11]),
    .i1(freqB[11]),
    .sel(\PWMB/n0 ),
    .o(\PWMB/n13 [11]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMB/mux0_b12  (
    .i0(\PWMB/n12 [12]),
    .i1(freqB[12]),
    .sel(\PWMB/n0 ),
    .o(\PWMB/n13 [12]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMB/mux0_b13  (
    .i0(\PWMB/n12 [13]),
    .i1(freqB[13]),
    .sel(\PWMB/n0 ),
    .o(\PWMB/n13 [13]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMB/mux0_b14  (
    .i0(\PWMB/n12 [14]),
    .i1(freqB[14]),
    .sel(\PWMB/n0 ),
    .o(\PWMB/n13 [14]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMB/mux0_b15  (
    .i0(\PWMB/n12 [15]),
    .i1(freqB[15]),
    .sel(\PWMB/n0 ),
    .o(\PWMB/n13 [15]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMB/mux0_b16  (
    .i0(\PWMB/n12 [16]),
    .i1(freqB[16]),
    .sel(\PWMB/n0 ),
    .o(\PWMB/n13 [16]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMB/mux0_b17  (
    .i0(\PWMB/n12 [17]),
    .i1(freqB[17]),
    .sel(\PWMB/n0 ),
    .o(\PWMB/n13 [17]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMB/mux0_b18  (
    .i0(\PWMB/n12 [18]),
    .i1(freqB[18]),
    .sel(\PWMB/n0 ),
    .o(\PWMB/n13 [18]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMB/mux0_b19  (
    .i0(\PWMB/n12 [19]),
    .i1(freqB[19]),
    .sel(\PWMB/n0 ),
    .o(\PWMB/n13 [19]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMB/mux0_b2  (
    .i0(\PWMB/n12 [2]),
    .i1(freqB[2]),
    .sel(\PWMB/n0 ),
    .o(\PWMB/n13 [2]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMB/mux0_b20  (
    .i0(\PWMB/n12 [20]),
    .i1(freqB[20]),
    .sel(\PWMB/n0 ),
    .o(\PWMB/n13 [20]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMB/mux0_b21  (
    .i0(\PWMB/n12 [21]),
    .i1(freqB[21]),
    .sel(\PWMB/n0 ),
    .o(\PWMB/n13 [21]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMB/mux0_b22  (
    .i0(\PWMB/n12 [22]),
    .i1(freqB[22]),
    .sel(\PWMB/n0 ),
    .o(\PWMB/n13 [22]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMB/mux0_b23  (
    .i0(\PWMB/n12 [23]),
    .i1(freqB[23]),
    .sel(\PWMB/n0 ),
    .o(\PWMB/n13 [23]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMB/mux0_b24  (
    .i0(\PWMB/n12 [24]),
    .i1(freqB[24]),
    .sel(\PWMB/n0 ),
    .o(\PWMB/n13 [24]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMB/mux0_b25  (
    .i0(\PWMB/n12 [25]),
    .i1(freqB[25]),
    .sel(\PWMB/n0 ),
    .o(\PWMB/n13 [25]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMB/mux0_b26  (
    .i0(\PWMB/n12 [26]),
    .i1(freqB[26]),
    .sel(\PWMB/n0 ),
    .o(\PWMB/n13 [26]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMB/mux0_b3  (
    .i0(\PWMB/n12 [3]),
    .i1(freqB[3]),
    .sel(\PWMB/n0 ),
    .o(\PWMB/n13 [3]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMB/mux0_b4  (
    .i0(\PWMB/n12 [4]),
    .i1(freqB[4]),
    .sel(\PWMB/n0 ),
    .o(\PWMB/n13 [4]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMB/mux0_b5  (
    .i0(\PWMB/n12 [5]),
    .i1(freqB[5]),
    .sel(\PWMB/n0 ),
    .o(\PWMB/n13 [5]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMB/mux0_b6  (
    .i0(\PWMB/n12 [6]),
    .i1(freqB[6]),
    .sel(\PWMB/n0 ),
    .o(\PWMB/n13 [6]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMB/mux0_b7  (
    .i0(\PWMB/n12 [7]),
    .i1(freqB[7]),
    .sel(\PWMB/n0 ),
    .o(\PWMB/n13 [7]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMB/mux0_b8  (
    .i0(\PWMB/n12 [8]),
    .i1(freqB[8]),
    .sel(\PWMB/n0 ),
    .o(\PWMB/n13 [8]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMB/mux0_b9  (
    .i0(\PWMB/n12 [9]),
    .i1(freqB[9]),
    .sel(\PWMB/n0 ),
    .o(\PWMB/n13 [9]));  // src/OnePWM.v(32)
  and \PWMB/mux3_b0_sel_is_3  (\PWMB/mux3_b0_sel_is_3_o , \PWMB/n11 , \PWMB/n0 );
  binary_mux_s1_w1 \PWMB/mux4_b0  (
    .i0(\PWMB/pnumr [0]),
    .i1(1'b0),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n22 [0]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux4_b1  (
    .i0(\PWMB/pnumr [1]),
    .i1(1'b0),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n22 [1]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux4_b10  (
    .i0(\PWMB/pnumr [10]),
    .i1(1'b0),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n22 [10]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux4_b11  (
    .i0(\PWMB/pnumr [11]),
    .i1(1'b0),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n22 [11]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux4_b12  (
    .i0(\PWMB/pnumr [12]),
    .i1(1'b0),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n22 [12]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux4_b13  (
    .i0(\PWMB/pnumr [13]),
    .i1(1'b0),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n22 [13]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux4_b14  (
    .i0(\PWMB/pnumr [14]),
    .i1(1'b0),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n22 [14]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux4_b15  (
    .i0(\PWMB/pnumr [15]),
    .i1(1'b0),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n22 [15]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux4_b16  (
    .i0(\PWMB/pnumr [16]),
    .i1(1'b0),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n22 [16]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux4_b17  (
    .i0(\PWMB/pnumr [17]),
    .i1(1'b0),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n22 [17]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux4_b18  (
    .i0(\PWMB/pnumr [18]),
    .i1(1'b0),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n22 [18]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux4_b19  (
    .i0(\PWMB/pnumr [19]),
    .i1(1'b0),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n22 [19]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux4_b2  (
    .i0(\PWMB/pnumr [2]),
    .i1(1'b0),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n22 [2]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux4_b20  (
    .i0(\PWMB/pnumr [20]),
    .i1(1'b0),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n22 [20]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux4_b21  (
    .i0(\PWMB/pnumr [21]),
    .i1(1'b0),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n22 [21]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux4_b22  (
    .i0(\PWMB/pnumr [22]),
    .i1(1'b0),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n22 [22]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux4_b23  (
    .i0(\PWMB/pnumr [23]),
    .i1(1'b0),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n22 [23]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux4_b24  (
    .i0(\PWMB/pnumr [24]),
    .i1(1'b0),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n22 [24]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux4_b25  (
    .i0(\PWMB/pnumr [25]),
    .i1(1'b0),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n22 [25]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux4_b26  (
    .i0(\PWMB/pnumr [26]),
    .i1(1'b0),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n22 [26]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux4_b27  (
    .i0(\PWMB/pnumr [27]),
    .i1(1'b0),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n22 [27]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux4_b28  (
    .i0(\PWMB/pnumr [28]),
    .i1(1'b0),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n22 [28]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux4_b29  (
    .i0(\PWMB/pnumr [29]),
    .i1(1'b0),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n22 [29]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux4_b3  (
    .i0(\PWMB/pnumr [3]),
    .i1(1'b0),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n22 [3]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux4_b30  (
    .i0(\PWMB/pnumr [30]),
    .i1(1'b0),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n22 [30]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux4_b31  (
    .i0(\PWMB/pnumr [31]),
    .i1(1'b0),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n22 [31]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux4_b4  (
    .i0(\PWMB/pnumr [4]),
    .i1(1'b0),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n22 [4]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux4_b5  (
    .i0(\PWMB/pnumr [5]),
    .i1(1'b0),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n22 [5]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux4_b6  (
    .i0(\PWMB/pnumr [6]),
    .i1(1'b0),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n22 [6]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux4_b7  (
    .i0(\PWMB/pnumr [7]),
    .i1(1'b0),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n22 [7]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux4_b8  (
    .i0(\PWMB/pnumr [8]),
    .i1(1'b0),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n22 [8]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux4_b9  (
    .i0(\PWMB/pnumr [9]),
    .i1(1'b0),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n22 [9]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux5_b0  (
    .i0(\PWMB/n22 [0]),
    .i1(pnumB[0]),
    .sel(pnumB[32]),
    .o(\PWMB/n23 [0]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux5_b1  (
    .i0(\PWMB/n22 [1]),
    .i1(pnumB[1]),
    .sel(pnumB[32]),
    .o(\PWMB/n23 [1]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux5_b10  (
    .i0(\PWMB/n22 [10]),
    .i1(pnumB[10]),
    .sel(pnumB[32]),
    .o(\PWMB/n23 [10]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux5_b11  (
    .i0(\PWMB/n22 [11]),
    .i1(pnumB[11]),
    .sel(pnumB[32]),
    .o(\PWMB/n23 [11]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux5_b12  (
    .i0(\PWMB/n22 [12]),
    .i1(pnumB[12]),
    .sel(pnumB[32]),
    .o(\PWMB/n23 [12]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux5_b13  (
    .i0(\PWMB/n22 [13]),
    .i1(pnumB[13]),
    .sel(pnumB[32]),
    .o(\PWMB/n23 [13]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux5_b14  (
    .i0(\PWMB/n22 [14]),
    .i1(pnumB[14]),
    .sel(pnumB[32]),
    .o(\PWMB/n23 [14]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux5_b15  (
    .i0(\PWMB/n22 [15]),
    .i1(pnumB[15]),
    .sel(pnumB[32]),
    .o(\PWMB/n23 [15]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux5_b16  (
    .i0(\PWMB/n22 [16]),
    .i1(pnumB[16]),
    .sel(pnumB[32]),
    .o(\PWMB/n23 [16]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux5_b17  (
    .i0(\PWMB/n22 [17]),
    .i1(pnumB[17]),
    .sel(pnumB[32]),
    .o(\PWMB/n23 [17]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux5_b18  (
    .i0(\PWMB/n22 [18]),
    .i1(pnumB[18]),
    .sel(pnumB[32]),
    .o(\PWMB/n23 [18]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux5_b19  (
    .i0(\PWMB/n22 [19]),
    .i1(pnumB[19]),
    .sel(pnumB[32]),
    .o(\PWMB/n23 [19]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux5_b2  (
    .i0(\PWMB/n22 [2]),
    .i1(pnumB[2]),
    .sel(pnumB[32]),
    .o(\PWMB/n23 [2]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux5_b20  (
    .i0(\PWMB/n22 [20]),
    .i1(pnumB[20]),
    .sel(pnumB[32]),
    .o(\PWMB/n23 [20]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux5_b21  (
    .i0(\PWMB/n22 [21]),
    .i1(pnumB[21]),
    .sel(pnumB[32]),
    .o(\PWMB/n23 [21]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux5_b22  (
    .i0(\PWMB/n22 [22]),
    .i1(pnumB[22]),
    .sel(pnumB[32]),
    .o(\PWMB/n23 [22]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux5_b23  (
    .i0(\PWMB/n22 [23]),
    .i1(pnumB[23]),
    .sel(pnumB[32]),
    .o(\PWMB/n23 [23]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux5_b24  (
    .i0(\PWMB/n22 [24]),
    .i1(pnumB[24]),
    .sel(pnumB[32]),
    .o(\PWMB/n23 [24]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux5_b25  (
    .i0(\PWMB/n22 [25]),
    .i1(pnumB[25]),
    .sel(pnumB[32]),
    .o(\PWMB/n23 [25]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux5_b26  (
    .i0(\PWMB/n22 [26]),
    .i1(pnumB[26]),
    .sel(pnumB[32]),
    .o(\PWMB/n23 [26]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux5_b27  (
    .i0(\PWMB/n22 [27]),
    .i1(pnumB[27]),
    .sel(pnumB[32]),
    .o(\PWMB/n23 [27]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux5_b28  (
    .i0(\PWMB/n22 [28]),
    .i1(pnumB[28]),
    .sel(pnumB[32]),
    .o(\PWMB/n23 [28]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux5_b29  (
    .i0(\PWMB/n22 [29]),
    .i1(pnumB[29]),
    .sel(pnumB[32]),
    .o(\PWMB/n23 [29]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux5_b3  (
    .i0(\PWMB/n22 [3]),
    .i1(pnumB[3]),
    .sel(pnumB[32]),
    .o(\PWMB/n23 [3]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux5_b30  (
    .i0(\PWMB/n22 [30]),
    .i1(pnumB[30]),
    .sel(pnumB[32]),
    .o(\PWMB/n23 [30]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux5_b31  (
    .i0(\PWMB/n22 [31]),
    .i1(pnumB[31]),
    .sel(pnumB[32]),
    .o(\PWMB/n23 [31]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux5_b4  (
    .i0(\PWMB/n22 [4]),
    .i1(pnumB[4]),
    .sel(pnumB[32]),
    .o(\PWMB/n23 [4]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux5_b5  (
    .i0(\PWMB/n22 [5]),
    .i1(pnumB[5]),
    .sel(pnumB[32]),
    .o(\PWMB/n23 [5]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux5_b6  (
    .i0(\PWMB/n22 [6]),
    .i1(pnumB[6]),
    .sel(pnumB[32]),
    .o(\PWMB/n23 [6]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux5_b7  (
    .i0(\PWMB/n22 [7]),
    .i1(pnumB[7]),
    .sel(pnumB[32]),
    .o(\PWMB/n23 [7]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux5_b8  (
    .i0(\PWMB/n22 [8]),
    .i1(pnumB[8]),
    .sel(pnumB[32]),
    .o(\PWMB/n23 [8]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux5_b9  (
    .i0(\PWMB/n22 [9]),
    .i1(pnumB[9]),
    .sel(pnumB[32]),
    .o(\PWMB/n23 [9]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMB/mux6_b0  (
    .i0(\PWMB/pnumr [0]),
    .i1(\PWMB/n26 [0]),
    .sel(\PWMB/n25 ),
    .o(\PWMB/n27 [0]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMB/mux6_b1  (
    .i0(\PWMB/pnumr [1]),
    .i1(\PWMB/n26 [1]),
    .sel(\PWMB/n25 ),
    .o(\PWMB/n27 [1]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMB/mux6_b10  (
    .i0(\PWMB/pnumr [10]),
    .i1(\PWMB/n26 [10]),
    .sel(\PWMB/n25 ),
    .o(\PWMB/n27 [10]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMB/mux6_b11  (
    .i0(\PWMB/pnumr [11]),
    .i1(\PWMB/n26 [11]),
    .sel(\PWMB/n25 ),
    .o(\PWMB/n27 [11]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMB/mux6_b12  (
    .i0(\PWMB/pnumr [12]),
    .i1(\PWMB/n26 [12]),
    .sel(\PWMB/n25 ),
    .o(\PWMB/n27 [12]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMB/mux6_b13  (
    .i0(\PWMB/pnumr [13]),
    .i1(\PWMB/n26 [13]),
    .sel(\PWMB/n25 ),
    .o(\PWMB/n27 [13]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMB/mux6_b14  (
    .i0(\PWMB/pnumr [14]),
    .i1(\PWMB/n26 [14]),
    .sel(\PWMB/n25 ),
    .o(\PWMB/n27 [14]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMB/mux6_b15  (
    .i0(\PWMB/pnumr [15]),
    .i1(\PWMB/n26 [15]),
    .sel(\PWMB/n25 ),
    .o(\PWMB/n27 [15]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMB/mux6_b16  (
    .i0(\PWMB/pnumr [16]),
    .i1(\PWMB/n26 [16]),
    .sel(\PWMB/n25 ),
    .o(\PWMB/n27 [16]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMB/mux6_b17  (
    .i0(\PWMB/pnumr [17]),
    .i1(\PWMB/n26 [17]),
    .sel(\PWMB/n25 ),
    .o(\PWMB/n27 [17]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMB/mux6_b18  (
    .i0(\PWMB/pnumr [18]),
    .i1(\PWMB/n26 [18]),
    .sel(\PWMB/n25 ),
    .o(\PWMB/n27 [18]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMB/mux6_b19  (
    .i0(\PWMB/pnumr [19]),
    .i1(\PWMB/n26 [19]),
    .sel(\PWMB/n25 ),
    .o(\PWMB/n27 [19]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMB/mux6_b2  (
    .i0(\PWMB/pnumr [2]),
    .i1(\PWMB/n26 [2]),
    .sel(\PWMB/n25 ),
    .o(\PWMB/n27 [2]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMB/mux6_b20  (
    .i0(\PWMB/pnumr [20]),
    .i1(\PWMB/n26 [20]),
    .sel(\PWMB/n25 ),
    .o(\PWMB/n27 [20]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMB/mux6_b21  (
    .i0(\PWMB/pnumr [21]),
    .i1(\PWMB/n26 [21]),
    .sel(\PWMB/n25 ),
    .o(\PWMB/n27 [21]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMB/mux6_b22  (
    .i0(\PWMB/pnumr [22]),
    .i1(\PWMB/n26 [22]),
    .sel(\PWMB/n25 ),
    .o(\PWMB/n27 [22]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMB/mux6_b23  (
    .i0(\PWMB/pnumr [23]),
    .i1(\PWMB/n26 [23]),
    .sel(\PWMB/n25 ),
    .o(\PWMB/n27 [23]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMB/mux6_b3  (
    .i0(\PWMB/pnumr [3]),
    .i1(\PWMB/n26 [3]),
    .sel(\PWMB/n25 ),
    .o(\PWMB/n27 [3]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMB/mux6_b4  (
    .i0(\PWMB/pnumr [4]),
    .i1(\PWMB/n26 [4]),
    .sel(\PWMB/n25 ),
    .o(\PWMB/n27 [4]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMB/mux6_b5  (
    .i0(\PWMB/pnumr [5]),
    .i1(\PWMB/n26 [5]),
    .sel(\PWMB/n25 ),
    .o(\PWMB/n27 [5]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMB/mux6_b6  (
    .i0(\PWMB/pnumr [6]),
    .i1(\PWMB/n26 [6]),
    .sel(\PWMB/n25 ),
    .o(\PWMB/n27 [6]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMB/mux6_b7  (
    .i0(\PWMB/pnumr [7]),
    .i1(\PWMB/n26 [7]),
    .sel(\PWMB/n25 ),
    .o(\PWMB/n27 [7]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMB/mux6_b8  (
    .i0(\PWMB/pnumr [8]),
    .i1(\PWMB/n26 [8]),
    .sel(\PWMB/n25 ),
    .o(\PWMB/n27 [8]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMB/mux6_b9  (
    .i0(\PWMB/pnumr [9]),
    .i1(\PWMB/n26 [9]),
    .sel(\PWMB/n25 ),
    .o(\PWMB/n27 [9]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMB/mux7_b0  (
    .i0(pnumcntB[0]),
    .i1(\PWMB/n27 [0]),
    .sel(\PWMB/n24 ),
    .o(\PWMB/n29 [0]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux7_b1  (
    .i0(pnumcntB[1]),
    .i1(\PWMB/n27 [1]),
    .sel(\PWMB/n24 ),
    .o(\PWMB/n29 [1]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux7_b10  (
    .i0(pnumcntB[10]),
    .i1(\PWMB/n27 [10]),
    .sel(\PWMB/n24 ),
    .o(\PWMB/n29 [10]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux7_b11  (
    .i0(pnumcntB[11]),
    .i1(\PWMB/n27 [11]),
    .sel(\PWMB/n24 ),
    .o(\PWMB/n29 [11]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux7_b12  (
    .i0(pnumcntB[12]),
    .i1(\PWMB/n27 [12]),
    .sel(\PWMB/n24 ),
    .o(\PWMB/n29 [12]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux7_b13  (
    .i0(pnumcntB[13]),
    .i1(\PWMB/n27 [13]),
    .sel(\PWMB/n24 ),
    .o(\PWMB/n29 [13]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux7_b14  (
    .i0(pnumcntB[14]),
    .i1(\PWMB/n27 [14]),
    .sel(\PWMB/n24 ),
    .o(\PWMB/n29 [14]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux7_b15  (
    .i0(pnumcntB[15]),
    .i1(\PWMB/n27 [15]),
    .sel(\PWMB/n24 ),
    .o(\PWMB/n29 [15]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux7_b16  (
    .i0(pnumcntB[16]),
    .i1(\PWMB/n27 [16]),
    .sel(\PWMB/n24 ),
    .o(\PWMB/n29 [16]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux7_b17  (
    .i0(pnumcntB[17]),
    .i1(\PWMB/n27 [17]),
    .sel(\PWMB/n24 ),
    .o(\PWMB/n29 [17]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux7_b18  (
    .i0(pnumcntB[18]),
    .i1(\PWMB/n27 [18]),
    .sel(\PWMB/n24 ),
    .o(\PWMB/n29 [18]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux7_b19  (
    .i0(pnumcntB[19]),
    .i1(\PWMB/n27 [19]),
    .sel(\PWMB/n24 ),
    .o(\PWMB/n29 [19]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux7_b2  (
    .i0(pnumcntB[2]),
    .i1(\PWMB/n27 [2]),
    .sel(\PWMB/n24 ),
    .o(\PWMB/n29 [2]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux7_b20  (
    .i0(pnumcntB[20]),
    .i1(\PWMB/n27 [20]),
    .sel(\PWMB/n24 ),
    .o(\PWMB/n29 [20]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux7_b21  (
    .i0(pnumcntB[21]),
    .i1(\PWMB/n27 [21]),
    .sel(\PWMB/n24 ),
    .o(\PWMB/n29 [21]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux7_b22  (
    .i0(pnumcntB[22]),
    .i1(\PWMB/n27 [22]),
    .sel(\PWMB/n24 ),
    .o(\PWMB/n29 [22]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux7_b23  (
    .i0(pnumcntB[23]),
    .i1(\PWMB/n27 [23]),
    .sel(\PWMB/n24 ),
    .o(\PWMB/n29 [23]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux7_b3  (
    .i0(pnumcntB[3]),
    .i1(\PWMB/n27 [3]),
    .sel(\PWMB/n24 ),
    .o(\PWMB/n29 [3]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux7_b4  (
    .i0(pnumcntB[4]),
    .i1(\PWMB/n27 [4]),
    .sel(\PWMB/n24 ),
    .o(\PWMB/n29 [4]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux7_b5  (
    .i0(pnumcntB[5]),
    .i1(\PWMB/n27 [5]),
    .sel(\PWMB/n24 ),
    .o(\PWMB/n29 [5]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux7_b6  (
    .i0(pnumcntB[6]),
    .i1(\PWMB/n27 [6]),
    .sel(\PWMB/n24 ),
    .o(\PWMB/n29 [6]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux7_b7  (
    .i0(pnumcntB[7]),
    .i1(\PWMB/n27 [7]),
    .sel(\PWMB/n24 ),
    .o(\PWMB/n29 [7]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux7_b8  (
    .i0(pnumcntB[8]),
    .i1(\PWMB/n27 [8]),
    .sel(\PWMB/n24 ),
    .o(\PWMB/n29 [8]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux7_b9  (
    .i0(pnumcntB[9]),
    .i1(\PWMB/n27 [9]),
    .sel(\PWMB/n24 ),
    .o(\PWMB/n29 [9]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux8_b0  (
    .i0(\PWMB/n29 [0]),
    .i1(\PWMB/pnumr [0]),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n31 [0]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux8_b1  (
    .i0(\PWMB/n29 [1]),
    .i1(\PWMB/pnumr [1]),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n31 [1]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux8_b10  (
    .i0(\PWMB/n29 [10]),
    .i1(\PWMB/pnumr [10]),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n31 [10]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux8_b11  (
    .i0(\PWMB/n29 [11]),
    .i1(\PWMB/pnumr [11]),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n31 [11]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux8_b12  (
    .i0(\PWMB/n29 [12]),
    .i1(\PWMB/pnumr [12]),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n31 [12]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux8_b13  (
    .i0(\PWMB/n29 [13]),
    .i1(\PWMB/pnumr [13]),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n31 [13]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux8_b14  (
    .i0(\PWMB/n29 [14]),
    .i1(\PWMB/pnumr [14]),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n31 [14]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux8_b15  (
    .i0(\PWMB/n29 [15]),
    .i1(\PWMB/pnumr [15]),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n31 [15]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux8_b16  (
    .i0(\PWMB/n29 [16]),
    .i1(\PWMB/pnumr [16]),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n31 [16]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux8_b17  (
    .i0(\PWMB/n29 [17]),
    .i1(\PWMB/pnumr [17]),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n31 [17]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux8_b18  (
    .i0(\PWMB/n29 [18]),
    .i1(\PWMB/pnumr [18]),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n31 [18]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux8_b19  (
    .i0(\PWMB/n29 [19]),
    .i1(\PWMB/pnumr [19]),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n31 [19]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux8_b2  (
    .i0(\PWMB/n29 [2]),
    .i1(\PWMB/pnumr [2]),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n31 [2]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux8_b20  (
    .i0(\PWMB/n29 [20]),
    .i1(\PWMB/pnumr [20]),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n31 [20]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux8_b21  (
    .i0(\PWMB/n29 [21]),
    .i1(\PWMB/pnumr [21]),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n31 [21]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux8_b22  (
    .i0(\PWMB/n29 [22]),
    .i1(\PWMB/pnumr [22]),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n31 [22]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux8_b23  (
    .i0(\PWMB/n29 [23]),
    .i1(\PWMB/pnumr [23]),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n31 [23]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux8_b3  (
    .i0(\PWMB/n29 [3]),
    .i1(\PWMB/pnumr [3]),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n31 [3]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux8_b4  (
    .i0(\PWMB/n29 [4]),
    .i1(\PWMB/pnumr [4]),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n31 [4]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux8_b5  (
    .i0(\PWMB/n29 [5]),
    .i1(\PWMB/pnumr [5]),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n31 [5]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux8_b6  (
    .i0(\PWMB/n29 [6]),
    .i1(\PWMB/pnumr [6]),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n31 [6]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux8_b7  (
    .i0(\PWMB/n29 [7]),
    .i1(\PWMB/pnumr [7]),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n31 [7]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux8_b8  (
    .i0(\PWMB/n29 [8]),
    .i1(\PWMB/pnumr [8]),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n31 [8]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMB/mux8_b9  (
    .i0(\PWMB/n29 [9]),
    .i1(\PWMB/pnumr [9]),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n31 [9]));  // src/OnePWM.v(57)
  not \PWMB/n17_inv  (\PWMB/n17_neg , \PWMB/n17 );
  not \PWMB/n25_inv  (\PWMB/n25_neg , \PWMB/n25 );
  not \PWMB/n4_inv  (\PWMB/n4_neg , \PWMB/n4 );
  not \PWMB/n6_inv  (\PWMB/n6_neg , \PWMB/n6 );
  ne_w24 \PWMB/neq0  (
    .i0(pnumcntB),
    .i1(24'b000000000000000000000000),
    .o(\PWMB/n25 ));  // src/OnePWM.v(55)
  reg_sr_ss_w1 \PWMB/pwm_reg  (
    .clk(clk100m),
    .d(pwm[11]),
    .en(1'b1),
    .reset(~\PWMB/u14_sel_is_1_o ),
    .set(\PWMB/n18 ),
    .q(\PWMB/pwm_keep ));  // src/OnePWM.v(45)
  reg_sr_as_w1 \PWMB/reg0_b0  (
    .clk(clk100m),
    .d(\PWMB/n13 [0]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [0]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b1  (
    .clk(clk100m),
    .d(\PWMB/n13 [1]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [1]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b10  (
    .clk(clk100m),
    .d(\PWMB/n13 [10]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [10]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b11  (
    .clk(clk100m),
    .d(\PWMB/n13 [11]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [11]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b12  (
    .clk(clk100m),
    .d(\PWMB/n13 [12]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [12]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b13  (
    .clk(clk100m),
    .d(\PWMB/n13 [13]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [13]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b14  (
    .clk(clk100m),
    .d(\PWMB/n13 [14]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [14]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b15  (
    .clk(clk100m),
    .d(\PWMB/n13 [15]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [15]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b16  (
    .clk(clk100m),
    .d(\PWMB/n13 [16]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [16]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b17  (
    .clk(clk100m),
    .d(\PWMB/n13 [17]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [17]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b18  (
    .clk(clk100m),
    .d(\PWMB/n13 [18]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [18]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b19  (
    .clk(clk100m),
    .d(\PWMB/n13 [19]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [19]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b2  (
    .clk(clk100m),
    .d(\PWMB/n13 [2]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [2]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b20  (
    .clk(clk100m),
    .d(\PWMB/n13 [20]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [20]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b21  (
    .clk(clk100m),
    .d(\PWMB/n13 [21]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [21]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b22  (
    .clk(clk100m),
    .d(\PWMB/n13 [22]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [22]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b23  (
    .clk(clk100m),
    .d(\PWMB/n13 [23]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [23]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b24  (
    .clk(clk100m),
    .d(\PWMB/n13 [24]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [24]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b25  (
    .clk(clk100m),
    .d(\PWMB/n13 [25]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [25]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b26  (
    .clk(clk100m),
    .d(\PWMB/n13 [26]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [26]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b3  (
    .clk(clk100m),
    .d(\PWMB/n13 [3]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [3]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b4  (
    .clk(clk100m),
    .d(\PWMB/n13 [4]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [4]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b5  (
    .clk(clk100m),
    .d(\PWMB/n13 [5]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [5]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b6  (
    .clk(clk100m),
    .d(\PWMB/n13 [6]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [6]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b7  (
    .clk(clk100m),
    .d(\PWMB/n13 [7]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [7]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b8  (
    .clk(clk100m),
    .d(\PWMB/n13 [8]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [8]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMB/reg0_b9  (
    .clk(clk100m),
    .d(\PWMB/n13 [9]),
    .en(1'b1),
    .reset(~\PWMB/n11 ),
    .set(1'b0),
    .q(\PWMB/FreCnt [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b0  (
    .clk(clk100m),
    .d(freqB[0]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [0]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b1  (
    .clk(clk100m),
    .d(freqB[1]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [1]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b10  (
    .clk(clk100m),
    .d(freqB[10]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [10]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b11  (
    .clk(clk100m),
    .d(freqB[11]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [11]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b12  (
    .clk(clk100m),
    .d(freqB[12]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [12]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b13  (
    .clk(clk100m),
    .d(freqB[13]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [13]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b14  (
    .clk(clk100m),
    .d(freqB[14]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [14]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b15  (
    .clk(clk100m),
    .d(freqB[15]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [15]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b16  (
    .clk(clk100m),
    .d(freqB[16]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [16]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b17  (
    .clk(clk100m),
    .d(freqB[17]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [17]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b18  (
    .clk(clk100m),
    .d(freqB[18]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [18]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b19  (
    .clk(clk100m),
    .d(freqB[19]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [19]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b2  (
    .clk(clk100m),
    .d(freqB[2]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [2]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b20  (
    .clk(clk100m),
    .d(freqB[20]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [20]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b21  (
    .clk(clk100m),
    .d(freqB[21]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [21]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b22  (
    .clk(clk100m),
    .d(freqB[22]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [22]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b23  (
    .clk(clk100m),
    .d(freqB[23]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [23]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b24  (
    .clk(clk100m),
    .d(freqB[24]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [24]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b25  (
    .clk(clk100m),
    .d(freqB[25]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [25]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b26  (
    .clk(clk100m),
    .d(freqB[26]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [26]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b3  (
    .clk(clk100m),
    .d(freqB[3]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [3]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b4  (
    .clk(clk100m),
    .d(freqB[4]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [4]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b5  (
    .clk(clk100m),
    .d(freqB[5]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [5]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b6  (
    .clk(clk100m),
    .d(freqB[6]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [6]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b7  (
    .clk(clk100m),
    .d(freqB[7]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [7]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b8  (
    .clk(clk100m),
    .d(freqB[8]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [8]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg1_b9  (
    .clk(clk100m),
    .d(freqB[9]),
    .en(\PWMB/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/FreCntr [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMB/reg2_b0  (
    .clk(clk100m),
    .d(\PWMB/n23 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[0]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b1  (
    .clk(clk100m),
    .d(\PWMB/n23 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[1]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b10  (
    .clk(clk100m),
    .d(\PWMB/n23 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[10]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b11  (
    .clk(clk100m),
    .d(\PWMB/n23 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[11]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b12  (
    .clk(clk100m),
    .d(\PWMB/n23 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[12]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b13  (
    .clk(clk100m),
    .d(\PWMB/n23 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[13]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b14  (
    .clk(clk100m),
    .d(\PWMB/n23 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[14]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b15  (
    .clk(clk100m),
    .d(\PWMB/n23 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[15]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b16  (
    .clk(clk100m),
    .d(\PWMB/n23 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[16]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b17  (
    .clk(clk100m),
    .d(\PWMB/n23 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[17]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b18  (
    .clk(clk100m),
    .d(\PWMB/n23 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[18]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b19  (
    .clk(clk100m),
    .d(\PWMB/n23 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[19]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b2  (
    .clk(clk100m),
    .d(\PWMB/n23 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[2]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b20  (
    .clk(clk100m),
    .d(\PWMB/n23 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[20]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b21  (
    .clk(clk100m),
    .d(\PWMB/n23 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[21]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b22  (
    .clk(clk100m),
    .d(\PWMB/n23 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[22]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b23  (
    .clk(clk100m),
    .d(\PWMB/n23 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[23]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b24  (
    .clk(clk100m),
    .d(\PWMB/n23 [24]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[24]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b25  (
    .clk(clk100m),
    .d(\PWMB/n23 [25]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[25]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b26  (
    .clk(clk100m),
    .d(\PWMB/n23 [26]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[26]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b27  (
    .clk(clk100m),
    .d(\PWMB/n23 [27]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[27]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b28  (
    .clk(clk100m),
    .d(\PWMB/n23 [28]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[28]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b29  (
    .clk(clk100m),
    .d(\PWMB/n23 [29]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[29]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b3  (
    .clk(clk100m),
    .d(\PWMB/n23 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[3]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b30  (
    .clk(clk100m),
    .d(\PWMB/n23 [30]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[30]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b31  (
    .clk(clk100m),
    .d(\PWMB/n23 [31]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[31]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b4  (
    .clk(clk100m),
    .d(\PWMB/n23 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[4]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b5  (
    .clk(clk100m),
    .d(\PWMB/n23 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[5]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b6  (
    .clk(clk100m),
    .d(\PWMB/n23 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[6]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b7  (
    .clk(clk100m),
    .d(\PWMB/n23 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[7]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b8  (
    .clk(clk100m),
    .d(\PWMB/n23 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[8]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg2_b9  (
    .clk(clk100m),
    .d(\PWMB/n23 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/pnumr[9]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMB/reg3_b0  (
    .clk(clk100m),
    .d(\PWMB/n31 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[0]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b1  (
    .clk(clk100m),
    .d(\PWMB/n31 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[1]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b10  (
    .clk(clk100m),
    .d(\PWMB/n31 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[10]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b11  (
    .clk(clk100m),
    .d(\PWMB/n31 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[11]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b12  (
    .clk(clk100m),
    .d(\PWMB/n31 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[12]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b13  (
    .clk(clk100m),
    .d(\PWMB/n31 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[13]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b14  (
    .clk(clk100m),
    .d(\PWMB/n31 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[14]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b15  (
    .clk(clk100m),
    .d(\PWMB/n31 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[15]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b16  (
    .clk(clk100m),
    .d(\PWMB/n31 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[16]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b17  (
    .clk(clk100m),
    .d(\PWMB/n31 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[17]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b18  (
    .clk(clk100m),
    .d(\PWMB/n31 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[18]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b19  (
    .clk(clk100m),
    .d(\PWMB/n31 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[19]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b2  (
    .clk(clk100m),
    .d(\PWMB/n31 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[2]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b20  (
    .clk(clk100m),
    .d(\PWMB/n31 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[20]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b21  (
    .clk(clk100m),
    .d(\PWMB/n31 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[21]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b22  (
    .clk(clk100m),
    .d(\PWMB/n31 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[22]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b23  (
    .clk(clk100m),
    .d(\PWMB/n31 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[23]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b3  (
    .clk(clk100m),
    .d(\PWMB/n31 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[3]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b4  (
    .clk(clk100m),
    .d(\PWMB/n31 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[4]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b5  (
    .clk(clk100m),
    .d(\PWMB/n31 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[5]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b6  (
    .clk(clk100m),
    .d(\PWMB/n31 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[6]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b7  (
    .clk(clk100m),
    .d(\PWMB/n31 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[7]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b8  (
    .clk(clk100m),
    .d(\PWMB/n31 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[8]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMB/reg3_b9  (
    .clk(clk100m),
    .d(\PWMB/n31 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMB/RemaTxNum[9]_keep ));  // src/OnePWM.v(58)
  reg_ar_ss_w1 \PWMB/stopreq_reg  (
    .clk(clk100m),
    .d(\PWMB/n1 ),
    .en(1'b1),
    .reset(1'b0),
    .set(pwm_start_stop[11]),
    .q(\PWMB/stopreq_keep ));  // src/OnePWM.v(15)
  add_pu27_mu27_o27 \PWMB/sub0  (
    .i0(\PWMB/FreCnt ),
    .i1(27'b000000000000000000000000001),
    .o(\PWMB/n12 [26:0]));  // src/OnePWM.v(32)
  add_pu24_mu24_o24 \PWMB/sub1  (
    .i0(pnumcntB),
    .i1(24'b000000000000000000000001),
    .o(\PWMB/n26 [23:0]));  // src/OnePWM.v(55)
  AL_MUX \PWMB/u10  (
    .i0(1'b0),
    .i1(\PWMB/n9 ),
    .sel(n22),
    .o(\PWMB/n10 ));  // src/OnePWM.v(26)
  or \PWMB/u11  (\PWMB/n11 , pwm_state_read[11], pwm_start_stop[27]);  // src/OnePWM.v(30)
  and \PWMB/u14_sel_is_1  (\PWMB/u14_sel_is_1_o , pwm_state_read[11], \PWMB/n17_neg );
  and \PWMB/u15  (\PWMB/n24 , \PWMB/n0 , pwm_state_read[11]);  // src/OnePWM.v(54)
  and \PWMB/u17_sel_is_1  (\PWMB/u17_sel_is_1_o , \PWMB/n24 , \PWMB/n25_neg );
  not \PWMB/u17_sel_is_1_o_inv  (\PWMB/u17_sel_is_1_o_neg , \PWMB/u17_sel_is_1_o );
  AL_MUX \PWMB/u18  (
    .i0(\PWMB/pnumr [31]),
    .i1(dir[11]),
    .sel(\PWMB/u18_sel_is_0_o ),
    .o(\PWMB/n32 ));
  and \PWMB/u18_sel_is_0  (\PWMB/u18_sel_is_0_o , \pwm_start_stop[27]_neg , \PWMB/u17_sel_is_1_o_neg );
  AL_MUX \PWMB/u2  (
    .i0(\PWMB/stopreq ),
    .i1(1'b0),
    .sel(\PWMB/n0 ),
    .o(\PWMB/n1 ));  // src/OnePWM.v(15)
  and \PWMB/u5  (\PWMB/n4 , \PWMB/stopreq , \PWMB/n0 );  // src/OnePWM.v(23)
  and \PWMB/u6  (\PWMB/n6 , \PWMB/n5 , \PWMB/n0 );  // src/OnePWM.v(25)
  AL_MUX \PWMB/u8  (
    .i0(1'b0),
    .i1(pwm_state_read[11]),
    .sel(\PWMB/u8_sel_is_0_o ),
    .o(\PWMB/n8 ));
  and \PWMB/u8_sel_is_0  (\PWMB/u8_sel_is_0_o , \PWMB/n4_neg , \PWMB/n6_neg );
  AL_MUX \PWMB/u9  (
    .i0(\PWMB/n8 ),
    .i1(1'b1),
    .sel(pwm_start_stop[27]),
    .o(\PWMB/n9 ));  // src/OnePWM.v(26)
  reg_ar_as_w1 \PWMC/State_reg  (
    .clk(clk100m),
    .d(\PWMC/n10 ),
    .en(1'b1),
    .reset(~rstn),
    .set(1'b0),
    .q(pwm_state_read[12]));  // src/OnePWM.v(26)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[0]  (
    .i(\PWMC/RemaTxNum[0]_keep ),
    .o(pnumcntC[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[10]  (
    .i(\PWMC/RemaTxNum[10]_keep ),
    .o(pnumcntC[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[11]  (
    .i(\PWMC/RemaTxNum[11]_keep ),
    .o(pnumcntC[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[12]  (
    .i(\PWMC/RemaTxNum[12]_keep ),
    .o(pnumcntC[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[13]  (
    .i(\PWMC/RemaTxNum[13]_keep ),
    .o(pnumcntC[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[14]  (
    .i(\PWMC/RemaTxNum[14]_keep ),
    .o(pnumcntC[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[15]  (
    .i(\PWMC/RemaTxNum[15]_keep ),
    .o(pnumcntC[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[16]  (
    .i(\PWMC/RemaTxNum[16]_keep ),
    .o(pnumcntC[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[17]  (
    .i(\PWMC/RemaTxNum[17]_keep ),
    .o(pnumcntC[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[18]  (
    .i(\PWMC/RemaTxNum[18]_keep ),
    .o(pnumcntC[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[19]  (
    .i(\PWMC/RemaTxNum[19]_keep ),
    .o(pnumcntC[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[1]  (
    .i(\PWMC/RemaTxNum[1]_keep ),
    .o(pnumcntC[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[20]  (
    .i(\PWMC/RemaTxNum[20]_keep ),
    .o(pnumcntC[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[21]  (
    .i(\PWMC/RemaTxNum[21]_keep ),
    .o(pnumcntC[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[22]  (
    .i(\PWMC/RemaTxNum[22]_keep ),
    .o(pnumcntC[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[23]  (
    .i(\PWMC/RemaTxNum[23]_keep ),
    .o(pnumcntC[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[2]  (
    .i(\PWMC/RemaTxNum[2]_keep ),
    .o(pnumcntC[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[3]  (
    .i(\PWMC/RemaTxNum[3]_keep ),
    .o(pnumcntC[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[4]  (
    .i(\PWMC/RemaTxNum[4]_keep ),
    .o(pnumcntC[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[5]  (
    .i(\PWMC/RemaTxNum[5]_keep ),
    .o(pnumcntC[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[6]  (
    .i(\PWMC/RemaTxNum[6]_keep ),
    .o(pnumcntC[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[7]  (
    .i(\PWMC/RemaTxNum[7]_keep ),
    .o(pnumcntC[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[8]  (
    .i(\PWMC/RemaTxNum[8]_keep ),
    .o(pnumcntC[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_RemaTxNum[9]  (
    .i(\PWMC/RemaTxNum[9]_keep ),
    .o(pnumcntC[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_dir  (
    .i(\PWMC/dir_keep ),
    .o(dir[12]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[0]  (
    .i(\PWMC/pnumr[0]_keep ),
    .o(\PWMC/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[10]  (
    .i(\PWMC/pnumr[10]_keep ),
    .o(\PWMC/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[11]  (
    .i(\PWMC/pnumr[11]_keep ),
    .o(\PWMC/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[12]  (
    .i(\PWMC/pnumr[12]_keep ),
    .o(\PWMC/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[13]  (
    .i(\PWMC/pnumr[13]_keep ),
    .o(\PWMC/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[14]  (
    .i(\PWMC/pnumr[14]_keep ),
    .o(\PWMC/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[15]  (
    .i(\PWMC/pnumr[15]_keep ),
    .o(\PWMC/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[16]  (
    .i(\PWMC/pnumr[16]_keep ),
    .o(\PWMC/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[17]  (
    .i(\PWMC/pnumr[17]_keep ),
    .o(\PWMC/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[18]  (
    .i(\PWMC/pnumr[18]_keep ),
    .o(\PWMC/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[19]  (
    .i(\PWMC/pnumr[19]_keep ),
    .o(\PWMC/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[1]  (
    .i(\PWMC/pnumr[1]_keep ),
    .o(\PWMC/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[20]  (
    .i(\PWMC/pnumr[20]_keep ),
    .o(\PWMC/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[21]  (
    .i(\PWMC/pnumr[21]_keep ),
    .o(\PWMC/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[22]  (
    .i(\PWMC/pnumr[22]_keep ),
    .o(\PWMC/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[23]  (
    .i(\PWMC/pnumr[23]_keep ),
    .o(\PWMC/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[24]  (
    .i(\PWMC/pnumr[24]_keep ),
    .o(\PWMC/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[25]  (
    .i(\PWMC/pnumr[25]_keep ),
    .o(\PWMC/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[26]  (
    .i(\PWMC/pnumr[26]_keep ),
    .o(\PWMC/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[27]  (
    .i(\PWMC/pnumr[27]_keep ),
    .o(\PWMC/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[28]  (
    .i(\PWMC/pnumr[28]_keep ),
    .o(\PWMC/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[29]  (
    .i(\PWMC/pnumr[29]_keep ),
    .o(\PWMC/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[2]  (
    .i(\PWMC/pnumr[2]_keep ),
    .o(\PWMC/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[30]  (
    .i(\PWMC/pnumr[30]_keep ),
    .o(\PWMC/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[31]  (
    .i(\PWMC/pnumr[31]_keep ),
    .o(\PWMC/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[3]  (
    .i(\PWMC/pnumr[3]_keep ),
    .o(\PWMC/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[4]  (
    .i(\PWMC/pnumr[4]_keep ),
    .o(\PWMC/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[5]  (
    .i(\PWMC/pnumr[5]_keep ),
    .o(\PWMC/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[6]  (
    .i(\PWMC/pnumr[6]_keep ),
    .o(\PWMC/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[7]  (
    .i(\PWMC/pnumr[7]_keep ),
    .o(\PWMC/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[8]  (
    .i(\PWMC/pnumr[8]_keep ),
    .o(\PWMC/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pnumr[9]  (
    .i(\PWMC/pnumr[9]_keep ),
    .o(\PWMC/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_pwm  (
    .i(\PWMC/pwm_keep ),
    .o(pwm[12]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMC/_bufkeep_stopreq  (
    .i(\PWMC/stopreq_keep ),
    .o(\PWMC/stopreq ));  // src/OnePWM.v(14)
  reg_ar_as_w1 \PWMC/dir_reg  (
    .clk(clk100m),
    .d(\PWMC/n32 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/dir_keep ));  // src/OnePWM.v(58)
  eq_w27 \PWMC/eq0  (
    .i0(\PWMC/FreCnt ),
    .i1(27'b000000000000000000000000000),
    .o(\PWMC/n0 ));  // src/OnePWM.v(15)
  eq_w24 \PWMC/eq1  (
    .i0(pnumcntC),
    .i1(24'b000000000000000000000001),
    .o(\PWMC/n5 ));  // src/OnePWM.v(25)
  eq_w27 \PWMC/eq2  (
    .i0(\PWMC/FreCnt ),
    .i1({1'b0,\PWMC/FreCntr [26:1]}),
    .o(\PWMC/n17 ));  // src/OnePWM.v(41)
  eq_w27 \PWMC/eq3  (
    .i0(\PWMC/FreCnt ),
    .i1(\PWMC/FreCntr ),
    .o(\PWMC/n18 ));  // src/OnePWM.v(43)
  binary_mux_s1_w1 \PWMC/mux0_b0  (
    .i0(\PWMC/n12 [0]),
    .i1(freqC[0]),
    .sel(\PWMC/n0 ),
    .o(\PWMC/n13 [0]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMC/mux0_b1  (
    .i0(\PWMC/n12 [1]),
    .i1(freqC[1]),
    .sel(\PWMC/n0 ),
    .o(\PWMC/n13 [1]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMC/mux0_b10  (
    .i0(\PWMC/n12 [10]),
    .i1(freqC[10]),
    .sel(\PWMC/n0 ),
    .o(\PWMC/n13 [10]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMC/mux0_b11  (
    .i0(\PWMC/n12 [11]),
    .i1(freqC[11]),
    .sel(\PWMC/n0 ),
    .o(\PWMC/n13 [11]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMC/mux0_b12  (
    .i0(\PWMC/n12 [12]),
    .i1(freqC[12]),
    .sel(\PWMC/n0 ),
    .o(\PWMC/n13 [12]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMC/mux0_b13  (
    .i0(\PWMC/n12 [13]),
    .i1(freqC[13]),
    .sel(\PWMC/n0 ),
    .o(\PWMC/n13 [13]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMC/mux0_b14  (
    .i0(\PWMC/n12 [14]),
    .i1(freqC[14]),
    .sel(\PWMC/n0 ),
    .o(\PWMC/n13 [14]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMC/mux0_b15  (
    .i0(\PWMC/n12 [15]),
    .i1(freqC[15]),
    .sel(\PWMC/n0 ),
    .o(\PWMC/n13 [15]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMC/mux0_b16  (
    .i0(\PWMC/n12 [16]),
    .i1(freqC[16]),
    .sel(\PWMC/n0 ),
    .o(\PWMC/n13 [16]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMC/mux0_b17  (
    .i0(\PWMC/n12 [17]),
    .i1(freqC[17]),
    .sel(\PWMC/n0 ),
    .o(\PWMC/n13 [17]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMC/mux0_b18  (
    .i0(\PWMC/n12 [18]),
    .i1(freqC[18]),
    .sel(\PWMC/n0 ),
    .o(\PWMC/n13 [18]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMC/mux0_b19  (
    .i0(\PWMC/n12 [19]),
    .i1(freqC[19]),
    .sel(\PWMC/n0 ),
    .o(\PWMC/n13 [19]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMC/mux0_b2  (
    .i0(\PWMC/n12 [2]),
    .i1(freqC[2]),
    .sel(\PWMC/n0 ),
    .o(\PWMC/n13 [2]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMC/mux0_b20  (
    .i0(\PWMC/n12 [20]),
    .i1(freqC[20]),
    .sel(\PWMC/n0 ),
    .o(\PWMC/n13 [20]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMC/mux0_b21  (
    .i0(\PWMC/n12 [21]),
    .i1(freqC[21]),
    .sel(\PWMC/n0 ),
    .o(\PWMC/n13 [21]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMC/mux0_b22  (
    .i0(\PWMC/n12 [22]),
    .i1(freqC[22]),
    .sel(\PWMC/n0 ),
    .o(\PWMC/n13 [22]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMC/mux0_b23  (
    .i0(\PWMC/n12 [23]),
    .i1(freqC[23]),
    .sel(\PWMC/n0 ),
    .o(\PWMC/n13 [23]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMC/mux0_b24  (
    .i0(\PWMC/n12 [24]),
    .i1(freqC[24]),
    .sel(\PWMC/n0 ),
    .o(\PWMC/n13 [24]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMC/mux0_b25  (
    .i0(\PWMC/n12 [25]),
    .i1(freqC[25]),
    .sel(\PWMC/n0 ),
    .o(\PWMC/n13 [25]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMC/mux0_b26  (
    .i0(\PWMC/n12 [26]),
    .i1(freqC[26]),
    .sel(\PWMC/n0 ),
    .o(\PWMC/n13 [26]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMC/mux0_b3  (
    .i0(\PWMC/n12 [3]),
    .i1(freqC[3]),
    .sel(\PWMC/n0 ),
    .o(\PWMC/n13 [3]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMC/mux0_b4  (
    .i0(\PWMC/n12 [4]),
    .i1(freqC[4]),
    .sel(\PWMC/n0 ),
    .o(\PWMC/n13 [4]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMC/mux0_b5  (
    .i0(\PWMC/n12 [5]),
    .i1(freqC[5]),
    .sel(\PWMC/n0 ),
    .o(\PWMC/n13 [5]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMC/mux0_b6  (
    .i0(\PWMC/n12 [6]),
    .i1(freqC[6]),
    .sel(\PWMC/n0 ),
    .o(\PWMC/n13 [6]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMC/mux0_b7  (
    .i0(\PWMC/n12 [7]),
    .i1(freqC[7]),
    .sel(\PWMC/n0 ),
    .o(\PWMC/n13 [7]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMC/mux0_b8  (
    .i0(\PWMC/n12 [8]),
    .i1(freqC[8]),
    .sel(\PWMC/n0 ),
    .o(\PWMC/n13 [8]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMC/mux0_b9  (
    .i0(\PWMC/n12 [9]),
    .i1(freqC[9]),
    .sel(\PWMC/n0 ),
    .o(\PWMC/n13 [9]));  // src/OnePWM.v(32)
  and \PWMC/mux3_b0_sel_is_3  (\PWMC/mux3_b0_sel_is_3_o , \PWMC/n11 , \PWMC/n0 );
  binary_mux_s1_w1 \PWMC/mux4_b0  (
    .i0(\PWMC/pnumr [0]),
    .i1(1'b0),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n22 [0]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux4_b1  (
    .i0(\PWMC/pnumr [1]),
    .i1(1'b0),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n22 [1]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux4_b10  (
    .i0(\PWMC/pnumr [10]),
    .i1(1'b0),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n22 [10]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux4_b11  (
    .i0(\PWMC/pnumr [11]),
    .i1(1'b0),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n22 [11]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux4_b12  (
    .i0(\PWMC/pnumr [12]),
    .i1(1'b0),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n22 [12]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux4_b13  (
    .i0(\PWMC/pnumr [13]),
    .i1(1'b0),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n22 [13]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux4_b14  (
    .i0(\PWMC/pnumr [14]),
    .i1(1'b0),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n22 [14]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux4_b15  (
    .i0(\PWMC/pnumr [15]),
    .i1(1'b0),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n22 [15]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux4_b16  (
    .i0(\PWMC/pnumr [16]),
    .i1(1'b0),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n22 [16]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux4_b17  (
    .i0(\PWMC/pnumr [17]),
    .i1(1'b0),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n22 [17]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux4_b18  (
    .i0(\PWMC/pnumr [18]),
    .i1(1'b0),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n22 [18]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux4_b19  (
    .i0(\PWMC/pnumr [19]),
    .i1(1'b0),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n22 [19]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux4_b2  (
    .i0(\PWMC/pnumr [2]),
    .i1(1'b0),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n22 [2]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux4_b20  (
    .i0(\PWMC/pnumr [20]),
    .i1(1'b0),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n22 [20]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux4_b21  (
    .i0(\PWMC/pnumr [21]),
    .i1(1'b0),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n22 [21]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux4_b22  (
    .i0(\PWMC/pnumr [22]),
    .i1(1'b0),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n22 [22]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux4_b23  (
    .i0(\PWMC/pnumr [23]),
    .i1(1'b0),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n22 [23]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux4_b24  (
    .i0(\PWMC/pnumr [24]),
    .i1(1'b0),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n22 [24]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux4_b25  (
    .i0(\PWMC/pnumr [25]),
    .i1(1'b0),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n22 [25]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux4_b26  (
    .i0(\PWMC/pnumr [26]),
    .i1(1'b0),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n22 [26]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux4_b27  (
    .i0(\PWMC/pnumr [27]),
    .i1(1'b0),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n22 [27]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux4_b28  (
    .i0(\PWMC/pnumr [28]),
    .i1(1'b0),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n22 [28]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux4_b29  (
    .i0(\PWMC/pnumr [29]),
    .i1(1'b0),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n22 [29]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux4_b3  (
    .i0(\PWMC/pnumr [3]),
    .i1(1'b0),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n22 [3]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux4_b30  (
    .i0(\PWMC/pnumr [30]),
    .i1(1'b0),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n22 [30]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux4_b31  (
    .i0(\PWMC/pnumr [31]),
    .i1(1'b0),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n22 [31]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux4_b4  (
    .i0(\PWMC/pnumr [4]),
    .i1(1'b0),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n22 [4]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux4_b5  (
    .i0(\PWMC/pnumr [5]),
    .i1(1'b0),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n22 [5]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux4_b6  (
    .i0(\PWMC/pnumr [6]),
    .i1(1'b0),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n22 [6]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux4_b7  (
    .i0(\PWMC/pnumr [7]),
    .i1(1'b0),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n22 [7]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux4_b8  (
    .i0(\PWMC/pnumr [8]),
    .i1(1'b0),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n22 [8]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux4_b9  (
    .i0(\PWMC/pnumr [9]),
    .i1(1'b0),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n22 [9]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux5_b0  (
    .i0(\PWMC/n22 [0]),
    .i1(pnumC[0]),
    .sel(pnumC[32]),
    .o(\PWMC/n23 [0]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux5_b1  (
    .i0(\PWMC/n22 [1]),
    .i1(pnumC[1]),
    .sel(pnumC[32]),
    .o(\PWMC/n23 [1]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux5_b10  (
    .i0(\PWMC/n22 [10]),
    .i1(pnumC[10]),
    .sel(pnumC[32]),
    .o(\PWMC/n23 [10]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux5_b11  (
    .i0(\PWMC/n22 [11]),
    .i1(pnumC[11]),
    .sel(pnumC[32]),
    .o(\PWMC/n23 [11]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux5_b12  (
    .i0(\PWMC/n22 [12]),
    .i1(pnumC[12]),
    .sel(pnumC[32]),
    .o(\PWMC/n23 [12]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux5_b13  (
    .i0(\PWMC/n22 [13]),
    .i1(pnumC[13]),
    .sel(pnumC[32]),
    .o(\PWMC/n23 [13]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux5_b14  (
    .i0(\PWMC/n22 [14]),
    .i1(pnumC[14]),
    .sel(pnumC[32]),
    .o(\PWMC/n23 [14]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux5_b15  (
    .i0(\PWMC/n22 [15]),
    .i1(pnumC[15]),
    .sel(pnumC[32]),
    .o(\PWMC/n23 [15]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux5_b16  (
    .i0(\PWMC/n22 [16]),
    .i1(pnumC[16]),
    .sel(pnumC[32]),
    .o(\PWMC/n23 [16]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux5_b17  (
    .i0(\PWMC/n22 [17]),
    .i1(pnumC[17]),
    .sel(pnumC[32]),
    .o(\PWMC/n23 [17]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux5_b18  (
    .i0(\PWMC/n22 [18]),
    .i1(pnumC[18]),
    .sel(pnumC[32]),
    .o(\PWMC/n23 [18]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux5_b19  (
    .i0(\PWMC/n22 [19]),
    .i1(pnumC[19]),
    .sel(pnumC[32]),
    .o(\PWMC/n23 [19]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux5_b2  (
    .i0(\PWMC/n22 [2]),
    .i1(pnumC[2]),
    .sel(pnumC[32]),
    .o(\PWMC/n23 [2]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux5_b20  (
    .i0(\PWMC/n22 [20]),
    .i1(pnumC[20]),
    .sel(pnumC[32]),
    .o(\PWMC/n23 [20]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux5_b21  (
    .i0(\PWMC/n22 [21]),
    .i1(pnumC[21]),
    .sel(pnumC[32]),
    .o(\PWMC/n23 [21]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux5_b22  (
    .i0(\PWMC/n22 [22]),
    .i1(pnumC[22]),
    .sel(pnumC[32]),
    .o(\PWMC/n23 [22]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux5_b23  (
    .i0(\PWMC/n22 [23]),
    .i1(pnumC[23]),
    .sel(pnumC[32]),
    .o(\PWMC/n23 [23]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux5_b24  (
    .i0(\PWMC/n22 [24]),
    .i1(pnumC[24]),
    .sel(pnumC[32]),
    .o(\PWMC/n23 [24]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux5_b25  (
    .i0(\PWMC/n22 [25]),
    .i1(pnumC[25]),
    .sel(pnumC[32]),
    .o(\PWMC/n23 [25]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux5_b26  (
    .i0(\PWMC/n22 [26]),
    .i1(pnumC[26]),
    .sel(pnumC[32]),
    .o(\PWMC/n23 [26]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux5_b27  (
    .i0(\PWMC/n22 [27]),
    .i1(pnumC[27]),
    .sel(pnumC[32]),
    .o(\PWMC/n23 [27]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux5_b28  (
    .i0(\PWMC/n22 [28]),
    .i1(pnumC[28]),
    .sel(pnumC[32]),
    .o(\PWMC/n23 [28]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux5_b29  (
    .i0(\PWMC/n22 [29]),
    .i1(pnumC[29]),
    .sel(pnumC[32]),
    .o(\PWMC/n23 [29]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux5_b3  (
    .i0(\PWMC/n22 [3]),
    .i1(pnumC[3]),
    .sel(pnumC[32]),
    .o(\PWMC/n23 [3]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux5_b30  (
    .i0(\PWMC/n22 [30]),
    .i1(pnumC[30]),
    .sel(pnumC[32]),
    .o(\PWMC/n23 [30]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux5_b31  (
    .i0(\PWMC/n22 [31]),
    .i1(pnumC[31]),
    .sel(pnumC[32]),
    .o(\PWMC/n23 [31]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux5_b4  (
    .i0(\PWMC/n22 [4]),
    .i1(pnumC[4]),
    .sel(pnumC[32]),
    .o(\PWMC/n23 [4]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux5_b5  (
    .i0(\PWMC/n22 [5]),
    .i1(pnumC[5]),
    .sel(pnumC[32]),
    .o(\PWMC/n23 [5]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux5_b6  (
    .i0(\PWMC/n22 [6]),
    .i1(pnumC[6]),
    .sel(pnumC[32]),
    .o(\PWMC/n23 [6]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux5_b7  (
    .i0(\PWMC/n22 [7]),
    .i1(pnumC[7]),
    .sel(pnumC[32]),
    .o(\PWMC/n23 [7]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux5_b8  (
    .i0(\PWMC/n22 [8]),
    .i1(pnumC[8]),
    .sel(pnumC[32]),
    .o(\PWMC/n23 [8]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux5_b9  (
    .i0(\PWMC/n22 [9]),
    .i1(pnumC[9]),
    .sel(pnumC[32]),
    .o(\PWMC/n23 [9]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMC/mux6_b0  (
    .i0(\PWMC/pnumr [0]),
    .i1(\PWMC/n26 [0]),
    .sel(\PWMC/n25 ),
    .o(\PWMC/n27 [0]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMC/mux6_b1  (
    .i0(\PWMC/pnumr [1]),
    .i1(\PWMC/n26 [1]),
    .sel(\PWMC/n25 ),
    .o(\PWMC/n27 [1]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMC/mux6_b10  (
    .i0(\PWMC/pnumr [10]),
    .i1(\PWMC/n26 [10]),
    .sel(\PWMC/n25 ),
    .o(\PWMC/n27 [10]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMC/mux6_b11  (
    .i0(\PWMC/pnumr [11]),
    .i1(\PWMC/n26 [11]),
    .sel(\PWMC/n25 ),
    .o(\PWMC/n27 [11]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMC/mux6_b12  (
    .i0(\PWMC/pnumr [12]),
    .i1(\PWMC/n26 [12]),
    .sel(\PWMC/n25 ),
    .o(\PWMC/n27 [12]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMC/mux6_b13  (
    .i0(\PWMC/pnumr [13]),
    .i1(\PWMC/n26 [13]),
    .sel(\PWMC/n25 ),
    .o(\PWMC/n27 [13]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMC/mux6_b14  (
    .i0(\PWMC/pnumr [14]),
    .i1(\PWMC/n26 [14]),
    .sel(\PWMC/n25 ),
    .o(\PWMC/n27 [14]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMC/mux6_b15  (
    .i0(\PWMC/pnumr [15]),
    .i1(\PWMC/n26 [15]),
    .sel(\PWMC/n25 ),
    .o(\PWMC/n27 [15]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMC/mux6_b16  (
    .i0(\PWMC/pnumr [16]),
    .i1(\PWMC/n26 [16]),
    .sel(\PWMC/n25 ),
    .o(\PWMC/n27 [16]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMC/mux6_b17  (
    .i0(\PWMC/pnumr [17]),
    .i1(\PWMC/n26 [17]),
    .sel(\PWMC/n25 ),
    .o(\PWMC/n27 [17]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMC/mux6_b18  (
    .i0(\PWMC/pnumr [18]),
    .i1(\PWMC/n26 [18]),
    .sel(\PWMC/n25 ),
    .o(\PWMC/n27 [18]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMC/mux6_b19  (
    .i0(\PWMC/pnumr [19]),
    .i1(\PWMC/n26 [19]),
    .sel(\PWMC/n25 ),
    .o(\PWMC/n27 [19]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMC/mux6_b2  (
    .i0(\PWMC/pnumr [2]),
    .i1(\PWMC/n26 [2]),
    .sel(\PWMC/n25 ),
    .o(\PWMC/n27 [2]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMC/mux6_b20  (
    .i0(\PWMC/pnumr [20]),
    .i1(\PWMC/n26 [20]),
    .sel(\PWMC/n25 ),
    .o(\PWMC/n27 [20]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMC/mux6_b21  (
    .i0(\PWMC/pnumr [21]),
    .i1(\PWMC/n26 [21]),
    .sel(\PWMC/n25 ),
    .o(\PWMC/n27 [21]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMC/mux6_b22  (
    .i0(\PWMC/pnumr [22]),
    .i1(\PWMC/n26 [22]),
    .sel(\PWMC/n25 ),
    .o(\PWMC/n27 [22]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMC/mux6_b23  (
    .i0(\PWMC/pnumr [23]),
    .i1(\PWMC/n26 [23]),
    .sel(\PWMC/n25 ),
    .o(\PWMC/n27 [23]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMC/mux6_b3  (
    .i0(\PWMC/pnumr [3]),
    .i1(\PWMC/n26 [3]),
    .sel(\PWMC/n25 ),
    .o(\PWMC/n27 [3]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMC/mux6_b4  (
    .i0(\PWMC/pnumr [4]),
    .i1(\PWMC/n26 [4]),
    .sel(\PWMC/n25 ),
    .o(\PWMC/n27 [4]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMC/mux6_b5  (
    .i0(\PWMC/pnumr [5]),
    .i1(\PWMC/n26 [5]),
    .sel(\PWMC/n25 ),
    .o(\PWMC/n27 [5]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMC/mux6_b6  (
    .i0(\PWMC/pnumr [6]),
    .i1(\PWMC/n26 [6]),
    .sel(\PWMC/n25 ),
    .o(\PWMC/n27 [6]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMC/mux6_b7  (
    .i0(\PWMC/pnumr [7]),
    .i1(\PWMC/n26 [7]),
    .sel(\PWMC/n25 ),
    .o(\PWMC/n27 [7]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMC/mux6_b8  (
    .i0(\PWMC/pnumr [8]),
    .i1(\PWMC/n26 [8]),
    .sel(\PWMC/n25 ),
    .o(\PWMC/n27 [8]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMC/mux6_b9  (
    .i0(\PWMC/pnumr [9]),
    .i1(\PWMC/n26 [9]),
    .sel(\PWMC/n25 ),
    .o(\PWMC/n27 [9]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMC/mux7_b0  (
    .i0(pnumcntC[0]),
    .i1(\PWMC/n27 [0]),
    .sel(\PWMC/n24 ),
    .o(\PWMC/n29 [0]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux7_b1  (
    .i0(pnumcntC[1]),
    .i1(\PWMC/n27 [1]),
    .sel(\PWMC/n24 ),
    .o(\PWMC/n29 [1]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux7_b10  (
    .i0(pnumcntC[10]),
    .i1(\PWMC/n27 [10]),
    .sel(\PWMC/n24 ),
    .o(\PWMC/n29 [10]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux7_b11  (
    .i0(pnumcntC[11]),
    .i1(\PWMC/n27 [11]),
    .sel(\PWMC/n24 ),
    .o(\PWMC/n29 [11]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux7_b12  (
    .i0(pnumcntC[12]),
    .i1(\PWMC/n27 [12]),
    .sel(\PWMC/n24 ),
    .o(\PWMC/n29 [12]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux7_b13  (
    .i0(pnumcntC[13]),
    .i1(\PWMC/n27 [13]),
    .sel(\PWMC/n24 ),
    .o(\PWMC/n29 [13]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux7_b14  (
    .i0(pnumcntC[14]),
    .i1(\PWMC/n27 [14]),
    .sel(\PWMC/n24 ),
    .o(\PWMC/n29 [14]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux7_b15  (
    .i0(pnumcntC[15]),
    .i1(\PWMC/n27 [15]),
    .sel(\PWMC/n24 ),
    .o(\PWMC/n29 [15]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux7_b16  (
    .i0(pnumcntC[16]),
    .i1(\PWMC/n27 [16]),
    .sel(\PWMC/n24 ),
    .o(\PWMC/n29 [16]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux7_b17  (
    .i0(pnumcntC[17]),
    .i1(\PWMC/n27 [17]),
    .sel(\PWMC/n24 ),
    .o(\PWMC/n29 [17]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux7_b18  (
    .i0(pnumcntC[18]),
    .i1(\PWMC/n27 [18]),
    .sel(\PWMC/n24 ),
    .o(\PWMC/n29 [18]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux7_b19  (
    .i0(pnumcntC[19]),
    .i1(\PWMC/n27 [19]),
    .sel(\PWMC/n24 ),
    .o(\PWMC/n29 [19]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux7_b2  (
    .i0(pnumcntC[2]),
    .i1(\PWMC/n27 [2]),
    .sel(\PWMC/n24 ),
    .o(\PWMC/n29 [2]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux7_b20  (
    .i0(pnumcntC[20]),
    .i1(\PWMC/n27 [20]),
    .sel(\PWMC/n24 ),
    .o(\PWMC/n29 [20]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux7_b21  (
    .i0(pnumcntC[21]),
    .i1(\PWMC/n27 [21]),
    .sel(\PWMC/n24 ),
    .o(\PWMC/n29 [21]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux7_b22  (
    .i0(pnumcntC[22]),
    .i1(\PWMC/n27 [22]),
    .sel(\PWMC/n24 ),
    .o(\PWMC/n29 [22]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux7_b23  (
    .i0(pnumcntC[23]),
    .i1(\PWMC/n27 [23]),
    .sel(\PWMC/n24 ),
    .o(\PWMC/n29 [23]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux7_b3  (
    .i0(pnumcntC[3]),
    .i1(\PWMC/n27 [3]),
    .sel(\PWMC/n24 ),
    .o(\PWMC/n29 [3]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux7_b4  (
    .i0(pnumcntC[4]),
    .i1(\PWMC/n27 [4]),
    .sel(\PWMC/n24 ),
    .o(\PWMC/n29 [4]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux7_b5  (
    .i0(pnumcntC[5]),
    .i1(\PWMC/n27 [5]),
    .sel(\PWMC/n24 ),
    .o(\PWMC/n29 [5]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux7_b6  (
    .i0(pnumcntC[6]),
    .i1(\PWMC/n27 [6]),
    .sel(\PWMC/n24 ),
    .o(\PWMC/n29 [6]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux7_b7  (
    .i0(pnumcntC[7]),
    .i1(\PWMC/n27 [7]),
    .sel(\PWMC/n24 ),
    .o(\PWMC/n29 [7]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux7_b8  (
    .i0(pnumcntC[8]),
    .i1(\PWMC/n27 [8]),
    .sel(\PWMC/n24 ),
    .o(\PWMC/n29 [8]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux7_b9  (
    .i0(pnumcntC[9]),
    .i1(\PWMC/n27 [9]),
    .sel(\PWMC/n24 ),
    .o(\PWMC/n29 [9]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux8_b0  (
    .i0(\PWMC/n29 [0]),
    .i1(\PWMC/pnumr [0]),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n31 [0]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux8_b1  (
    .i0(\PWMC/n29 [1]),
    .i1(\PWMC/pnumr [1]),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n31 [1]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux8_b10  (
    .i0(\PWMC/n29 [10]),
    .i1(\PWMC/pnumr [10]),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n31 [10]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux8_b11  (
    .i0(\PWMC/n29 [11]),
    .i1(\PWMC/pnumr [11]),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n31 [11]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux8_b12  (
    .i0(\PWMC/n29 [12]),
    .i1(\PWMC/pnumr [12]),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n31 [12]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux8_b13  (
    .i0(\PWMC/n29 [13]),
    .i1(\PWMC/pnumr [13]),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n31 [13]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux8_b14  (
    .i0(\PWMC/n29 [14]),
    .i1(\PWMC/pnumr [14]),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n31 [14]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux8_b15  (
    .i0(\PWMC/n29 [15]),
    .i1(\PWMC/pnumr [15]),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n31 [15]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux8_b16  (
    .i0(\PWMC/n29 [16]),
    .i1(\PWMC/pnumr [16]),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n31 [16]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux8_b17  (
    .i0(\PWMC/n29 [17]),
    .i1(\PWMC/pnumr [17]),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n31 [17]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux8_b18  (
    .i0(\PWMC/n29 [18]),
    .i1(\PWMC/pnumr [18]),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n31 [18]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux8_b19  (
    .i0(\PWMC/n29 [19]),
    .i1(\PWMC/pnumr [19]),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n31 [19]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux8_b2  (
    .i0(\PWMC/n29 [2]),
    .i1(\PWMC/pnumr [2]),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n31 [2]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux8_b20  (
    .i0(\PWMC/n29 [20]),
    .i1(\PWMC/pnumr [20]),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n31 [20]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux8_b21  (
    .i0(\PWMC/n29 [21]),
    .i1(\PWMC/pnumr [21]),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n31 [21]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux8_b22  (
    .i0(\PWMC/n29 [22]),
    .i1(\PWMC/pnumr [22]),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n31 [22]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux8_b23  (
    .i0(\PWMC/n29 [23]),
    .i1(\PWMC/pnumr [23]),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n31 [23]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux8_b3  (
    .i0(\PWMC/n29 [3]),
    .i1(\PWMC/pnumr [3]),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n31 [3]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux8_b4  (
    .i0(\PWMC/n29 [4]),
    .i1(\PWMC/pnumr [4]),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n31 [4]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux8_b5  (
    .i0(\PWMC/n29 [5]),
    .i1(\PWMC/pnumr [5]),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n31 [5]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux8_b6  (
    .i0(\PWMC/n29 [6]),
    .i1(\PWMC/pnumr [6]),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n31 [6]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux8_b7  (
    .i0(\PWMC/n29 [7]),
    .i1(\PWMC/pnumr [7]),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n31 [7]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux8_b8  (
    .i0(\PWMC/n29 [8]),
    .i1(\PWMC/pnumr [8]),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n31 [8]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMC/mux8_b9  (
    .i0(\PWMC/n29 [9]),
    .i1(\PWMC/pnumr [9]),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n31 [9]));  // src/OnePWM.v(57)
  not \PWMC/n17_inv  (\PWMC/n17_neg , \PWMC/n17 );
  not \PWMC/n25_inv  (\PWMC/n25_neg , \PWMC/n25 );
  not \PWMC/n4_inv  (\PWMC/n4_neg , \PWMC/n4 );
  not \PWMC/n6_inv  (\PWMC/n6_neg , \PWMC/n6 );
  ne_w24 \PWMC/neq0  (
    .i0(pnumcntC),
    .i1(24'b000000000000000000000000),
    .o(\PWMC/n25 ));  // src/OnePWM.v(55)
  reg_sr_ss_w1 \PWMC/pwm_reg  (
    .clk(clk100m),
    .d(pwm[12]),
    .en(1'b1),
    .reset(~\PWMC/u14_sel_is_1_o ),
    .set(\PWMC/n18 ),
    .q(\PWMC/pwm_keep ));  // src/OnePWM.v(45)
  reg_sr_as_w1 \PWMC/reg0_b0  (
    .clk(clk100m),
    .d(\PWMC/n13 [0]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [0]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b1  (
    .clk(clk100m),
    .d(\PWMC/n13 [1]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [1]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b10  (
    .clk(clk100m),
    .d(\PWMC/n13 [10]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [10]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b11  (
    .clk(clk100m),
    .d(\PWMC/n13 [11]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [11]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b12  (
    .clk(clk100m),
    .d(\PWMC/n13 [12]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [12]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b13  (
    .clk(clk100m),
    .d(\PWMC/n13 [13]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [13]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b14  (
    .clk(clk100m),
    .d(\PWMC/n13 [14]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [14]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b15  (
    .clk(clk100m),
    .d(\PWMC/n13 [15]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [15]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b16  (
    .clk(clk100m),
    .d(\PWMC/n13 [16]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [16]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b17  (
    .clk(clk100m),
    .d(\PWMC/n13 [17]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [17]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b18  (
    .clk(clk100m),
    .d(\PWMC/n13 [18]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [18]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b19  (
    .clk(clk100m),
    .d(\PWMC/n13 [19]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [19]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b2  (
    .clk(clk100m),
    .d(\PWMC/n13 [2]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [2]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b20  (
    .clk(clk100m),
    .d(\PWMC/n13 [20]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [20]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b21  (
    .clk(clk100m),
    .d(\PWMC/n13 [21]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [21]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b22  (
    .clk(clk100m),
    .d(\PWMC/n13 [22]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [22]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b23  (
    .clk(clk100m),
    .d(\PWMC/n13 [23]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [23]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b24  (
    .clk(clk100m),
    .d(\PWMC/n13 [24]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [24]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b25  (
    .clk(clk100m),
    .d(\PWMC/n13 [25]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [25]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b26  (
    .clk(clk100m),
    .d(\PWMC/n13 [26]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [26]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b3  (
    .clk(clk100m),
    .d(\PWMC/n13 [3]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [3]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b4  (
    .clk(clk100m),
    .d(\PWMC/n13 [4]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [4]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b5  (
    .clk(clk100m),
    .d(\PWMC/n13 [5]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [5]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b6  (
    .clk(clk100m),
    .d(\PWMC/n13 [6]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [6]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b7  (
    .clk(clk100m),
    .d(\PWMC/n13 [7]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [7]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b8  (
    .clk(clk100m),
    .d(\PWMC/n13 [8]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [8]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMC/reg0_b9  (
    .clk(clk100m),
    .d(\PWMC/n13 [9]),
    .en(1'b1),
    .reset(~\PWMC/n11 ),
    .set(1'b0),
    .q(\PWMC/FreCnt [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b0  (
    .clk(clk100m),
    .d(freqC[0]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [0]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b1  (
    .clk(clk100m),
    .d(freqC[1]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [1]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b10  (
    .clk(clk100m),
    .d(freqC[10]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [10]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b11  (
    .clk(clk100m),
    .d(freqC[11]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [11]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b12  (
    .clk(clk100m),
    .d(freqC[12]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [12]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b13  (
    .clk(clk100m),
    .d(freqC[13]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [13]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b14  (
    .clk(clk100m),
    .d(freqC[14]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [14]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b15  (
    .clk(clk100m),
    .d(freqC[15]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [15]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b16  (
    .clk(clk100m),
    .d(freqC[16]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [16]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b17  (
    .clk(clk100m),
    .d(freqC[17]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [17]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b18  (
    .clk(clk100m),
    .d(freqC[18]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [18]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b19  (
    .clk(clk100m),
    .d(freqC[19]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [19]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b2  (
    .clk(clk100m),
    .d(freqC[2]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [2]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b20  (
    .clk(clk100m),
    .d(freqC[20]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [20]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b21  (
    .clk(clk100m),
    .d(freqC[21]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [21]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b22  (
    .clk(clk100m),
    .d(freqC[22]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [22]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b23  (
    .clk(clk100m),
    .d(freqC[23]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [23]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b24  (
    .clk(clk100m),
    .d(freqC[24]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [24]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b25  (
    .clk(clk100m),
    .d(freqC[25]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [25]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b26  (
    .clk(clk100m),
    .d(freqC[26]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [26]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b3  (
    .clk(clk100m),
    .d(freqC[3]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [3]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b4  (
    .clk(clk100m),
    .d(freqC[4]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [4]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b5  (
    .clk(clk100m),
    .d(freqC[5]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [5]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b6  (
    .clk(clk100m),
    .d(freqC[6]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [6]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b7  (
    .clk(clk100m),
    .d(freqC[7]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [7]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b8  (
    .clk(clk100m),
    .d(freqC[8]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [8]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg1_b9  (
    .clk(clk100m),
    .d(freqC[9]),
    .en(\PWMC/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/FreCntr [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMC/reg2_b0  (
    .clk(clk100m),
    .d(\PWMC/n23 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[0]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b1  (
    .clk(clk100m),
    .d(\PWMC/n23 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[1]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b10  (
    .clk(clk100m),
    .d(\PWMC/n23 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[10]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b11  (
    .clk(clk100m),
    .d(\PWMC/n23 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[11]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b12  (
    .clk(clk100m),
    .d(\PWMC/n23 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[12]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b13  (
    .clk(clk100m),
    .d(\PWMC/n23 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[13]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b14  (
    .clk(clk100m),
    .d(\PWMC/n23 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[14]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b15  (
    .clk(clk100m),
    .d(\PWMC/n23 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[15]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b16  (
    .clk(clk100m),
    .d(\PWMC/n23 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[16]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b17  (
    .clk(clk100m),
    .d(\PWMC/n23 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[17]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b18  (
    .clk(clk100m),
    .d(\PWMC/n23 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[18]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b19  (
    .clk(clk100m),
    .d(\PWMC/n23 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[19]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b2  (
    .clk(clk100m),
    .d(\PWMC/n23 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[2]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b20  (
    .clk(clk100m),
    .d(\PWMC/n23 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[20]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b21  (
    .clk(clk100m),
    .d(\PWMC/n23 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[21]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b22  (
    .clk(clk100m),
    .d(\PWMC/n23 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[22]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b23  (
    .clk(clk100m),
    .d(\PWMC/n23 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[23]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b24  (
    .clk(clk100m),
    .d(\PWMC/n23 [24]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[24]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b25  (
    .clk(clk100m),
    .d(\PWMC/n23 [25]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[25]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b26  (
    .clk(clk100m),
    .d(\PWMC/n23 [26]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[26]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b27  (
    .clk(clk100m),
    .d(\PWMC/n23 [27]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[27]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b28  (
    .clk(clk100m),
    .d(\PWMC/n23 [28]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[28]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b29  (
    .clk(clk100m),
    .d(\PWMC/n23 [29]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[29]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b3  (
    .clk(clk100m),
    .d(\PWMC/n23 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[3]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b30  (
    .clk(clk100m),
    .d(\PWMC/n23 [30]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[30]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b31  (
    .clk(clk100m),
    .d(\PWMC/n23 [31]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[31]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b4  (
    .clk(clk100m),
    .d(\PWMC/n23 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[4]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b5  (
    .clk(clk100m),
    .d(\PWMC/n23 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[5]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b6  (
    .clk(clk100m),
    .d(\PWMC/n23 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[6]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b7  (
    .clk(clk100m),
    .d(\PWMC/n23 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[7]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b8  (
    .clk(clk100m),
    .d(\PWMC/n23 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[8]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg2_b9  (
    .clk(clk100m),
    .d(\PWMC/n23 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/pnumr[9]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMC/reg3_b0  (
    .clk(clk100m),
    .d(\PWMC/n31 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[0]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b1  (
    .clk(clk100m),
    .d(\PWMC/n31 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[1]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b10  (
    .clk(clk100m),
    .d(\PWMC/n31 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[10]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b11  (
    .clk(clk100m),
    .d(\PWMC/n31 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[11]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b12  (
    .clk(clk100m),
    .d(\PWMC/n31 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[12]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b13  (
    .clk(clk100m),
    .d(\PWMC/n31 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[13]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b14  (
    .clk(clk100m),
    .d(\PWMC/n31 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[14]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b15  (
    .clk(clk100m),
    .d(\PWMC/n31 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[15]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b16  (
    .clk(clk100m),
    .d(\PWMC/n31 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[16]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b17  (
    .clk(clk100m),
    .d(\PWMC/n31 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[17]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b18  (
    .clk(clk100m),
    .d(\PWMC/n31 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[18]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b19  (
    .clk(clk100m),
    .d(\PWMC/n31 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[19]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b2  (
    .clk(clk100m),
    .d(\PWMC/n31 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[2]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b20  (
    .clk(clk100m),
    .d(\PWMC/n31 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[20]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b21  (
    .clk(clk100m),
    .d(\PWMC/n31 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[21]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b22  (
    .clk(clk100m),
    .d(\PWMC/n31 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[22]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b23  (
    .clk(clk100m),
    .d(\PWMC/n31 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[23]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b3  (
    .clk(clk100m),
    .d(\PWMC/n31 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[3]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b4  (
    .clk(clk100m),
    .d(\PWMC/n31 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[4]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b5  (
    .clk(clk100m),
    .d(\PWMC/n31 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[5]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b6  (
    .clk(clk100m),
    .d(\PWMC/n31 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[6]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b7  (
    .clk(clk100m),
    .d(\PWMC/n31 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[7]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b8  (
    .clk(clk100m),
    .d(\PWMC/n31 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[8]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMC/reg3_b9  (
    .clk(clk100m),
    .d(\PWMC/n31 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMC/RemaTxNum[9]_keep ));  // src/OnePWM.v(58)
  reg_ar_ss_w1 \PWMC/stopreq_reg  (
    .clk(clk100m),
    .d(\PWMC/n1 ),
    .en(1'b1),
    .reset(1'b0),
    .set(pwm_start_stop[12]),
    .q(\PWMC/stopreq_keep ));  // src/OnePWM.v(15)
  add_pu27_mu27_o27 \PWMC/sub0  (
    .i0(\PWMC/FreCnt ),
    .i1(27'b000000000000000000000000001),
    .o(\PWMC/n12 [26:0]));  // src/OnePWM.v(32)
  add_pu24_mu24_o24 \PWMC/sub1  (
    .i0(pnumcntC),
    .i1(24'b000000000000000000000001),
    .o(\PWMC/n26 [23:0]));  // src/OnePWM.v(55)
  AL_MUX \PWMC/u10  (
    .i0(1'b0),
    .i1(\PWMC/n9 ),
    .sel(n23),
    .o(\PWMC/n10 ));  // src/OnePWM.v(26)
  or \PWMC/u11  (\PWMC/n11 , pwm_state_read[12], pwm_start_stop[28]);  // src/OnePWM.v(30)
  and \PWMC/u14_sel_is_1  (\PWMC/u14_sel_is_1_o , pwm_state_read[12], \PWMC/n17_neg );
  and \PWMC/u15  (\PWMC/n24 , \PWMC/n0 , pwm_state_read[12]);  // src/OnePWM.v(54)
  and \PWMC/u17_sel_is_1  (\PWMC/u17_sel_is_1_o , \PWMC/n24 , \PWMC/n25_neg );
  not \PWMC/u17_sel_is_1_o_inv  (\PWMC/u17_sel_is_1_o_neg , \PWMC/u17_sel_is_1_o );
  AL_MUX \PWMC/u18  (
    .i0(\PWMC/pnumr [31]),
    .i1(dir[12]),
    .sel(\PWMC/u18_sel_is_0_o ),
    .o(\PWMC/n32 ));
  and \PWMC/u18_sel_is_0  (\PWMC/u18_sel_is_0_o , \pwm_start_stop[28]_neg , \PWMC/u17_sel_is_1_o_neg );
  AL_MUX \PWMC/u2  (
    .i0(\PWMC/stopreq ),
    .i1(1'b0),
    .sel(\PWMC/n0 ),
    .o(\PWMC/n1 ));  // src/OnePWM.v(15)
  and \PWMC/u5  (\PWMC/n4 , \PWMC/stopreq , \PWMC/n0 );  // src/OnePWM.v(23)
  and \PWMC/u6  (\PWMC/n6 , \PWMC/n5 , \PWMC/n0 );  // src/OnePWM.v(25)
  AL_MUX \PWMC/u8  (
    .i0(1'b0),
    .i1(pwm_state_read[12]),
    .sel(\PWMC/u8_sel_is_0_o ),
    .o(\PWMC/n8 ));
  and \PWMC/u8_sel_is_0  (\PWMC/u8_sel_is_0_o , \PWMC/n4_neg , \PWMC/n6_neg );
  AL_MUX \PWMC/u9  (
    .i0(\PWMC/n8 ),
    .i1(1'b1),
    .sel(pwm_start_stop[28]),
    .o(\PWMC/n9 ));  // src/OnePWM.v(26)
  reg_ar_as_w1 \PWMD/State_reg  (
    .clk(clk100m),
    .d(\PWMD/n10 ),
    .en(1'b1),
    .reset(~rstn),
    .set(1'b0),
    .q(pwm_state_read[13]));  // src/OnePWM.v(26)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[0]  (
    .i(\PWMD/RemaTxNum[0]_keep ),
    .o(pnumcntD[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[10]  (
    .i(\PWMD/RemaTxNum[10]_keep ),
    .o(pnumcntD[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[11]  (
    .i(\PWMD/RemaTxNum[11]_keep ),
    .o(pnumcntD[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[12]  (
    .i(\PWMD/RemaTxNum[12]_keep ),
    .o(pnumcntD[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[13]  (
    .i(\PWMD/RemaTxNum[13]_keep ),
    .o(pnumcntD[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[14]  (
    .i(\PWMD/RemaTxNum[14]_keep ),
    .o(pnumcntD[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[15]  (
    .i(\PWMD/RemaTxNum[15]_keep ),
    .o(pnumcntD[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[16]  (
    .i(\PWMD/RemaTxNum[16]_keep ),
    .o(pnumcntD[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[17]  (
    .i(\PWMD/RemaTxNum[17]_keep ),
    .o(pnumcntD[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[18]  (
    .i(\PWMD/RemaTxNum[18]_keep ),
    .o(pnumcntD[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[19]  (
    .i(\PWMD/RemaTxNum[19]_keep ),
    .o(pnumcntD[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[1]  (
    .i(\PWMD/RemaTxNum[1]_keep ),
    .o(pnumcntD[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[20]  (
    .i(\PWMD/RemaTxNum[20]_keep ),
    .o(pnumcntD[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[21]  (
    .i(\PWMD/RemaTxNum[21]_keep ),
    .o(pnumcntD[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[22]  (
    .i(\PWMD/RemaTxNum[22]_keep ),
    .o(pnumcntD[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[23]  (
    .i(\PWMD/RemaTxNum[23]_keep ),
    .o(pnumcntD[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[2]  (
    .i(\PWMD/RemaTxNum[2]_keep ),
    .o(pnumcntD[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[3]  (
    .i(\PWMD/RemaTxNum[3]_keep ),
    .o(pnumcntD[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[4]  (
    .i(\PWMD/RemaTxNum[4]_keep ),
    .o(pnumcntD[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[5]  (
    .i(\PWMD/RemaTxNum[5]_keep ),
    .o(pnumcntD[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[6]  (
    .i(\PWMD/RemaTxNum[6]_keep ),
    .o(pnumcntD[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[7]  (
    .i(\PWMD/RemaTxNum[7]_keep ),
    .o(pnumcntD[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[8]  (
    .i(\PWMD/RemaTxNum[8]_keep ),
    .o(pnumcntD[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_RemaTxNum[9]  (
    .i(\PWMD/RemaTxNum[9]_keep ),
    .o(pnumcntD[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_dir  (
    .i(\PWMD/dir_keep ),
    .o(dir[13]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[0]  (
    .i(\PWMD/pnumr[0]_keep ),
    .o(\PWMD/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[10]  (
    .i(\PWMD/pnumr[10]_keep ),
    .o(\PWMD/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[11]  (
    .i(\PWMD/pnumr[11]_keep ),
    .o(\PWMD/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[12]  (
    .i(\PWMD/pnumr[12]_keep ),
    .o(\PWMD/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[13]  (
    .i(\PWMD/pnumr[13]_keep ),
    .o(\PWMD/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[14]  (
    .i(\PWMD/pnumr[14]_keep ),
    .o(\PWMD/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[15]  (
    .i(\PWMD/pnumr[15]_keep ),
    .o(\PWMD/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[16]  (
    .i(\PWMD/pnumr[16]_keep ),
    .o(\PWMD/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[17]  (
    .i(\PWMD/pnumr[17]_keep ),
    .o(\PWMD/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[18]  (
    .i(\PWMD/pnumr[18]_keep ),
    .o(\PWMD/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[19]  (
    .i(\PWMD/pnumr[19]_keep ),
    .o(\PWMD/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[1]  (
    .i(\PWMD/pnumr[1]_keep ),
    .o(\PWMD/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[20]  (
    .i(\PWMD/pnumr[20]_keep ),
    .o(\PWMD/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[21]  (
    .i(\PWMD/pnumr[21]_keep ),
    .o(\PWMD/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[22]  (
    .i(\PWMD/pnumr[22]_keep ),
    .o(\PWMD/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[23]  (
    .i(\PWMD/pnumr[23]_keep ),
    .o(\PWMD/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[24]  (
    .i(\PWMD/pnumr[24]_keep ),
    .o(\PWMD/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[25]  (
    .i(\PWMD/pnumr[25]_keep ),
    .o(\PWMD/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[26]  (
    .i(\PWMD/pnumr[26]_keep ),
    .o(\PWMD/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[27]  (
    .i(\PWMD/pnumr[27]_keep ),
    .o(\PWMD/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[28]  (
    .i(\PWMD/pnumr[28]_keep ),
    .o(\PWMD/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[29]  (
    .i(\PWMD/pnumr[29]_keep ),
    .o(\PWMD/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[2]  (
    .i(\PWMD/pnumr[2]_keep ),
    .o(\PWMD/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[30]  (
    .i(\PWMD/pnumr[30]_keep ),
    .o(\PWMD/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[31]  (
    .i(\PWMD/pnumr[31]_keep ),
    .o(\PWMD/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[3]  (
    .i(\PWMD/pnumr[3]_keep ),
    .o(\PWMD/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[4]  (
    .i(\PWMD/pnumr[4]_keep ),
    .o(\PWMD/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[5]  (
    .i(\PWMD/pnumr[5]_keep ),
    .o(\PWMD/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[6]  (
    .i(\PWMD/pnumr[6]_keep ),
    .o(\PWMD/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[7]  (
    .i(\PWMD/pnumr[7]_keep ),
    .o(\PWMD/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[8]  (
    .i(\PWMD/pnumr[8]_keep ),
    .o(\PWMD/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pnumr[9]  (
    .i(\PWMD/pnumr[9]_keep ),
    .o(\PWMD/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_pwm  (
    .i(\PWMD/pwm_keep ),
    .o(pwm[13]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMD/_bufkeep_stopreq  (
    .i(\PWMD/stopreq_keep ),
    .o(\PWMD/stopreq ));  // src/OnePWM.v(14)
  reg_ar_as_w1 \PWMD/dir_reg  (
    .clk(clk100m),
    .d(\PWMD/n32 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/dir_keep ));  // src/OnePWM.v(58)
  eq_w27 \PWMD/eq0  (
    .i0(\PWMD/FreCnt ),
    .i1(27'b000000000000000000000000000),
    .o(\PWMD/n0 ));  // src/OnePWM.v(15)
  eq_w24 \PWMD/eq1  (
    .i0(pnumcntD),
    .i1(24'b000000000000000000000001),
    .o(\PWMD/n5 ));  // src/OnePWM.v(25)
  eq_w27 \PWMD/eq2  (
    .i0(\PWMD/FreCnt ),
    .i1({1'b0,\PWMD/FreCntr [26:1]}),
    .o(\PWMD/n17 ));  // src/OnePWM.v(41)
  eq_w27 \PWMD/eq3  (
    .i0(\PWMD/FreCnt ),
    .i1(\PWMD/FreCntr ),
    .o(\PWMD/n18 ));  // src/OnePWM.v(43)
  binary_mux_s1_w1 \PWMD/mux0_b0  (
    .i0(\PWMD/n12 [0]),
    .i1(freqD[0]),
    .sel(\PWMD/n0 ),
    .o(\PWMD/n13 [0]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMD/mux0_b1  (
    .i0(\PWMD/n12 [1]),
    .i1(freqD[1]),
    .sel(\PWMD/n0 ),
    .o(\PWMD/n13 [1]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMD/mux0_b10  (
    .i0(\PWMD/n12 [10]),
    .i1(freqD[10]),
    .sel(\PWMD/n0 ),
    .o(\PWMD/n13 [10]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMD/mux0_b11  (
    .i0(\PWMD/n12 [11]),
    .i1(freqD[11]),
    .sel(\PWMD/n0 ),
    .o(\PWMD/n13 [11]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMD/mux0_b12  (
    .i0(\PWMD/n12 [12]),
    .i1(freqD[12]),
    .sel(\PWMD/n0 ),
    .o(\PWMD/n13 [12]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMD/mux0_b13  (
    .i0(\PWMD/n12 [13]),
    .i1(freqD[13]),
    .sel(\PWMD/n0 ),
    .o(\PWMD/n13 [13]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMD/mux0_b14  (
    .i0(\PWMD/n12 [14]),
    .i1(freqD[14]),
    .sel(\PWMD/n0 ),
    .o(\PWMD/n13 [14]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMD/mux0_b15  (
    .i0(\PWMD/n12 [15]),
    .i1(freqD[15]),
    .sel(\PWMD/n0 ),
    .o(\PWMD/n13 [15]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMD/mux0_b16  (
    .i0(\PWMD/n12 [16]),
    .i1(freqD[16]),
    .sel(\PWMD/n0 ),
    .o(\PWMD/n13 [16]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMD/mux0_b17  (
    .i0(\PWMD/n12 [17]),
    .i1(freqD[17]),
    .sel(\PWMD/n0 ),
    .o(\PWMD/n13 [17]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMD/mux0_b18  (
    .i0(\PWMD/n12 [18]),
    .i1(freqD[18]),
    .sel(\PWMD/n0 ),
    .o(\PWMD/n13 [18]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMD/mux0_b19  (
    .i0(\PWMD/n12 [19]),
    .i1(freqD[19]),
    .sel(\PWMD/n0 ),
    .o(\PWMD/n13 [19]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMD/mux0_b2  (
    .i0(\PWMD/n12 [2]),
    .i1(freqD[2]),
    .sel(\PWMD/n0 ),
    .o(\PWMD/n13 [2]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMD/mux0_b20  (
    .i0(\PWMD/n12 [20]),
    .i1(freqD[20]),
    .sel(\PWMD/n0 ),
    .o(\PWMD/n13 [20]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMD/mux0_b21  (
    .i0(\PWMD/n12 [21]),
    .i1(freqD[21]),
    .sel(\PWMD/n0 ),
    .o(\PWMD/n13 [21]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMD/mux0_b22  (
    .i0(\PWMD/n12 [22]),
    .i1(freqD[22]),
    .sel(\PWMD/n0 ),
    .o(\PWMD/n13 [22]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMD/mux0_b23  (
    .i0(\PWMD/n12 [23]),
    .i1(freqD[23]),
    .sel(\PWMD/n0 ),
    .o(\PWMD/n13 [23]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMD/mux0_b24  (
    .i0(\PWMD/n12 [24]),
    .i1(freqD[24]),
    .sel(\PWMD/n0 ),
    .o(\PWMD/n13 [24]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMD/mux0_b25  (
    .i0(\PWMD/n12 [25]),
    .i1(freqD[25]),
    .sel(\PWMD/n0 ),
    .o(\PWMD/n13 [25]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMD/mux0_b26  (
    .i0(\PWMD/n12 [26]),
    .i1(freqD[26]),
    .sel(\PWMD/n0 ),
    .o(\PWMD/n13 [26]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMD/mux0_b3  (
    .i0(\PWMD/n12 [3]),
    .i1(freqD[3]),
    .sel(\PWMD/n0 ),
    .o(\PWMD/n13 [3]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMD/mux0_b4  (
    .i0(\PWMD/n12 [4]),
    .i1(freqD[4]),
    .sel(\PWMD/n0 ),
    .o(\PWMD/n13 [4]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMD/mux0_b5  (
    .i0(\PWMD/n12 [5]),
    .i1(freqD[5]),
    .sel(\PWMD/n0 ),
    .o(\PWMD/n13 [5]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMD/mux0_b6  (
    .i0(\PWMD/n12 [6]),
    .i1(freqD[6]),
    .sel(\PWMD/n0 ),
    .o(\PWMD/n13 [6]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMD/mux0_b7  (
    .i0(\PWMD/n12 [7]),
    .i1(freqD[7]),
    .sel(\PWMD/n0 ),
    .o(\PWMD/n13 [7]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMD/mux0_b8  (
    .i0(\PWMD/n12 [8]),
    .i1(freqD[8]),
    .sel(\PWMD/n0 ),
    .o(\PWMD/n13 [8]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMD/mux0_b9  (
    .i0(\PWMD/n12 [9]),
    .i1(freqD[9]),
    .sel(\PWMD/n0 ),
    .o(\PWMD/n13 [9]));  // src/OnePWM.v(32)
  and \PWMD/mux3_b0_sel_is_3  (\PWMD/mux3_b0_sel_is_3_o , \PWMD/n11 , \PWMD/n0 );
  binary_mux_s1_w1 \PWMD/mux4_b0  (
    .i0(\PWMD/pnumr [0]),
    .i1(1'b0),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n22 [0]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux4_b1  (
    .i0(\PWMD/pnumr [1]),
    .i1(1'b0),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n22 [1]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux4_b10  (
    .i0(\PWMD/pnumr [10]),
    .i1(1'b0),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n22 [10]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux4_b11  (
    .i0(\PWMD/pnumr [11]),
    .i1(1'b0),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n22 [11]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux4_b12  (
    .i0(\PWMD/pnumr [12]),
    .i1(1'b0),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n22 [12]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux4_b13  (
    .i0(\PWMD/pnumr [13]),
    .i1(1'b0),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n22 [13]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux4_b14  (
    .i0(\PWMD/pnumr [14]),
    .i1(1'b0),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n22 [14]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux4_b15  (
    .i0(\PWMD/pnumr [15]),
    .i1(1'b0),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n22 [15]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux4_b16  (
    .i0(\PWMD/pnumr [16]),
    .i1(1'b0),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n22 [16]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux4_b17  (
    .i0(\PWMD/pnumr [17]),
    .i1(1'b0),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n22 [17]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux4_b18  (
    .i0(\PWMD/pnumr [18]),
    .i1(1'b0),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n22 [18]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux4_b19  (
    .i0(\PWMD/pnumr [19]),
    .i1(1'b0),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n22 [19]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux4_b2  (
    .i0(\PWMD/pnumr [2]),
    .i1(1'b0),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n22 [2]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux4_b20  (
    .i0(\PWMD/pnumr [20]),
    .i1(1'b0),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n22 [20]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux4_b21  (
    .i0(\PWMD/pnumr [21]),
    .i1(1'b0),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n22 [21]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux4_b22  (
    .i0(\PWMD/pnumr [22]),
    .i1(1'b0),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n22 [22]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux4_b23  (
    .i0(\PWMD/pnumr [23]),
    .i1(1'b0),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n22 [23]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux4_b24  (
    .i0(\PWMD/pnumr [24]),
    .i1(1'b0),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n22 [24]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux4_b25  (
    .i0(\PWMD/pnumr [25]),
    .i1(1'b0),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n22 [25]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux4_b26  (
    .i0(\PWMD/pnumr [26]),
    .i1(1'b0),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n22 [26]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux4_b27  (
    .i0(\PWMD/pnumr [27]),
    .i1(1'b0),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n22 [27]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux4_b28  (
    .i0(\PWMD/pnumr [28]),
    .i1(1'b0),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n22 [28]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux4_b29  (
    .i0(\PWMD/pnumr [29]),
    .i1(1'b0),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n22 [29]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux4_b3  (
    .i0(\PWMD/pnumr [3]),
    .i1(1'b0),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n22 [3]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux4_b30  (
    .i0(\PWMD/pnumr [30]),
    .i1(1'b0),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n22 [30]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux4_b31  (
    .i0(\PWMD/pnumr [31]),
    .i1(1'b0),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n22 [31]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux4_b4  (
    .i0(\PWMD/pnumr [4]),
    .i1(1'b0),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n22 [4]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux4_b5  (
    .i0(\PWMD/pnumr [5]),
    .i1(1'b0),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n22 [5]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux4_b6  (
    .i0(\PWMD/pnumr [6]),
    .i1(1'b0),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n22 [6]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux4_b7  (
    .i0(\PWMD/pnumr [7]),
    .i1(1'b0),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n22 [7]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux4_b8  (
    .i0(\PWMD/pnumr [8]),
    .i1(1'b0),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n22 [8]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux4_b9  (
    .i0(\PWMD/pnumr [9]),
    .i1(1'b0),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n22 [9]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux5_b0  (
    .i0(\PWMD/n22 [0]),
    .i1(pnumD[0]),
    .sel(pnumD[32]),
    .o(\PWMD/n23 [0]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux5_b1  (
    .i0(\PWMD/n22 [1]),
    .i1(pnumD[1]),
    .sel(pnumD[32]),
    .o(\PWMD/n23 [1]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux5_b10  (
    .i0(\PWMD/n22 [10]),
    .i1(pnumD[10]),
    .sel(pnumD[32]),
    .o(\PWMD/n23 [10]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux5_b11  (
    .i0(\PWMD/n22 [11]),
    .i1(pnumD[11]),
    .sel(pnumD[32]),
    .o(\PWMD/n23 [11]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux5_b12  (
    .i0(\PWMD/n22 [12]),
    .i1(pnumD[12]),
    .sel(pnumD[32]),
    .o(\PWMD/n23 [12]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux5_b13  (
    .i0(\PWMD/n22 [13]),
    .i1(pnumD[13]),
    .sel(pnumD[32]),
    .o(\PWMD/n23 [13]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux5_b14  (
    .i0(\PWMD/n22 [14]),
    .i1(pnumD[14]),
    .sel(pnumD[32]),
    .o(\PWMD/n23 [14]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux5_b15  (
    .i0(\PWMD/n22 [15]),
    .i1(pnumD[15]),
    .sel(pnumD[32]),
    .o(\PWMD/n23 [15]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux5_b16  (
    .i0(\PWMD/n22 [16]),
    .i1(pnumD[16]),
    .sel(pnumD[32]),
    .o(\PWMD/n23 [16]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux5_b17  (
    .i0(\PWMD/n22 [17]),
    .i1(pnumD[17]),
    .sel(pnumD[32]),
    .o(\PWMD/n23 [17]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux5_b18  (
    .i0(\PWMD/n22 [18]),
    .i1(pnumD[18]),
    .sel(pnumD[32]),
    .o(\PWMD/n23 [18]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux5_b19  (
    .i0(\PWMD/n22 [19]),
    .i1(pnumD[19]),
    .sel(pnumD[32]),
    .o(\PWMD/n23 [19]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux5_b2  (
    .i0(\PWMD/n22 [2]),
    .i1(pnumD[2]),
    .sel(pnumD[32]),
    .o(\PWMD/n23 [2]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux5_b20  (
    .i0(\PWMD/n22 [20]),
    .i1(pnumD[20]),
    .sel(pnumD[32]),
    .o(\PWMD/n23 [20]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux5_b21  (
    .i0(\PWMD/n22 [21]),
    .i1(pnumD[21]),
    .sel(pnumD[32]),
    .o(\PWMD/n23 [21]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux5_b22  (
    .i0(\PWMD/n22 [22]),
    .i1(pnumD[22]),
    .sel(pnumD[32]),
    .o(\PWMD/n23 [22]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux5_b23  (
    .i0(\PWMD/n22 [23]),
    .i1(pnumD[23]),
    .sel(pnumD[32]),
    .o(\PWMD/n23 [23]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux5_b24  (
    .i0(\PWMD/n22 [24]),
    .i1(pnumD[24]),
    .sel(pnumD[32]),
    .o(\PWMD/n23 [24]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux5_b25  (
    .i0(\PWMD/n22 [25]),
    .i1(pnumD[25]),
    .sel(pnumD[32]),
    .o(\PWMD/n23 [25]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux5_b26  (
    .i0(\PWMD/n22 [26]),
    .i1(pnumD[26]),
    .sel(pnumD[32]),
    .o(\PWMD/n23 [26]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux5_b27  (
    .i0(\PWMD/n22 [27]),
    .i1(pnumD[27]),
    .sel(pnumD[32]),
    .o(\PWMD/n23 [27]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux5_b28  (
    .i0(\PWMD/n22 [28]),
    .i1(pnumD[28]),
    .sel(pnumD[32]),
    .o(\PWMD/n23 [28]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux5_b29  (
    .i0(\PWMD/n22 [29]),
    .i1(pnumD[29]),
    .sel(pnumD[32]),
    .o(\PWMD/n23 [29]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux5_b3  (
    .i0(\PWMD/n22 [3]),
    .i1(pnumD[3]),
    .sel(pnumD[32]),
    .o(\PWMD/n23 [3]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux5_b30  (
    .i0(\PWMD/n22 [30]),
    .i1(pnumD[30]),
    .sel(pnumD[32]),
    .o(\PWMD/n23 [30]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux5_b31  (
    .i0(\PWMD/n22 [31]),
    .i1(pnumD[31]),
    .sel(pnumD[32]),
    .o(\PWMD/n23 [31]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux5_b4  (
    .i0(\PWMD/n22 [4]),
    .i1(pnumD[4]),
    .sel(pnumD[32]),
    .o(\PWMD/n23 [4]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux5_b5  (
    .i0(\PWMD/n22 [5]),
    .i1(pnumD[5]),
    .sel(pnumD[32]),
    .o(\PWMD/n23 [5]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux5_b6  (
    .i0(\PWMD/n22 [6]),
    .i1(pnumD[6]),
    .sel(pnumD[32]),
    .o(\PWMD/n23 [6]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux5_b7  (
    .i0(\PWMD/n22 [7]),
    .i1(pnumD[7]),
    .sel(pnumD[32]),
    .o(\PWMD/n23 [7]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux5_b8  (
    .i0(\PWMD/n22 [8]),
    .i1(pnumD[8]),
    .sel(pnumD[32]),
    .o(\PWMD/n23 [8]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux5_b9  (
    .i0(\PWMD/n22 [9]),
    .i1(pnumD[9]),
    .sel(pnumD[32]),
    .o(\PWMD/n23 [9]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMD/mux6_b0  (
    .i0(\PWMD/pnumr [0]),
    .i1(\PWMD/n26 [0]),
    .sel(\PWMD/n25 ),
    .o(\PWMD/n27 [0]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMD/mux6_b1  (
    .i0(\PWMD/pnumr [1]),
    .i1(\PWMD/n26 [1]),
    .sel(\PWMD/n25 ),
    .o(\PWMD/n27 [1]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMD/mux6_b10  (
    .i0(\PWMD/pnumr [10]),
    .i1(\PWMD/n26 [10]),
    .sel(\PWMD/n25 ),
    .o(\PWMD/n27 [10]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMD/mux6_b11  (
    .i0(\PWMD/pnumr [11]),
    .i1(\PWMD/n26 [11]),
    .sel(\PWMD/n25 ),
    .o(\PWMD/n27 [11]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMD/mux6_b12  (
    .i0(\PWMD/pnumr [12]),
    .i1(\PWMD/n26 [12]),
    .sel(\PWMD/n25 ),
    .o(\PWMD/n27 [12]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMD/mux6_b13  (
    .i0(\PWMD/pnumr [13]),
    .i1(\PWMD/n26 [13]),
    .sel(\PWMD/n25 ),
    .o(\PWMD/n27 [13]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMD/mux6_b14  (
    .i0(\PWMD/pnumr [14]),
    .i1(\PWMD/n26 [14]),
    .sel(\PWMD/n25 ),
    .o(\PWMD/n27 [14]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMD/mux6_b15  (
    .i0(\PWMD/pnumr [15]),
    .i1(\PWMD/n26 [15]),
    .sel(\PWMD/n25 ),
    .o(\PWMD/n27 [15]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMD/mux6_b16  (
    .i0(\PWMD/pnumr [16]),
    .i1(\PWMD/n26 [16]),
    .sel(\PWMD/n25 ),
    .o(\PWMD/n27 [16]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMD/mux6_b17  (
    .i0(\PWMD/pnumr [17]),
    .i1(\PWMD/n26 [17]),
    .sel(\PWMD/n25 ),
    .o(\PWMD/n27 [17]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMD/mux6_b18  (
    .i0(\PWMD/pnumr [18]),
    .i1(\PWMD/n26 [18]),
    .sel(\PWMD/n25 ),
    .o(\PWMD/n27 [18]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMD/mux6_b19  (
    .i0(\PWMD/pnumr [19]),
    .i1(\PWMD/n26 [19]),
    .sel(\PWMD/n25 ),
    .o(\PWMD/n27 [19]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMD/mux6_b2  (
    .i0(\PWMD/pnumr [2]),
    .i1(\PWMD/n26 [2]),
    .sel(\PWMD/n25 ),
    .o(\PWMD/n27 [2]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMD/mux6_b20  (
    .i0(\PWMD/pnumr [20]),
    .i1(\PWMD/n26 [20]),
    .sel(\PWMD/n25 ),
    .o(\PWMD/n27 [20]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMD/mux6_b21  (
    .i0(\PWMD/pnumr [21]),
    .i1(\PWMD/n26 [21]),
    .sel(\PWMD/n25 ),
    .o(\PWMD/n27 [21]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMD/mux6_b22  (
    .i0(\PWMD/pnumr [22]),
    .i1(\PWMD/n26 [22]),
    .sel(\PWMD/n25 ),
    .o(\PWMD/n27 [22]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMD/mux6_b23  (
    .i0(\PWMD/pnumr [23]),
    .i1(\PWMD/n26 [23]),
    .sel(\PWMD/n25 ),
    .o(\PWMD/n27 [23]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMD/mux6_b3  (
    .i0(\PWMD/pnumr [3]),
    .i1(\PWMD/n26 [3]),
    .sel(\PWMD/n25 ),
    .o(\PWMD/n27 [3]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMD/mux6_b4  (
    .i0(\PWMD/pnumr [4]),
    .i1(\PWMD/n26 [4]),
    .sel(\PWMD/n25 ),
    .o(\PWMD/n27 [4]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMD/mux6_b5  (
    .i0(\PWMD/pnumr [5]),
    .i1(\PWMD/n26 [5]),
    .sel(\PWMD/n25 ),
    .o(\PWMD/n27 [5]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMD/mux6_b6  (
    .i0(\PWMD/pnumr [6]),
    .i1(\PWMD/n26 [6]),
    .sel(\PWMD/n25 ),
    .o(\PWMD/n27 [6]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMD/mux6_b7  (
    .i0(\PWMD/pnumr [7]),
    .i1(\PWMD/n26 [7]),
    .sel(\PWMD/n25 ),
    .o(\PWMD/n27 [7]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMD/mux6_b8  (
    .i0(\PWMD/pnumr [8]),
    .i1(\PWMD/n26 [8]),
    .sel(\PWMD/n25 ),
    .o(\PWMD/n27 [8]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMD/mux6_b9  (
    .i0(\PWMD/pnumr [9]),
    .i1(\PWMD/n26 [9]),
    .sel(\PWMD/n25 ),
    .o(\PWMD/n27 [9]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMD/mux7_b0  (
    .i0(pnumcntD[0]),
    .i1(\PWMD/n27 [0]),
    .sel(\PWMD/n24 ),
    .o(\PWMD/n29 [0]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux7_b1  (
    .i0(pnumcntD[1]),
    .i1(\PWMD/n27 [1]),
    .sel(\PWMD/n24 ),
    .o(\PWMD/n29 [1]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux7_b10  (
    .i0(pnumcntD[10]),
    .i1(\PWMD/n27 [10]),
    .sel(\PWMD/n24 ),
    .o(\PWMD/n29 [10]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux7_b11  (
    .i0(pnumcntD[11]),
    .i1(\PWMD/n27 [11]),
    .sel(\PWMD/n24 ),
    .o(\PWMD/n29 [11]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux7_b12  (
    .i0(pnumcntD[12]),
    .i1(\PWMD/n27 [12]),
    .sel(\PWMD/n24 ),
    .o(\PWMD/n29 [12]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux7_b13  (
    .i0(pnumcntD[13]),
    .i1(\PWMD/n27 [13]),
    .sel(\PWMD/n24 ),
    .o(\PWMD/n29 [13]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux7_b14  (
    .i0(pnumcntD[14]),
    .i1(\PWMD/n27 [14]),
    .sel(\PWMD/n24 ),
    .o(\PWMD/n29 [14]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux7_b15  (
    .i0(pnumcntD[15]),
    .i1(\PWMD/n27 [15]),
    .sel(\PWMD/n24 ),
    .o(\PWMD/n29 [15]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux7_b16  (
    .i0(pnumcntD[16]),
    .i1(\PWMD/n27 [16]),
    .sel(\PWMD/n24 ),
    .o(\PWMD/n29 [16]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux7_b17  (
    .i0(pnumcntD[17]),
    .i1(\PWMD/n27 [17]),
    .sel(\PWMD/n24 ),
    .o(\PWMD/n29 [17]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux7_b18  (
    .i0(pnumcntD[18]),
    .i1(\PWMD/n27 [18]),
    .sel(\PWMD/n24 ),
    .o(\PWMD/n29 [18]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux7_b19  (
    .i0(pnumcntD[19]),
    .i1(\PWMD/n27 [19]),
    .sel(\PWMD/n24 ),
    .o(\PWMD/n29 [19]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux7_b2  (
    .i0(pnumcntD[2]),
    .i1(\PWMD/n27 [2]),
    .sel(\PWMD/n24 ),
    .o(\PWMD/n29 [2]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux7_b20  (
    .i0(pnumcntD[20]),
    .i1(\PWMD/n27 [20]),
    .sel(\PWMD/n24 ),
    .o(\PWMD/n29 [20]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux7_b21  (
    .i0(pnumcntD[21]),
    .i1(\PWMD/n27 [21]),
    .sel(\PWMD/n24 ),
    .o(\PWMD/n29 [21]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux7_b22  (
    .i0(pnumcntD[22]),
    .i1(\PWMD/n27 [22]),
    .sel(\PWMD/n24 ),
    .o(\PWMD/n29 [22]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux7_b23  (
    .i0(pnumcntD[23]),
    .i1(\PWMD/n27 [23]),
    .sel(\PWMD/n24 ),
    .o(\PWMD/n29 [23]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux7_b3  (
    .i0(pnumcntD[3]),
    .i1(\PWMD/n27 [3]),
    .sel(\PWMD/n24 ),
    .o(\PWMD/n29 [3]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux7_b4  (
    .i0(pnumcntD[4]),
    .i1(\PWMD/n27 [4]),
    .sel(\PWMD/n24 ),
    .o(\PWMD/n29 [4]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux7_b5  (
    .i0(pnumcntD[5]),
    .i1(\PWMD/n27 [5]),
    .sel(\PWMD/n24 ),
    .o(\PWMD/n29 [5]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux7_b6  (
    .i0(pnumcntD[6]),
    .i1(\PWMD/n27 [6]),
    .sel(\PWMD/n24 ),
    .o(\PWMD/n29 [6]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux7_b7  (
    .i0(pnumcntD[7]),
    .i1(\PWMD/n27 [7]),
    .sel(\PWMD/n24 ),
    .o(\PWMD/n29 [7]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux7_b8  (
    .i0(pnumcntD[8]),
    .i1(\PWMD/n27 [8]),
    .sel(\PWMD/n24 ),
    .o(\PWMD/n29 [8]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux7_b9  (
    .i0(pnumcntD[9]),
    .i1(\PWMD/n27 [9]),
    .sel(\PWMD/n24 ),
    .o(\PWMD/n29 [9]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux8_b0  (
    .i0(\PWMD/n29 [0]),
    .i1(\PWMD/pnumr [0]),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n31 [0]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux8_b1  (
    .i0(\PWMD/n29 [1]),
    .i1(\PWMD/pnumr [1]),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n31 [1]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux8_b10  (
    .i0(\PWMD/n29 [10]),
    .i1(\PWMD/pnumr [10]),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n31 [10]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux8_b11  (
    .i0(\PWMD/n29 [11]),
    .i1(\PWMD/pnumr [11]),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n31 [11]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux8_b12  (
    .i0(\PWMD/n29 [12]),
    .i1(\PWMD/pnumr [12]),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n31 [12]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux8_b13  (
    .i0(\PWMD/n29 [13]),
    .i1(\PWMD/pnumr [13]),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n31 [13]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux8_b14  (
    .i0(\PWMD/n29 [14]),
    .i1(\PWMD/pnumr [14]),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n31 [14]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux8_b15  (
    .i0(\PWMD/n29 [15]),
    .i1(\PWMD/pnumr [15]),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n31 [15]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux8_b16  (
    .i0(\PWMD/n29 [16]),
    .i1(\PWMD/pnumr [16]),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n31 [16]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux8_b17  (
    .i0(\PWMD/n29 [17]),
    .i1(\PWMD/pnumr [17]),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n31 [17]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux8_b18  (
    .i0(\PWMD/n29 [18]),
    .i1(\PWMD/pnumr [18]),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n31 [18]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux8_b19  (
    .i0(\PWMD/n29 [19]),
    .i1(\PWMD/pnumr [19]),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n31 [19]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux8_b2  (
    .i0(\PWMD/n29 [2]),
    .i1(\PWMD/pnumr [2]),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n31 [2]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux8_b20  (
    .i0(\PWMD/n29 [20]),
    .i1(\PWMD/pnumr [20]),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n31 [20]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux8_b21  (
    .i0(\PWMD/n29 [21]),
    .i1(\PWMD/pnumr [21]),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n31 [21]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux8_b22  (
    .i0(\PWMD/n29 [22]),
    .i1(\PWMD/pnumr [22]),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n31 [22]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux8_b23  (
    .i0(\PWMD/n29 [23]),
    .i1(\PWMD/pnumr [23]),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n31 [23]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux8_b3  (
    .i0(\PWMD/n29 [3]),
    .i1(\PWMD/pnumr [3]),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n31 [3]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux8_b4  (
    .i0(\PWMD/n29 [4]),
    .i1(\PWMD/pnumr [4]),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n31 [4]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux8_b5  (
    .i0(\PWMD/n29 [5]),
    .i1(\PWMD/pnumr [5]),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n31 [5]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux8_b6  (
    .i0(\PWMD/n29 [6]),
    .i1(\PWMD/pnumr [6]),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n31 [6]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux8_b7  (
    .i0(\PWMD/n29 [7]),
    .i1(\PWMD/pnumr [7]),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n31 [7]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux8_b8  (
    .i0(\PWMD/n29 [8]),
    .i1(\PWMD/pnumr [8]),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n31 [8]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMD/mux8_b9  (
    .i0(\PWMD/n29 [9]),
    .i1(\PWMD/pnumr [9]),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n31 [9]));  // src/OnePWM.v(57)
  not \PWMD/n17_inv  (\PWMD/n17_neg , \PWMD/n17 );
  not \PWMD/n25_inv  (\PWMD/n25_neg , \PWMD/n25 );
  not \PWMD/n4_inv  (\PWMD/n4_neg , \PWMD/n4 );
  not \PWMD/n6_inv  (\PWMD/n6_neg , \PWMD/n6 );
  ne_w24 \PWMD/neq0  (
    .i0(pnumcntD),
    .i1(24'b000000000000000000000000),
    .o(\PWMD/n25 ));  // src/OnePWM.v(55)
  reg_sr_ss_w1 \PWMD/pwm_reg  (
    .clk(clk100m),
    .d(pwm[13]),
    .en(1'b1),
    .reset(~\PWMD/u14_sel_is_1_o ),
    .set(\PWMD/n18 ),
    .q(\PWMD/pwm_keep ));  // src/OnePWM.v(45)
  reg_sr_as_w1 \PWMD/reg0_b0  (
    .clk(clk100m),
    .d(\PWMD/n13 [0]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [0]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b1  (
    .clk(clk100m),
    .d(\PWMD/n13 [1]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [1]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b10  (
    .clk(clk100m),
    .d(\PWMD/n13 [10]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [10]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b11  (
    .clk(clk100m),
    .d(\PWMD/n13 [11]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [11]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b12  (
    .clk(clk100m),
    .d(\PWMD/n13 [12]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [12]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b13  (
    .clk(clk100m),
    .d(\PWMD/n13 [13]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [13]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b14  (
    .clk(clk100m),
    .d(\PWMD/n13 [14]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [14]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b15  (
    .clk(clk100m),
    .d(\PWMD/n13 [15]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [15]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b16  (
    .clk(clk100m),
    .d(\PWMD/n13 [16]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [16]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b17  (
    .clk(clk100m),
    .d(\PWMD/n13 [17]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [17]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b18  (
    .clk(clk100m),
    .d(\PWMD/n13 [18]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [18]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b19  (
    .clk(clk100m),
    .d(\PWMD/n13 [19]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [19]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b2  (
    .clk(clk100m),
    .d(\PWMD/n13 [2]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [2]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b20  (
    .clk(clk100m),
    .d(\PWMD/n13 [20]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [20]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b21  (
    .clk(clk100m),
    .d(\PWMD/n13 [21]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [21]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b22  (
    .clk(clk100m),
    .d(\PWMD/n13 [22]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [22]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b23  (
    .clk(clk100m),
    .d(\PWMD/n13 [23]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [23]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b24  (
    .clk(clk100m),
    .d(\PWMD/n13 [24]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [24]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b25  (
    .clk(clk100m),
    .d(\PWMD/n13 [25]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [25]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b26  (
    .clk(clk100m),
    .d(\PWMD/n13 [26]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [26]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b3  (
    .clk(clk100m),
    .d(\PWMD/n13 [3]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [3]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b4  (
    .clk(clk100m),
    .d(\PWMD/n13 [4]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [4]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b5  (
    .clk(clk100m),
    .d(\PWMD/n13 [5]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [5]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b6  (
    .clk(clk100m),
    .d(\PWMD/n13 [6]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [6]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b7  (
    .clk(clk100m),
    .d(\PWMD/n13 [7]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [7]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b8  (
    .clk(clk100m),
    .d(\PWMD/n13 [8]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [8]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMD/reg0_b9  (
    .clk(clk100m),
    .d(\PWMD/n13 [9]),
    .en(1'b1),
    .reset(~\PWMD/n11 ),
    .set(1'b0),
    .q(\PWMD/FreCnt [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b0  (
    .clk(clk100m),
    .d(freqD[0]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [0]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b1  (
    .clk(clk100m),
    .d(freqD[1]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [1]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b10  (
    .clk(clk100m),
    .d(freqD[10]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [10]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b11  (
    .clk(clk100m),
    .d(freqD[11]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [11]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b12  (
    .clk(clk100m),
    .d(freqD[12]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [12]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b13  (
    .clk(clk100m),
    .d(freqD[13]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [13]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b14  (
    .clk(clk100m),
    .d(freqD[14]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [14]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b15  (
    .clk(clk100m),
    .d(freqD[15]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [15]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b16  (
    .clk(clk100m),
    .d(freqD[16]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [16]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b17  (
    .clk(clk100m),
    .d(freqD[17]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [17]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b18  (
    .clk(clk100m),
    .d(freqD[18]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [18]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b19  (
    .clk(clk100m),
    .d(freqD[19]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [19]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b2  (
    .clk(clk100m),
    .d(freqD[2]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [2]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b20  (
    .clk(clk100m),
    .d(freqD[20]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [20]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b21  (
    .clk(clk100m),
    .d(freqD[21]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [21]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b22  (
    .clk(clk100m),
    .d(freqD[22]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [22]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b23  (
    .clk(clk100m),
    .d(freqD[23]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [23]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b24  (
    .clk(clk100m),
    .d(freqD[24]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [24]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b25  (
    .clk(clk100m),
    .d(freqD[25]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [25]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b26  (
    .clk(clk100m),
    .d(freqD[26]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [26]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b3  (
    .clk(clk100m),
    .d(freqD[3]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [3]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b4  (
    .clk(clk100m),
    .d(freqD[4]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [4]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b5  (
    .clk(clk100m),
    .d(freqD[5]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [5]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b6  (
    .clk(clk100m),
    .d(freqD[6]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [6]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b7  (
    .clk(clk100m),
    .d(freqD[7]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [7]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b8  (
    .clk(clk100m),
    .d(freqD[8]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [8]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg1_b9  (
    .clk(clk100m),
    .d(freqD[9]),
    .en(\PWMD/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/FreCntr [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMD/reg2_b0  (
    .clk(clk100m),
    .d(\PWMD/n23 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[0]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b1  (
    .clk(clk100m),
    .d(\PWMD/n23 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[1]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b10  (
    .clk(clk100m),
    .d(\PWMD/n23 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[10]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b11  (
    .clk(clk100m),
    .d(\PWMD/n23 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[11]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b12  (
    .clk(clk100m),
    .d(\PWMD/n23 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[12]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b13  (
    .clk(clk100m),
    .d(\PWMD/n23 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[13]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b14  (
    .clk(clk100m),
    .d(\PWMD/n23 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[14]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b15  (
    .clk(clk100m),
    .d(\PWMD/n23 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[15]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b16  (
    .clk(clk100m),
    .d(\PWMD/n23 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[16]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b17  (
    .clk(clk100m),
    .d(\PWMD/n23 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[17]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b18  (
    .clk(clk100m),
    .d(\PWMD/n23 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[18]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b19  (
    .clk(clk100m),
    .d(\PWMD/n23 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[19]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b2  (
    .clk(clk100m),
    .d(\PWMD/n23 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[2]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b20  (
    .clk(clk100m),
    .d(\PWMD/n23 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[20]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b21  (
    .clk(clk100m),
    .d(\PWMD/n23 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[21]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b22  (
    .clk(clk100m),
    .d(\PWMD/n23 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[22]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b23  (
    .clk(clk100m),
    .d(\PWMD/n23 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[23]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b24  (
    .clk(clk100m),
    .d(\PWMD/n23 [24]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[24]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b25  (
    .clk(clk100m),
    .d(\PWMD/n23 [25]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[25]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b26  (
    .clk(clk100m),
    .d(\PWMD/n23 [26]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[26]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b27  (
    .clk(clk100m),
    .d(\PWMD/n23 [27]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[27]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b28  (
    .clk(clk100m),
    .d(\PWMD/n23 [28]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[28]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b29  (
    .clk(clk100m),
    .d(\PWMD/n23 [29]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[29]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b3  (
    .clk(clk100m),
    .d(\PWMD/n23 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[3]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b30  (
    .clk(clk100m),
    .d(\PWMD/n23 [30]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[30]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b31  (
    .clk(clk100m),
    .d(\PWMD/n23 [31]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[31]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b4  (
    .clk(clk100m),
    .d(\PWMD/n23 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[4]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b5  (
    .clk(clk100m),
    .d(\PWMD/n23 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[5]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b6  (
    .clk(clk100m),
    .d(\PWMD/n23 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[6]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b7  (
    .clk(clk100m),
    .d(\PWMD/n23 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[7]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b8  (
    .clk(clk100m),
    .d(\PWMD/n23 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[8]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg2_b9  (
    .clk(clk100m),
    .d(\PWMD/n23 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/pnumr[9]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMD/reg3_b0  (
    .clk(clk100m),
    .d(\PWMD/n31 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[0]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b1  (
    .clk(clk100m),
    .d(\PWMD/n31 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[1]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b10  (
    .clk(clk100m),
    .d(\PWMD/n31 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[10]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b11  (
    .clk(clk100m),
    .d(\PWMD/n31 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[11]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b12  (
    .clk(clk100m),
    .d(\PWMD/n31 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[12]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b13  (
    .clk(clk100m),
    .d(\PWMD/n31 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[13]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b14  (
    .clk(clk100m),
    .d(\PWMD/n31 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[14]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b15  (
    .clk(clk100m),
    .d(\PWMD/n31 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[15]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b16  (
    .clk(clk100m),
    .d(\PWMD/n31 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[16]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b17  (
    .clk(clk100m),
    .d(\PWMD/n31 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[17]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b18  (
    .clk(clk100m),
    .d(\PWMD/n31 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[18]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b19  (
    .clk(clk100m),
    .d(\PWMD/n31 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[19]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b2  (
    .clk(clk100m),
    .d(\PWMD/n31 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[2]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b20  (
    .clk(clk100m),
    .d(\PWMD/n31 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[20]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b21  (
    .clk(clk100m),
    .d(\PWMD/n31 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[21]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b22  (
    .clk(clk100m),
    .d(\PWMD/n31 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[22]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b23  (
    .clk(clk100m),
    .d(\PWMD/n31 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[23]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b3  (
    .clk(clk100m),
    .d(\PWMD/n31 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[3]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b4  (
    .clk(clk100m),
    .d(\PWMD/n31 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[4]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b5  (
    .clk(clk100m),
    .d(\PWMD/n31 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[5]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b6  (
    .clk(clk100m),
    .d(\PWMD/n31 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[6]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b7  (
    .clk(clk100m),
    .d(\PWMD/n31 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[7]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b8  (
    .clk(clk100m),
    .d(\PWMD/n31 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[8]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMD/reg3_b9  (
    .clk(clk100m),
    .d(\PWMD/n31 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMD/RemaTxNum[9]_keep ));  // src/OnePWM.v(58)
  reg_ar_ss_w1 \PWMD/stopreq_reg  (
    .clk(clk100m),
    .d(\PWMD/n1 ),
    .en(1'b1),
    .reset(1'b0),
    .set(pwm_start_stop[13]),
    .q(\PWMD/stopreq_keep ));  // src/OnePWM.v(15)
  add_pu27_mu27_o27 \PWMD/sub0  (
    .i0(\PWMD/FreCnt ),
    .i1(27'b000000000000000000000000001),
    .o(\PWMD/n12 [26:0]));  // src/OnePWM.v(32)
  add_pu24_mu24_o24 \PWMD/sub1  (
    .i0(pnumcntD),
    .i1(24'b000000000000000000000001),
    .o(\PWMD/n26 [23:0]));  // src/OnePWM.v(55)
  AL_MUX \PWMD/u10  (
    .i0(1'b0),
    .i1(\PWMD/n9 ),
    .sel(n24),
    .o(\PWMD/n10 ));  // src/OnePWM.v(26)
  or \PWMD/u11  (\PWMD/n11 , pwm_state_read[13], pwm_start_stop[29]);  // src/OnePWM.v(30)
  and \PWMD/u14_sel_is_1  (\PWMD/u14_sel_is_1_o , pwm_state_read[13], \PWMD/n17_neg );
  and \PWMD/u15  (\PWMD/n24 , \PWMD/n0 , pwm_state_read[13]);  // src/OnePWM.v(54)
  and \PWMD/u17_sel_is_1  (\PWMD/u17_sel_is_1_o , \PWMD/n24 , \PWMD/n25_neg );
  not \PWMD/u17_sel_is_1_o_inv  (\PWMD/u17_sel_is_1_o_neg , \PWMD/u17_sel_is_1_o );
  AL_MUX \PWMD/u18  (
    .i0(\PWMD/pnumr [31]),
    .i1(dir[13]),
    .sel(\PWMD/u18_sel_is_0_o ),
    .o(\PWMD/n32 ));
  and \PWMD/u18_sel_is_0  (\PWMD/u18_sel_is_0_o , \pwm_start_stop[29]_neg , \PWMD/u17_sel_is_1_o_neg );
  AL_MUX \PWMD/u2  (
    .i0(\PWMD/stopreq ),
    .i1(1'b0),
    .sel(\PWMD/n0 ),
    .o(\PWMD/n1 ));  // src/OnePWM.v(15)
  and \PWMD/u5  (\PWMD/n4 , \PWMD/stopreq , \PWMD/n0 );  // src/OnePWM.v(23)
  and \PWMD/u6  (\PWMD/n6 , \PWMD/n5 , \PWMD/n0 );  // src/OnePWM.v(25)
  AL_MUX \PWMD/u8  (
    .i0(1'b0),
    .i1(pwm_state_read[13]),
    .sel(\PWMD/u8_sel_is_0_o ),
    .o(\PWMD/n8 ));
  and \PWMD/u8_sel_is_0  (\PWMD/u8_sel_is_0_o , \PWMD/n4_neg , \PWMD/n6_neg );
  AL_MUX \PWMD/u9  (
    .i0(\PWMD/n8 ),
    .i1(1'b1),
    .sel(pwm_start_stop[29]),
    .o(\PWMD/n9 ));  // src/OnePWM.v(26)
  reg_ar_as_w1 \PWME/State_reg  (
    .clk(clk100m),
    .d(\PWME/n10 ),
    .en(1'b1),
    .reset(~rstn),
    .set(1'b0),
    .q(pwm_state_read[14]));  // src/OnePWM.v(26)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[0]  (
    .i(\PWME/RemaTxNum[0]_keep ),
    .o(pnumcntE[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[10]  (
    .i(\PWME/RemaTxNum[10]_keep ),
    .o(pnumcntE[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[11]  (
    .i(\PWME/RemaTxNum[11]_keep ),
    .o(pnumcntE[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[12]  (
    .i(\PWME/RemaTxNum[12]_keep ),
    .o(pnumcntE[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[13]  (
    .i(\PWME/RemaTxNum[13]_keep ),
    .o(pnumcntE[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[14]  (
    .i(\PWME/RemaTxNum[14]_keep ),
    .o(pnumcntE[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[15]  (
    .i(\PWME/RemaTxNum[15]_keep ),
    .o(pnumcntE[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[16]  (
    .i(\PWME/RemaTxNum[16]_keep ),
    .o(pnumcntE[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[17]  (
    .i(\PWME/RemaTxNum[17]_keep ),
    .o(pnumcntE[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[18]  (
    .i(\PWME/RemaTxNum[18]_keep ),
    .o(pnumcntE[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[19]  (
    .i(\PWME/RemaTxNum[19]_keep ),
    .o(pnumcntE[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[1]  (
    .i(\PWME/RemaTxNum[1]_keep ),
    .o(pnumcntE[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[20]  (
    .i(\PWME/RemaTxNum[20]_keep ),
    .o(pnumcntE[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[21]  (
    .i(\PWME/RemaTxNum[21]_keep ),
    .o(pnumcntE[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[22]  (
    .i(\PWME/RemaTxNum[22]_keep ),
    .o(pnumcntE[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[23]  (
    .i(\PWME/RemaTxNum[23]_keep ),
    .o(pnumcntE[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[2]  (
    .i(\PWME/RemaTxNum[2]_keep ),
    .o(pnumcntE[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[3]  (
    .i(\PWME/RemaTxNum[3]_keep ),
    .o(pnumcntE[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[4]  (
    .i(\PWME/RemaTxNum[4]_keep ),
    .o(pnumcntE[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[5]  (
    .i(\PWME/RemaTxNum[5]_keep ),
    .o(pnumcntE[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[6]  (
    .i(\PWME/RemaTxNum[6]_keep ),
    .o(pnumcntE[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[7]  (
    .i(\PWME/RemaTxNum[7]_keep ),
    .o(pnumcntE[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[8]  (
    .i(\PWME/RemaTxNum[8]_keep ),
    .o(pnumcntE[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_RemaTxNum[9]  (
    .i(\PWME/RemaTxNum[9]_keep ),
    .o(pnumcntE[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_dir  (
    .i(\PWME/dir_keep ),
    .o(dir[14]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[0]  (
    .i(\PWME/pnumr[0]_keep ),
    .o(\PWME/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[10]  (
    .i(\PWME/pnumr[10]_keep ),
    .o(\PWME/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[11]  (
    .i(\PWME/pnumr[11]_keep ),
    .o(\PWME/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[12]  (
    .i(\PWME/pnumr[12]_keep ),
    .o(\PWME/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[13]  (
    .i(\PWME/pnumr[13]_keep ),
    .o(\PWME/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[14]  (
    .i(\PWME/pnumr[14]_keep ),
    .o(\PWME/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[15]  (
    .i(\PWME/pnumr[15]_keep ),
    .o(\PWME/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[16]  (
    .i(\PWME/pnumr[16]_keep ),
    .o(\PWME/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[17]  (
    .i(\PWME/pnumr[17]_keep ),
    .o(\PWME/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[18]  (
    .i(\PWME/pnumr[18]_keep ),
    .o(\PWME/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[19]  (
    .i(\PWME/pnumr[19]_keep ),
    .o(\PWME/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[1]  (
    .i(\PWME/pnumr[1]_keep ),
    .o(\PWME/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[20]  (
    .i(\PWME/pnumr[20]_keep ),
    .o(\PWME/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[21]  (
    .i(\PWME/pnumr[21]_keep ),
    .o(\PWME/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[22]  (
    .i(\PWME/pnumr[22]_keep ),
    .o(\PWME/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[23]  (
    .i(\PWME/pnumr[23]_keep ),
    .o(\PWME/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[24]  (
    .i(\PWME/pnumr[24]_keep ),
    .o(\PWME/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[25]  (
    .i(\PWME/pnumr[25]_keep ),
    .o(\PWME/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[26]  (
    .i(\PWME/pnumr[26]_keep ),
    .o(\PWME/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[27]  (
    .i(\PWME/pnumr[27]_keep ),
    .o(\PWME/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[28]  (
    .i(\PWME/pnumr[28]_keep ),
    .o(\PWME/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[29]  (
    .i(\PWME/pnumr[29]_keep ),
    .o(\PWME/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[2]  (
    .i(\PWME/pnumr[2]_keep ),
    .o(\PWME/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[30]  (
    .i(\PWME/pnumr[30]_keep ),
    .o(\PWME/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[31]  (
    .i(\PWME/pnumr[31]_keep ),
    .o(\PWME/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[3]  (
    .i(\PWME/pnumr[3]_keep ),
    .o(\PWME/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[4]  (
    .i(\PWME/pnumr[4]_keep ),
    .o(\PWME/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[5]  (
    .i(\PWME/pnumr[5]_keep ),
    .o(\PWME/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[6]  (
    .i(\PWME/pnumr[6]_keep ),
    .o(\PWME/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[7]  (
    .i(\PWME/pnumr[7]_keep ),
    .o(\PWME/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[8]  (
    .i(\PWME/pnumr[8]_keep ),
    .o(\PWME/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pnumr[9]  (
    .i(\PWME/pnumr[9]_keep ),
    .o(\PWME/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_pwm  (
    .i(\PWME/pwm_keep ),
    .o(pwm[14]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWME/_bufkeep_stopreq  (
    .i(\PWME/stopreq_keep ),
    .o(\PWME/stopreq ));  // src/OnePWM.v(14)
  reg_ar_as_w1 \PWME/dir_reg  (
    .clk(clk100m),
    .d(\PWME/n32 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/dir_keep ));  // src/OnePWM.v(58)
  eq_w27 \PWME/eq0  (
    .i0(\PWME/FreCnt ),
    .i1(27'b000000000000000000000000000),
    .o(\PWME/n0 ));  // src/OnePWM.v(15)
  eq_w24 \PWME/eq1  (
    .i0(pnumcntE),
    .i1(24'b000000000000000000000001),
    .o(\PWME/n5 ));  // src/OnePWM.v(25)
  eq_w27 \PWME/eq2  (
    .i0(\PWME/FreCnt ),
    .i1({1'b0,\PWME/FreCntr [26:1]}),
    .o(\PWME/n17 ));  // src/OnePWM.v(41)
  eq_w27 \PWME/eq3  (
    .i0(\PWME/FreCnt ),
    .i1(\PWME/FreCntr ),
    .o(\PWME/n18 ));  // src/OnePWM.v(43)
  binary_mux_s1_w1 \PWME/mux0_b0  (
    .i0(\PWME/n12 [0]),
    .i1(freqE[0]),
    .sel(\PWME/n0 ),
    .o(\PWME/n13 [0]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWME/mux0_b1  (
    .i0(\PWME/n12 [1]),
    .i1(freqE[1]),
    .sel(\PWME/n0 ),
    .o(\PWME/n13 [1]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWME/mux0_b10  (
    .i0(\PWME/n12 [10]),
    .i1(freqE[10]),
    .sel(\PWME/n0 ),
    .o(\PWME/n13 [10]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWME/mux0_b11  (
    .i0(\PWME/n12 [11]),
    .i1(freqE[11]),
    .sel(\PWME/n0 ),
    .o(\PWME/n13 [11]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWME/mux0_b12  (
    .i0(\PWME/n12 [12]),
    .i1(freqE[12]),
    .sel(\PWME/n0 ),
    .o(\PWME/n13 [12]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWME/mux0_b13  (
    .i0(\PWME/n12 [13]),
    .i1(freqE[13]),
    .sel(\PWME/n0 ),
    .o(\PWME/n13 [13]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWME/mux0_b14  (
    .i0(\PWME/n12 [14]),
    .i1(freqE[14]),
    .sel(\PWME/n0 ),
    .o(\PWME/n13 [14]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWME/mux0_b15  (
    .i0(\PWME/n12 [15]),
    .i1(freqE[15]),
    .sel(\PWME/n0 ),
    .o(\PWME/n13 [15]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWME/mux0_b16  (
    .i0(\PWME/n12 [16]),
    .i1(freqE[16]),
    .sel(\PWME/n0 ),
    .o(\PWME/n13 [16]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWME/mux0_b17  (
    .i0(\PWME/n12 [17]),
    .i1(freqE[17]),
    .sel(\PWME/n0 ),
    .o(\PWME/n13 [17]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWME/mux0_b18  (
    .i0(\PWME/n12 [18]),
    .i1(freqE[18]),
    .sel(\PWME/n0 ),
    .o(\PWME/n13 [18]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWME/mux0_b19  (
    .i0(\PWME/n12 [19]),
    .i1(freqE[19]),
    .sel(\PWME/n0 ),
    .o(\PWME/n13 [19]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWME/mux0_b2  (
    .i0(\PWME/n12 [2]),
    .i1(freqE[2]),
    .sel(\PWME/n0 ),
    .o(\PWME/n13 [2]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWME/mux0_b20  (
    .i0(\PWME/n12 [20]),
    .i1(freqE[20]),
    .sel(\PWME/n0 ),
    .o(\PWME/n13 [20]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWME/mux0_b21  (
    .i0(\PWME/n12 [21]),
    .i1(freqE[21]),
    .sel(\PWME/n0 ),
    .o(\PWME/n13 [21]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWME/mux0_b22  (
    .i0(\PWME/n12 [22]),
    .i1(freqE[22]),
    .sel(\PWME/n0 ),
    .o(\PWME/n13 [22]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWME/mux0_b23  (
    .i0(\PWME/n12 [23]),
    .i1(freqE[23]),
    .sel(\PWME/n0 ),
    .o(\PWME/n13 [23]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWME/mux0_b24  (
    .i0(\PWME/n12 [24]),
    .i1(freqE[24]),
    .sel(\PWME/n0 ),
    .o(\PWME/n13 [24]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWME/mux0_b25  (
    .i0(\PWME/n12 [25]),
    .i1(freqE[25]),
    .sel(\PWME/n0 ),
    .o(\PWME/n13 [25]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWME/mux0_b26  (
    .i0(\PWME/n12 [26]),
    .i1(freqE[26]),
    .sel(\PWME/n0 ),
    .o(\PWME/n13 [26]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWME/mux0_b3  (
    .i0(\PWME/n12 [3]),
    .i1(freqE[3]),
    .sel(\PWME/n0 ),
    .o(\PWME/n13 [3]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWME/mux0_b4  (
    .i0(\PWME/n12 [4]),
    .i1(freqE[4]),
    .sel(\PWME/n0 ),
    .o(\PWME/n13 [4]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWME/mux0_b5  (
    .i0(\PWME/n12 [5]),
    .i1(freqE[5]),
    .sel(\PWME/n0 ),
    .o(\PWME/n13 [5]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWME/mux0_b6  (
    .i0(\PWME/n12 [6]),
    .i1(freqE[6]),
    .sel(\PWME/n0 ),
    .o(\PWME/n13 [6]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWME/mux0_b7  (
    .i0(\PWME/n12 [7]),
    .i1(freqE[7]),
    .sel(\PWME/n0 ),
    .o(\PWME/n13 [7]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWME/mux0_b8  (
    .i0(\PWME/n12 [8]),
    .i1(freqE[8]),
    .sel(\PWME/n0 ),
    .o(\PWME/n13 [8]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWME/mux0_b9  (
    .i0(\PWME/n12 [9]),
    .i1(freqE[9]),
    .sel(\PWME/n0 ),
    .o(\PWME/n13 [9]));  // src/OnePWM.v(32)
  and \PWME/mux3_b0_sel_is_3  (\PWME/mux3_b0_sel_is_3_o , \PWME/n11 , \PWME/n0 );
  binary_mux_s1_w1 \PWME/mux4_b0  (
    .i0(\PWME/pnumr [0]),
    .i1(1'b0),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n22 [0]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux4_b1  (
    .i0(\PWME/pnumr [1]),
    .i1(1'b0),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n22 [1]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux4_b10  (
    .i0(\PWME/pnumr [10]),
    .i1(1'b0),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n22 [10]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux4_b11  (
    .i0(\PWME/pnumr [11]),
    .i1(1'b0),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n22 [11]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux4_b12  (
    .i0(\PWME/pnumr [12]),
    .i1(1'b0),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n22 [12]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux4_b13  (
    .i0(\PWME/pnumr [13]),
    .i1(1'b0),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n22 [13]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux4_b14  (
    .i0(\PWME/pnumr [14]),
    .i1(1'b0),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n22 [14]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux4_b15  (
    .i0(\PWME/pnumr [15]),
    .i1(1'b0),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n22 [15]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux4_b16  (
    .i0(\PWME/pnumr [16]),
    .i1(1'b0),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n22 [16]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux4_b17  (
    .i0(\PWME/pnumr [17]),
    .i1(1'b0),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n22 [17]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux4_b18  (
    .i0(\PWME/pnumr [18]),
    .i1(1'b0),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n22 [18]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux4_b19  (
    .i0(\PWME/pnumr [19]),
    .i1(1'b0),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n22 [19]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux4_b2  (
    .i0(\PWME/pnumr [2]),
    .i1(1'b0),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n22 [2]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux4_b20  (
    .i0(\PWME/pnumr [20]),
    .i1(1'b0),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n22 [20]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux4_b21  (
    .i0(\PWME/pnumr [21]),
    .i1(1'b0),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n22 [21]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux4_b22  (
    .i0(\PWME/pnumr [22]),
    .i1(1'b0),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n22 [22]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux4_b23  (
    .i0(\PWME/pnumr [23]),
    .i1(1'b0),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n22 [23]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux4_b24  (
    .i0(\PWME/pnumr [24]),
    .i1(1'b0),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n22 [24]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux4_b25  (
    .i0(\PWME/pnumr [25]),
    .i1(1'b0),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n22 [25]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux4_b26  (
    .i0(\PWME/pnumr [26]),
    .i1(1'b0),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n22 [26]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux4_b27  (
    .i0(\PWME/pnumr [27]),
    .i1(1'b0),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n22 [27]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux4_b28  (
    .i0(\PWME/pnumr [28]),
    .i1(1'b0),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n22 [28]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux4_b29  (
    .i0(\PWME/pnumr [29]),
    .i1(1'b0),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n22 [29]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux4_b3  (
    .i0(\PWME/pnumr [3]),
    .i1(1'b0),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n22 [3]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux4_b30  (
    .i0(\PWME/pnumr [30]),
    .i1(1'b0),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n22 [30]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux4_b31  (
    .i0(\PWME/pnumr [31]),
    .i1(1'b0),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n22 [31]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux4_b4  (
    .i0(\PWME/pnumr [4]),
    .i1(1'b0),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n22 [4]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux4_b5  (
    .i0(\PWME/pnumr [5]),
    .i1(1'b0),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n22 [5]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux4_b6  (
    .i0(\PWME/pnumr [6]),
    .i1(1'b0),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n22 [6]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux4_b7  (
    .i0(\PWME/pnumr [7]),
    .i1(1'b0),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n22 [7]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux4_b8  (
    .i0(\PWME/pnumr [8]),
    .i1(1'b0),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n22 [8]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux4_b9  (
    .i0(\PWME/pnumr [9]),
    .i1(1'b0),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n22 [9]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux5_b0  (
    .i0(\PWME/n22 [0]),
    .i1(pnumE[0]),
    .sel(pnumE[32]),
    .o(\PWME/n23 [0]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux5_b1  (
    .i0(\PWME/n22 [1]),
    .i1(pnumE[1]),
    .sel(pnumE[32]),
    .o(\PWME/n23 [1]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux5_b10  (
    .i0(\PWME/n22 [10]),
    .i1(pnumE[10]),
    .sel(pnumE[32]),
    .o(\PWME/n23 [10]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux5_b11  (
    .i0(\PWME/n22 [11]),
    .i1(pnumE[11]),
    .sel(pnumE[32]),
    .o(\PWME/n23 [11]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux5_b12  (
    .i0(\PWME/n22 [12]),
    .i1(pnumE[12]),
    .sel(pnumE[32]),
    .o(\PWME/n23 [12]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux5_b13  (
    .i0(\PWME/n22 [13]),
    .i1(pnumE[13]),
    .sel(pnumE[32]),
    .o(\PWME/n23 [13]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux5_b14  (
    .i0(\PWME/n22 [14]),
    .i1(pnumE[14]),
    .sel(pnumE[32]),
    .o(\PWME/n23 [14]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux5_b15  (
    .i0(\PWME/n22 [15]),
    .i1(pnumE[15]),
    .sel(pnumE[32]),
    .o(\PWME/n23 [15]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux5_b16  (
    .i0(\PWME/n22 [16]),
    .i1(pnumE[16]),
    .sel(pnumE[32]),
    .o(\PWME/n23 [16]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux5_b17  (
    .i0(\PWME/n22 [17]),
    .i1(pnumE[17]),
    .sel(pnumE[32]),
    .o(\PWME/n23 [17]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux5_b18  (
    .i0(\PWME/n22 [18]),
    .i1(pnumE[18]),
    .sel(pnumE[32]),
    .o(\PWME/n23 [18]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux5_b19  (
    .i0(\PWME/n22 [19]),
    .i1(pnumE[19]),
    .sel(pnumE[32]),
    .o(\PWME/n23 [19]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux5_b2  (
    .i0(\PWME/n22 [2]),
    .i1(pnumE[2]),
    .sel(pnumE[32]),
    .o(\PWME/n23 [2]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux5_b20  (
    .i0(\PWME/n22 [20]),
    .i1(pnumE[20]),
    .sel(pnumE[32]),
    .o(\PWME/n23 [20]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux5_b21  (
    .i0(\PWME/n22 [21]),
    .i1(pnumE[21]),
    .sel(pnumE[32]),
    .o(\PWME/n23 [21]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux5_b22  (
    .i0(\PWME/n22 [22]),
    .i1(pnumE[22]),
    .sel(pnumE[32]),
    .o(\PWME/n23 [22]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux5_b23  (
    .i0(\PWME/n22 [23]),
    .i1(pnumE[23]),
    .sel(pnumE[32]),
    .o(\PWME/n23 [23]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux5_b24  (
    .i0(\PWME/n22 [24]),
    .i1(pnumE[24]),
    .sel(pnumE[32]),
    .o(\PWME/n23 [24]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux5_b25  (
    .i0(\PWME/n22 [25]),
    .i1(pnumE[25]),
    .sel(pnumE[32]),
    .o(\PWME/n23 [25]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux5_b26  (
    .i0(\PWME/n22 [26]),
    .i1(pnumE[26]),
    .sel(pnumE[32]),
    .o(\PWME/n23 [26]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux5_b27  (
    .i0(\PWME/n22 [27]),
    .i1(pnumE[27]),
    .sel(pnumE[32]),
    .o(\PWME/n23 [27]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux5_b28  (
    .i0(\PWME/n22 [28]),
    .i1(pnumE[28]),
    .sel(pnumE[32]),
    .o(\PWME/n23 [28]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux5_b29  (
    .i0(\PWME/n22 [29]),
    .i1(pnumE[29]),
    .sel(pnumE[32]),
    .o(\PWME/n23 [29]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux5_b3  (
    .i0(\PWME/n22 [3]),
    .i1(pnumE[3]),
    .sel(pnumE[32]),
    .o(\PWME/n23 [3]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux5_b30  (
    .i0(\PWME/n22 [30]),
    .i1(pnumE[30]),
    .sel(pnumE[32]),
    .o(\PWME/n23 [30]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux5_b31  (
    .i0(\PWME/n22 [31]),
    .i1(pnumE[31]),
    .sel(pnumE[32]),
    .o(\PWME/n23 [31]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux5_b4  (
    .i0(\PWME/n22 [4]),
    .i1(pnumE[4]),
    .sel(pnumE[32]),
    .o(\PWME/n23 [4]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux5_b5  (
    .i0(\PWME/n22 [5]),
    .i1(pnumE[5]),
    .sel(pnumE[32]),
    .o(\PWME/n23 [5]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux5_b6  (
    .i0(\PWME/n22 [6]),
    .i1(pnumE[6]),
    .sel(pnumE[32]),
    .o(\PWME/n23 [6]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux5_b7  (
    .i0(\PWME/n22 [7]),
    .i1(pnumE[7]),
    .sel(pnumE[32]),
    .o(\PWME/n23 [7]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux5_b8  (
    .i0(\PWME/n22 [8]),
    .i1(pnumE[8]),
    .sel(pnumE[32]),
    .o(\PWME/n23 [8]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux5_b9  (
    .i0(\PWME/n22 [9]),
    .i1(pnumE[9]),
    .sel(pnumE[32]),
    .o(\PWME/n23 [9]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWME/mux6_b0  (
    .i0(\PWME/pnumr [0]),
    .i1(\PWME/n26 [0]),
    .sel(\PWME/n25 ),
    .o(\PWME/n27 [0]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWME/mux6_b1  (
    .i0(\PWME/pnumr [1]),
    .i1(\PWME/n26 [1]),
    .sel(\PWME/n25 ),
    .o(\PWME/n27 [1]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWME/mux6_b10  (
    .i0(\PWME/pnumr [10]),
    .i1(\PWME/n26 [10]),
    .sel(\PWME/n25 ),
    .o(\PWME/n27 [10]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWME/mux6_b11  (
    .i0(\PWME/pnumr [11]),
    .i1(\PWME/n26 [11]),
    .sel(\PWME/n25 ),
    .o(\PWME/n27 [11]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWME/mux6_b12  (
    .i0(\PWME/pnumr [12]),
    .i1(\PWME/n26 [12]),
    .sel(\PWME/n25 ),
    .o(\PWME/n27 [12]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWME/mux6_b13  (
    .i0(\PWME/pnumr [13]),
    .i1(\PWME/n26 [13]),
    .sel(\PWME/n25 ),
    .o(\PWME/n27 [13]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWME/mux6_b14  (
    .i0(\PWME/pnumr [14]),
    .i1(\PWME/n26 [14]),
    .sel(\PWME/n25 ),
    .o(\PWME/n27 [14]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWME/mux6_b15  (
    .i0(\PWME/pnumr [15]),
    .i1(\PWME/n26 [15]),
    .sel(\PWME/n25 ),
    .o(\PWME/n27 [15]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWME/mux6_b16  (
    .i0(\PWME/pnumr [16]),
    .i1(\PWME/n26 [16]),
    .sel(\PWME/n25 ),
    .o(\PWME/n27 [16]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWME/mux6_b17  (
    .i0(\PWME/pnumr [17]),
    .i1(\PWME/n26 [17]),
    .sel(\PWME/n25 ),
    .o(\PWME/n27 [17]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWME/mux6_b18  (
    .i0(\PWME/pnumr [18]),
    .i1(\PWME/n26 [18]),
    .sel(\PWME/n25 ),
    .o(\PWME/n27 [18]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWME/mux6_b19  (
    .i0(\PWME/pnumr [19]),
    .i1(\PWME/n26 [19]),
    .sel(\PWME/n25 ),
    .o(\PWME/n27 [19]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWME/mux6_b2  (
    .i0(\PWME/pnumr [2]),
    .i1(\PWME/n26 [2]),
    .sel(\PWME/n25 ),
    .o(\PWME/n27 [2]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWME/mux6_b20  (
    .i0(\PWME/pnumr [20]),
    .i1(\PWME/n26 [20]),
    .sel(\PWME/n25 ),
    .o(\PWME/n27 [20]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWME/mux6_b21  (
    .i0(\PWME/pnumr [21]),
    .i1(\PWME/n26 [21]),
    .sel(\PWME/n25 ),
    .o(\PWME/n27 [21]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWME/mux6_b22  (
    .i0(\PWME/pnumr [22]),
    .i1(\PWME/n26 [22]),
    .sel(\PWME/n25 ),
    .o(\PWME/n27 [22]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWME/mux6_b23  (
    .i0(\PWME/pnumr [23]),
    .i1(\PWME/n26 [23]),
    .sel(\PWME/n25 ),
    .o(\PWME/n27 [23]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWME/mux6_b3  (
    .i0(\PWME/pnumr [3]),
    .i1(\PWME/n26 [3]),
    .sel(\PWME/n25 ),
    .o(\PWME/n27 [3]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWME/mux6_b4  (
    .i0(\PWME/pnumr [4]),
    .i1(\PWME/n26 [4]),
    .sel(\PWME/n25 ),
    .o(\PWME/n27 [4]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWME/mux6_b5  (
    .i0(\PWME/pnumr [5]),
    .i1(\PWME/n26 [5]),
    .sel(\PWME/n25 ),
    .o(\PWME/n27 [5]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWME/mux6_b6  (
    .i0(\PWME/pnumr [6]),
    .i1(\PWME/n26 [6]),
    .sel(\PWME/n25 ),
    .o(\PWME/n27 [6]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWME/mux6_b7  (
    .i0(\PWME/pnumr [7]),
    .i1(\PWME/n26 [7]),
    .sel(\PWME/n25 ),
    .o(\PWME/n27 [7]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWME/mux6_b8  (
    .i0(\PWME/pnumr [8]),
    .i1(\PWME/n26 [8]),
    .sel(\PWME/n25 ),
    .o(\PWME/n27 [8]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWME/mux6_b9  (
    .i0(\PWME/pnumr [9]),
    .i1(\PWME/n26 [9]),
    .sel(\PWME/n25 ),
    .o(\PWME/n27 [9]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWME/mux7_b0  (
    .i0(pnumcntE[0]),
    .i1(\PWME/n27 [0]),
    .sel(\PWME/n24 ),
    .o(\PWME/n29 [0]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux7_b1  (
    .i0(pnumcntE[1]),
    .i1(\PWME/n27 [1]),
    .sel(\PWME/n24 ),
    .o(\PWME/n29 [1]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux7_b10  (
    .i0(pnumcntE[10]),
    .i1(\PWME/n27 [10]),
    .sel(\PWME/n24 ),
    .o(\PWME/n29 [10]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux7_b11  (
    .i0(pnumcntE[11]),
    .i1(\PWME/n27 [11]),
    .sel(\PWME/n24 ),
    .o(\PWME/n29 [11]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux7_b12  (
    .i0(pnumcntE[12]),
    .i1(\PWME/n27 [12]),
    .sel(\PWME/n24 ),
    .o(\PWME/n29 [12]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux7_b13  (
    .i0(pnumcntE[13]),
    .i1(\PWME/n27 [13]),
    .sel(\PWME/n24 ),
    .o(\PWME/n29 [13]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux7_b14  (
    .i0(pnumcntE[14]),
    .i1(\PWME/n27 [14]),
    .sel(\PWME/n24 ),
    .o(\PWME/n29 [14]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux7_b15  (
    .i0(pnumcntE[15]),
    .i1(\PWME/n27 [15]),
    .sel(\PWME/n24 ),
    .o(\PWME/n29 [15]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux7_b16  (
    .i0(pnumcntE[16]),
    .i1(\PWME/n27 [16]),
    .sel(\PWME/n24 ),
    .o(\PWME/n29 [16]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux7_b17  (
    .i0(pnumcntE[17]),
    .i1(\PWME/n27 [17]),
    .sel(\PWME/n24 ),
    .o(\PWME/n29 [17]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux7_b18  (
    .i0(pnumcntE[18]),
    .i1(\PWME/n27 [18]),
    .sel(\PWME/n24 ),
    .o(\PWME/n29 [18]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux7_b19  (
    .i0(pnumcntE[19]),
    .i1(\PWME/n27 [19]),
    .sel(\PWME/n24 ),
    .o(\PWME/n29 [19]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux7_b2  (
    .i0(pnumcntE[2]),
    .i1(\PWME/n27 [2]),
    .sel(\PWME/n24 ),
    .o(\PWME/n29 [2]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux7_b20  (
    .i0(pnumcntE[20]),
    .i1(\PWME/n27 [20]),
    .sel(\PWME/n24 ),
    .o(\PWME/n29 [20]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux7_b21  (
    .i0(pnumcntE[21]),
    .i1(\PWME/n27 [21]),
    .sel(\PWME/n24 ),
    .o(\PWME/n29 [21]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux7_b22  (
    .i0(pnumcntE[22]),
    .i1(\PWME/n27 [22]),
    .sel(\PWME/n24 ),
    .o(\PWME/n29 [22]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux7_b23  (
    .i0(pnumcntE[23]),
    .i1(\PWME/n27 [23]),
    .sel(\PWME/n24 ),
    .o(\PWME/n29 [23]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux7_b3  (
    .i0(pnumcntE[3]),
    .i1(\PWME/n27 [3]),
    .sel(\PWME/n24 ),
    .o(\PWME/n29 [3]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux7_b4  (
    .i0(pnumcntE[4]),
    .i1(\PWME/n27 [4]),
    .sel(\PWME/n24 ),
    .o(\PWME/n29 [4]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux7_b5  (
    .i0(pnumcntE[5]),
    .i1(\PWME/n27 [5]),
    .sel(\PWME/n24 ),
    .o(\PWME/n29 [5]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux7_b6  (
    .i0(pnumcntE[6]),
    .i1(\PWME/n27 [6]),
    .sel(\PWME/n24 ),
    .o(\PWME/n29 [6]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux7_b7  (
    .i0(pnumcntE[7]),
    .i1(\PWME/n27 [7]),
    .sel(\PWME/n24 ),
    .o(\PWME/n29 [7]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux7_b8  (
    .i0(pnumcntE[8]),
    .i1(\PWME/n27 [8]),
    .sel(\PWME/n24 ),
    .o(\PWME/n29 [8]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux7_b9  (
    .i0(pnumcntE[9]),
    .i1(\PWME/n27 [9]),
    .sel(\PWME/n24 ),
    .o(\PWME/n29 [9]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux8_b0  (
    .i0(\PWME/n29 [0]),
    .i1(\PWME/pnumr [0]),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n31 [0]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux8_b1  (
    .i0(\PWME/n29 [1]),
    .i1(\PWME/pnumr [1]),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n31 [1]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux8_b10  (
    .i0(\PWME/n29 [10]),
    .i1(\PWME/pnumr [10]),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n31 [10]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux8_b11  (
    .i0(\PWME/n29 [11]),
    .i1(\PWME/pnumr [11]),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n31 [11]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux8_b12  (
    .i0(\PWME/n29 [12]),
    .i1(\PWME/pnumr [12]),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n31 [12]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux8_b13  (
    .i0(\PWME/n29 [13]),
    .i1(\PWME/pnumr [13]),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n31 [13]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux8_b14  (
    .i0(\PWME/n29 [14]),
    .i1(\PWME/pnumr [14]),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n31 [14]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux8_b15  (
    .i0(\PWME/n29 [15]),
    .i1(\PWME/pnumr [15]),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n31 [15]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux8_b16  (
    .i0(\PWME/n29 [16]),
    .i1(\PWME/pnumr [16]),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n31 [16]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux8_b17  (
    .i0(\PWME/n29 [17]),
    .i1(\PWME/pnumr [17]),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n31 [17]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux8_b18  (
    .i0(\PWME/n29 [18]),
    .i1(\PWME/pnumr [18]),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n31 [18]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux8_b19  (
    .i0(\PWME/n29 [19]),
    .i1(\PWME/pnumr [19]),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n31 [19]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux8_b2  (
    .i0(\PWME/n29 [2]),
    .i1(\PWME/pnumr [2]),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n31 [2]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux8_b20  (
    .i0(\PWME/n29 [20]),
    .i1(\PWME/pnumr [20]),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n31 [20]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux8_b21  (
    .i0(\PWME/n29 [21]),
    .i1(\PWME/pnumr [21]),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n31 [21]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux8_b22  (
    .i0(\PWME/n29 [22]),
    .i1(\PWME/pnumr [22]),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n31 [22]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux8_b23  (
    .i0(\PWME/n29 [23]),
    .i1(\PWME/pnumr [23]),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n31 [23]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux8_b3  (
    .i0(\PWME/n29 [3]),
    .i1(\PWME/pnumr [3]),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n31 [3]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux8_b4  (
    .i0(\PWME/n29 [4]),
    .i1(\PWME/pnumr [4]),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n31 [4]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux8_b5  (
    .i0(\PWME/n29 [5]),
    .i1(\PWME/pnumr [5]),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n31 [5]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux8_b6  (
    .i0(\PWME/n29 [6]),
    .i1(\PWME/pnumr [6]),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n31 [6]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux8_b7  (
    .i0(\PWME/n29 [7]),
    .i1(\PWME/pnumr [7]),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n31 [7]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux8_b8  (
    .i0(\PWME/n29 [8]),
    .i1(\PWME/pnumr [8]),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n31 [8]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWME/mux8_b9  (
    .i0(\PWME/n29 [9]),
    .i1(\PWME/pnumr [9]),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n31 [9]));  // src/OnePWM.v(57)
  not \PWME/n17_inv  (\PWME/n17_neg , \PWME/n17 );
  not \PWME/n25_inv  (\PWME/n25_neg , \PWME/n25 );
  not \PWME/n4_inv  (\PWME/n4_neg , \PWME/n4 );
  not \PWME/n6_inv  (\PWME/n6_neg , \PWME/n6 );
  ne_w24 \PWME/neq0  (
    .i0(pnumcntE),
    .i1(24'b000000000000000000000000),
    .o(\PWME/n25 ));  // src/OnePWM.v(55)
  reg_sr_ss_w1 \PWME/pwm_reg  (
    .clk(clk100m),
    .d(pwm[14]),
    .en(1'b1),
    .reset(~\PWME/u14_sel_is_1_o ),
    .set(\PWME/n18 ),
    .q(\PWME/pwm_keep ));  // src/OnePWM.v(45)
  reg_sr_as_w1 \PWME/reg0_b0  (
    .clk(clk100m),
    .d(\PWME/n13 [0]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [0]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b1  (
    .clk(clk100m),
    .d(\PWME/n13 [1]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [1]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b10  (
    .clk(clk100m),
    .d(\PWME/n13 [10]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [10]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b11  (
    .clk(clk100m),
    .d(\PWME/n13 [11]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [11]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b12  (
    .clk(clk100m),
    .d(\PWME/n13 [12]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [12]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b13  (
    .clk(clk100m),
    .d(\PWME/n13 [13]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [13]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b14  (
    .clk(clk100m),
    .d(\PWME/n13 [14]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [14]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b15  (
    .clk(clk100m),
    .d(\PWME/n13 [15]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [15]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b16  (
    .clk(clk100m),
    .d(\PWME/n13 [16]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [16]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b17  (
    .clk(clk100m),
    .d(\PWME/n13 [17]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [17]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b18  (
    .clk(clk100m),
    .d(\PWME/n13 [18]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [18]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b19  (
    .clk(clk100m),
    .d(\PWME/n13 [19]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [19]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b2  (
    .clk(clk100m),
    .d(\PWME/n13 [2]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [2]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b20  (
    .clk(clk100m),
    .d(\PWME/n13 [20]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [20]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b21  (
    .clk(clk100m),
    .d(\PWME/n13 [21]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [21]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b22  (
    .clk(clk100m),
    .d(\PWME/n13 [22]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [22]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b23  (
    .clk(clk100m),
    .d(\PWME/n13 [23]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [23]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b24  (
    .clk(clk100m),
    .d(\PWME/n13 [24]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [24]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b25  (
    .clk(clk100m),
    .d(\PWME/n13 [25]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [25]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b26  (
    .clk(clk100m),
    .d(\PWME/n13 [26]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [26]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b3  (
    .clk(clk100m),
    .d(\PWME/n13 [3]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [3]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b4  (
    .clk(clk100m),
    .d(\PWME/n13 [4]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [4]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b5  (
    .clk(clk100m),
    .d(\PWME/n13 [5]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [5]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b6  (
    .clk(clk100m),
    .d(\PWME/n13 [6]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [6]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b7  (
    .clk(clk100m),
    .d(\PWME/n13 [7]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [7]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b8  (
    .clk(clk100m),
    .d(\PWME/n13 [8]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [8]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWME/reg0_b9  (
    .clk(clk100m),
    .d(\PWME/n13 [9]),
    .en(1'b1),
    .reset(~\PWME/n11 ),
    .set(1'b0),
    .q(\PWME/FreCnt [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b0  (
    .clk(clk100m),
    .d(freqE[0]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [0]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b1  (
    .clk(clk100m),
    .d(freqE[1]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [1]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b10  (
    .clk(clk100m),
    .d(freqE[10]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [10]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b11  (
    .clk(clk100m),
    .d(freqE[11]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [11]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b12  (
    .clk(clk100m),
    .d(freqE[12]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [12]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b13  (
    .clk(clk100m),
    .d(freqE[13]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [13]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b14  (
    .clk(clk100m),
    .d(freqE[14]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [14]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b15  (
    .clk(clk100m),
    .d(freqE[15]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [15]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b16  (
    .clk(clk100m),
    .d(freqE[16]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [16]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b17  (
    .clk(clk100m),
    .d(freqE[17]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [17]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b18  (
    .clk(clk100m),
    .d(freqE[18]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [18]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b19  (
    .clk(clk100m),
    .d(freqE[19]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [19]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b2  (
    .clk(clk100m),
    .d(freqE[2]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [2]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b20  (
    .clk(clk100m),
    .d(freqE[20]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [20]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b21  (
    .clk(clk100m),
    .d(freqE[21]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [21]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b22  (
    .clk(clk100m),
    .d(freqE[22]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [22]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b23  (
    .clk(clk100m),
    .d(freqE[23]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [23]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b24  (
    .clk(clk100m),
    .d(freqE[24]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [24]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b25  (
    .clk(clk100m),
    .d(freqE[25]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [25]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b26  (
    .clk(clk100m),
    .d(freqE[26]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [26]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b3  (
    .clk(clk100m),
    .d(freqE[3]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [3]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b4  (
    .clk(clk100m),
    .d(freqE[4]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [4]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b5  (
    .clk(clk100m),
    .d(freqE[5]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [5]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b6  (
    .clk(clk100m),
    .d(freqE[6]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [6]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b7  (
    .clk(clk100m),
    .d(freqE[7]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [7]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b8  (
    .clk(clk100m),
    .d(freqE[8]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [8]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg1_b9  (
    .clk(clk100m),
    .d(freqE[9]),
    .en(\PWME/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/FreCntr [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWME/reg2_b0  (
    .clk(clk100m),
    .d(\PWME/n23 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[0]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b1  (
    .clk(clk100m),
    .d(\PWME/n23 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[1]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b10  (
    .clk(clk100m),
    .d(\PWME/n23 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[10]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b11  (
    .clk(clk100m),
    .d(\PWME/n23 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[11]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b12  (
    .clk(clk100m),
    .d(\PWME/n23 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[12]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b13  (
    .clk(clk100m),
    .d(\PWME/n23 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[13]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b14  (
    .clk(clk100m),
    .d(\PWME/n23 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[14]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b15  (
    .clk(clk100m),
    .d(\PWME/n23 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[15]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b16  (
    .clk(clk100m),
    .d(\PWME/n23 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[16]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b17  (
    .clk(clk100m),
    .d(\PWME/n23 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[17]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b18  (
    .clk(clk100m),
    .d(\PWME/n23 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[18]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b19  (
    .clk(clk100m),
    .d(\PWME/n23 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[19]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b2  (
    .clk(clk100m),
    .d(\PWME/n23 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[2]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b20  (
    .clk(clk100m),
    .d(\PWME/n23 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[20]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b21  (
    .clk(clk100m),
    .d(\PWME/n23 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[21]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b22  (
    .clk(clk100m),
    .d(\PWME/n23 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[22]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b23  (
    .clk(clk100m),
    .d(\PWME/n23 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[23]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b24  (
    .clk(clk100m),
    .d(\PWME/n23 [24]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[24]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b25  (
    .clk(clk100m),
    .d(\PWME/n23 [25]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[25]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b26  (
    .clk(clk100m),
    .d(\PWME/n23 [26]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[26]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b27  (
    .clk(clk100m),
    .d(\PWME/n23 [27]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[27]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b28  (
    .clk(clk100m),
    .d(\PWME/n23 [28]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[28]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b29  (
    .clk(clk100m),
    .d(\PWME/n23 [29]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[29]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b3  (
    .clk(clk100m),
    .d(\PWME/n23 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[3]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b30  (
    .clk(clk100m),
    .d(\PWME/n23 [30]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[30]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b31  (
    .clk(clk100m),
    .d(\PWME/n23 [31]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[31]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b4  (
    .clk(clk100m),
    .d(\PWME/n23 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[4]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b5  (
    .clk(clk100m),
    .d(\PWME/n23 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[5]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b6  (
    .clk(clk100m),
    .d(\PWME/n23 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[6]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b7  (
    .clk(clk100m),
    .d(\PWME/n23 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[7]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b8  (
    .clk(clk100m),
    .d(\PWME/n23 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[8]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg2_b9  (
    .clk(clk100m),
    .d(\PWME/n23 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/pnumr[9]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWME/reg3_b0  (
    .clk(clk100m),
    .d(\PWME/n31 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[0]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b1  (
    .clk(clk100m),
    .d(\PWME/n31 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[1]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b10  (
    .clk(clk100m),
    .d(\PWME/n31 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[10]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b11  (
    .clk(clk100m),
    .d(\PWME/n31 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[11]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b12  (
    .clk(clk100m),
    .d(\PWME/n31 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[12]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b13  (
    .clk(clk100m),
    .d(\PWME/n31 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[13]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b14  (
    .clk(clk100m),
    .d(\PWME/n31 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[14]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b15  (
    .clk(clk100m),
    .d(\PWME/n31 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[15]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b16  (
    .clk(clk100m),
    .d(\PWME/n31 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[16]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b17  (
    .clk(clk100m),
    .d(\PWME/n31 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[17]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b18  (
    .clk(clk100m),
    .d(\PWME/n31 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[18]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b19  (
    .clk(clk100m),
    .d(\PWME/n31 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[19]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b2  (
    .clk(clk100m),
    .d(\PWME/n31 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[2]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b20  (
    .clk(clk100m),
    .d(\PWME/n31 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[20]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b21  (
    .clk(clk100m),
    .d(\PWME/n31 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[21]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b22  (
    .clk(clk100m),
    .d(\PWME/n31 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[22]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b23  (
    .clk(clk100m),
    .d(\PWME/n31 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[23]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b3  (
    .clk(clk100m),
    .d(\PWME/n31 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[3]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b4  (
    .clk(clk100m),
    .d(\PWME/n31 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[4]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b5  (
    .clk(clk100m),
    .d(\PWME/n31 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[5]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b6  (
    .clk(clk100m),
    .d(\PWME/n31 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[6]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b7  (
    .clk(clk100m),
    .d(\PWME/n31 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[7]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b8  (
    .clk(clk100m),
    .d(\PWME/n31 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[8]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWME/reg3_b9  (
    .clk(clk100m),
    .d(\PWME/n31 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWME/RemaTxNum[9]_keep ));  // src/OnePWM.v(58)
  reg_ar_ss_w1 \PWME/stopreq_reg  (
    .clk(clk100m),
    .d(\PWME/n1 ),
    .en(1'b1),
    .reset(1'b0),
    .set(pwm_start_stop[14]),
    .q(\PWME/stopreq_keep ));  // src/OnePWM.v(15)
  add_pu27_mu27_o27 \PWME/sub0  (
    .i0(\PWME/FreCnt ),
    .i1(27'b000000000000000000000000001),
    .o(\PWME/n12 [26:0]));  // src/OnePWM.v(32)
  add_pu24_mu24_o24 \PWME/sub1  (
    .i0(pnumcntE),
    .i1(24'b000000000000000000000001),
    .o(\PWME/n26 [23:0]));  // src/OnePWM.v(55)
  AL_MUX \PWME/u10  (
    .i0(1'b0),
    .i1(\PWME/n9 ),
    .sel(n25),
    .o(\PWME/n10 ));  // src/OnePWM.v(26)
  or \PWME/u11  (\PWME/n11 , pwm_state_read[14], pwm_start_stop[30]);  // src/OnePWM.v(30)
  and \PWME/u14_sel_is_1  (\PWME/u14_sel_is_1_o , pwm_state_read[14], \PWME/n17_neg );
  and \PWME/u15  (\PWME/n24 , \PWME/n0 , pwm_state_read[14]);  // src/OnePWM.v(54)
  and \PWME/u17_sel_is_1  (\PWME/u17_sel_is_1_o , \PWME/n24 , \PWME/n25_neg );
  not \PWME/u17_sel_is_1_o_inv  (\PWME/u17_sel_is_1_o_neg , \PWME/u17_sel_is_1_o );
  AL_MUX \PWME/u18  (
    .i0(\PWME/pnumr [31]),
    .i1(dir[14]),
    .sel(\PWME/u18_sel_is_0_o ),
    .o(\PWME/n32 ));
  and \PWME/u18_sel_is_0  (\PWME/u18_sel_is_0_o , \pwm_start_stop[30]_neg , \PWME/u17_sel_is_1_o_neg );
  AL_MUX \PWME/u2  (
    .i0(\PWME/stopreq ),
    .i1(1'b0),
    .sel(\PWME/n0 ),
    .o(\PWME/n1 ));  // src/OnePWM.v(15)
  and \PWME/u5  (\PWME/n4 , \PWME/stopreq , \PWME/n0 );  // src/OnePWM.v(23)
  and \PWME/u6  (\PWME/n6 , \PWME/n5 , \PWME/n0 );  // src/OnePWM.v(25)
  AL_MUX \PWME/u8  (
    .i0(1'b0),
    .i1(pwm_state_read[14]),
    .sel(\PWME/u8_sel_is_0_o ),
    .o(\PWME/n8 ));
  and \PWME/u8_sel_is_0  (\PWME/u8_sel_is_0_o , \PWME/n4_neg , \PWME/n6_neg );
  AL_MUX \PWME/u9  (
    .i0(\PWME/n8 ),
    .i1(1'b1),
    .sel(pwm_start_stop[30]),
    .o(\PWME/n9 ));  // src/OnePWM.v(26)
  reg_ar_as_w1 \PWMF/State_reg  (
    .clk(clk100m),
    .d(\PWMF/n10 ),
    .en(1'b1),
    .reset(~rstn),
    .set(1'b0),
    .q(pwm_state_read[15]));  // src/OnePWM.v(26)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[0]  (
    .i(\PWMF/RemaTxNum[0]_keep ),
    .o(pnumcntF[0]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[10]  (
    .i(\PWMF/RemaTxNum[10]_keep ),
    .o(pnumcntF[10]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[11]  (
    .i(\PWMF/RemaTxNum[11]_keep ),
    .o(pnumcntF[11]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[12]  (
    .i(\PWMF/RemaTxNum[12]_keep ),
    .o(pnumcntF[12]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[13]  (
    .i(\PWMF/RemaTxNum[13]_keep ),
    .o(pnumcntF[13]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[14]  (
    .i(\PWMF/RemaTxNum[14]_keep ),
    .o(pnumcntF[14]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[15]  (
    .i(\PWMF/RemaTxNum[15]_keep ),
    .o(pnumcntF[15]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[16]  (
    .i(\PWMF/RemaTxNum[16]_keep ),
    .o(pnumcntF[16]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[17]  (
    .i(\PWMF/RemaTxNum[17]_keep ),
    .o(pnumcntF[17]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[18]  (
    .i(\PWMF/RemaTxNum[18]_keep ),
    .o(pnumcntF[18]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[19]  (
    .i(\PWMF/RemaTxNum[19]_keep ),
    .o(pnumcntF[19]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[1]  (
    .i(\PWMF/RemaTxNum[1]_keep ),
    .o(pnumcntF[1]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[20]  (
    .i(\PWMF/RemaTxNum[20]_keep ),
    .o(pnumcntF[20]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[21]  (
    .i(\PWMF/RemaTxNum[21]_keep ),
    .o(pnumcntF[21]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[22]  (
    .i(\PWMF/RemaTxNum[22]_keep ),
    .o(pnumcntF[22]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[23]  (
    .i(\PWMF/RemaTxNum[23]_keep ),
    .o(pnumcntF[23]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[2]  (
    .i(\PWMF/RemaTxNum[2]_keep ),
    .o(pnumcntF[2]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[3]  (
    .i(\PWMF/RemaTxNum[3]_keep ),
    .o(pnumcntF[3]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[4]  (
    .i(\PWMF/RemaTxNum[4]_keep ),
    .o(pnumcntF[4]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[5]  (
    .i(\PWMF/RemaTxNum[5]_keep ),
    .o(pnumcntF[5]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[6]  (
    .i(\PWMF/RemaTxNum[6]_keep ),
    .o(pnumcntF[6]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[7]  (
    .i(\PWMF/RemaTxNum[7]_keep ),
    .o(pnumcntF[7]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[8]  (
    .i(\PWMF/RemaTxNum[8]_keep ),
    .o(pnumcntF[8]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_RemaTxNum[9]  (
    .i(\PWMF/RemaTxNum[9]_keep ),
    .o(pnumcntF[9]));  // src/OnePWM.v(8)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_dir  (
    .i(\PWMF/dir_keep ),
    .o(dir[15]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[0]  (
    .i(\PWMF/pnumr[0]_keep ),
    .o(\PWMF/pnumr [0]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[10]  (
    .i(\PWMF/pnumr[10]_keep ),
    .o(\PWMF/pnumr [10]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[11]  (
    .i(\PWMF/pnumr[11]_keep ),
    .o(\PWMF/pnumr [11]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[12]  (
    .i(\PWMF/pnumr[12]_keep ),
    .o(\PWMF/pnumr [12]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[13]  (
    .i(\PWMF/pnumr[13]_keep ),
    .o(\PWMF/pnumr [13]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[14]  (
    .i(\PWMF/pnumr[14]_keep ),
    .o(\PWMF/pnumr [14]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[15]  (
    .i(\PWMF/pnumr[15]_keep ),
    .o(\PWMF/pnumr [15]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[16]  (
    .i(\PWMF/pnumr[16]_keep ),
    .o(\PWMF/pnumr [16]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[17]  (
    .i(\PWMF/pnumr[17]_keep ),
    .o(\PWMF/pnumr [17]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[18]  (
    .i(\PWMF/pnumr[18]_keep ),
    .o(\PWMF/pnumr [18]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[19]  (
    .i(\PWMF/pnumr[19]_keep ),
    .o(\PWMF/pnumr [19]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[1]  (
    .i(\PWMF/pnumr[1]_keep ),
    .o(\PWMF/pnumr [1]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[20]  (
    .i(\PWMF/pnumr[20]_keep ),
    .o(\PWMF/pnumr [20]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[21]  (
    .i(\PWMF/pnumr[21]_keep ),
    .o(\PWMF/pnumr [21]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[22]  (
    .i(\PWMF/pnumr[22]_keep ),
    .o(\PWMF/pnumr [22]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[23]  (
    .i(\PWMF/pnumr[23]_keep ),
    .o(\PWMF/pnumr [23]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[24]  (
    .i(\PWMF/pnumr[24]_keep ),
    .o(\PWMF/pnumr [24]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[25]  (
    .i(\PWMF/pnumr[25]_keep ),
    .o(\PWMF/pnumr [25]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[26]  (
    .i(\PWMF/pnumr[26]_keep ),
    .o(\PWMF/pnumr [26]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[27]  (
    .i(\PWMF/pnumr[27]_keep ),
    .o(\PWMF/pnumr [27]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[28]  (
    .i(\PWMF/pnumr[28]_keep ),
    .o(\PWMF/pnumr [28]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[29]  (
    .i(\PWMF/pnumr[29]_keep ),
    .o(\PWMF/pnumr [29]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[2]  (
    .i(\PWMF/pnumr[2]_keep ),
    .o(\PWMF/pnumr [2]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[30]  (
    .i(\PWMF/pnumr[30]_keep ),
    .o(\PWMF/pnumr [30]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[31]  (
    .i(\PWMF/pnumr[31]_keep ),
    .o(\PWMF/pnumr [31]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[3]  (
    .i(\PWMF/pnumr[3]_keep ),
    .o(\PWMF/pnumr [3]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[4]  (
    .i(\PWMF/pnumr[4]_keep ),
    .o(\PWMF/pnumr [4]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[5]  (
    .i(\PWMF/pnumr[5]_keep ),
    .o(\PWMF/pnumr [5]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[6]  (
    .i(\PWMF/pnumr[6]_keep ),
    .o(\PWMF/pnumr [6]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[7]  (
    .i(\PWMF/pnumr[7]_keep ),
    .o(\PWMF/pnumr [7]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[8]  (
    .i(\PWMF/pnumr[8]_keep ),
    .o(\PWMF/pnumr [8]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pnumr[9]  (
    .i(\PWMF/pnumr[9]_keep ),
    .o(\PWMF/pnumr [9]));  // src/OnePWM.v(47)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_pwm  (
    .i(\PWMF/pwm_keep ),
    .o(pwm[15]));  // src/OnePWM.v(9)
  AL_BUFKEEP #(
    .KEEP("OUT"))
    \PWMF/_bufkeep_stopreq  (
    .i(\PWMF/stopreq_keep ),
    .o(\PWMF/stopreq ));  // src/OnePWM.v(14)
  reg_ar_as_w1 \PWMF/dir_reg  (
    .clk(clk100m),
    .d(\PWMF/n32 ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/dir_keep ));  // src/OnePWM.v(58)
  eq_w27 \PWMF/eq0  (
    .i0(\PWMF/FreCnt ),
    .i1(27'b000000000000000000000000000),
    .o(\PWMF/n0 ));  // src/OnePWM.v(15)
  eq_w24 \PWMF/eq1  (
    .i0(pnumcntF),
    .i1(24'b000000000000000000000001),
    .o(\PWMF/n5 ));  // src/OnePWM.v(25)
  eq_w27 \PWMF/eq2  (
    .i0(\PWMF/FreCnt ),
    .i1({1'b0,\PWMF/FreCntr [26:1]}),
    .o(\PWMF/n17 ));  // src/OnePWM.v(41)
  eq_w27 \PWMF/eq3  (
    .i0(\PWMF/FreCnt ),
    .i1(\PWMF/FreCntr ),
    .o(\PWMF/n18 ));  // src/OnePWM.v(43)
  binary_mux_s1_w1 \PWMF/mux0_b0  (
    .i0(\PWMF/n12 [0]),
    .i1(freqF[0]),
    .sel(\PWMF/n0 ),
    .o(\PWMF/n13 [0]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMF/mux0_b1  (
    .i0(\PWMF/n12 [1]),
    .i1(freqF[1]),
    .sel(\PWMF/n0 ),
    .o(\PWMF/n13 [1]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMF/mux0_b10  (
    .i0(\PWMF/n12 [10]),
    .i1(freqF[10]),
    .sel(\PWMF/n0 ),
    .o(\PWMF/n13 [10]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMF/mux0_b11  (
    .i0(\PWMF/n12 [11]),
    .i1(freqF[11]),
    .sel(\PWMF/n0 ),
    .o(\PWMF/n13 [11]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMF/mux0_b12  (
    .i0(\PWMF/n12 [12]),
    .i1(freqF[12]),
    .sel(\PWMF/n0 ),
    .o(\PWMF/n13 [12]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMF/mux0_b13  (
    .i0(\PWMF/n12 [13]),
    .i1(freqF[13]),
    .sel(\PWMF/n0 ),
    .o(\PWMF/n13 [13]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMF/mux0_b14  (
    .i0(\PWMF/n12 [14]),
    .i1(freqF[14]),
    .sel(\PWMF/n0 ),
    .o(\PWMF/n13 [14]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMF/mux0_b15  (
    .i0(\PWMF/n12 [15]),
    .i1(freqF[15]),
    .sel(\PWMF/n0 ),
    .o(\PWMF/n13 [15]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMF/mux0_b16  (
    .i0(\PWMF/n12 [16]),
    .i1(freqF[16]),
    .sel(\PWMF/n0 ),
    .o(\PWMF/n13 [16]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMF/mux0_b17  (
    .i0(\PWMF/n12 [17]),
    .i1(freqF[17]),
    .sel(\PWMF/n0 ),
    .o(\PWMF/n13 [17]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMF/mux0_b18  (
    .i0(\PWMF/n12 [18]),
    .i1(freqF[18]),
    .sel(\PWMF/n0 ),
    .o(\PWMF/n13 [18]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMF/mux0_b19  (
    .i0(\PWMF/n12 [19]),
    .i1(freqF[19]),
    .sel(\PWMF/n0 ),
    .o(\PWMF/n13 [19]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMF/mux0_b2  (
    .i0(\PWMF/n12 [2]),
    .i1(freqF[2]),
    .sel(\PWMF/n0 ),
    .o(\PWMF/n13 [2]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMF/mux0_b20  (
    .i0(\PWMF/n12 [20]),
    .i1(freqF[20]),
    .sel(\PWMF/n0 ),
    .o(\PWMF/n13 [20]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMF/mux0_b21  (
    .i0(\PWMF/n12 [21]),
    .i1(freqF[21]),
    .sel(\PWMF/n0 ),
    .o(\PWMF/n13 [21]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMF/mux0_b22  (
    .i0(\PWMF/n12 [22]),
    .i1(freqF[22]),
    .sel(\PWMF/n0 ),
    .o(\PWMF/n13 [22]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMF/mux0_b23  (
    .i0(\PWMF/n12 [23]),
    .i1(freqF[23]),
    .sel(\PWMF/n0 ),
    .o(\PWMF/n13 [23]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMF/mux0_b24  (
    .i0(\PWMF/n12 [24]),
    .i1(freqF[24]),
    .sel(\PWMF/n0 ),
    .o(\PWMF/n13 [24]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMF/mux0_b25  (
    .i0(\PWMF/n12 [25]),
    .i1(freqF[25]),
    .sel(\PWMF/n0 ),
    .o(\PWMF/n13 [25]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMF/mux0_b26  (
    .i0(\PWMF/n12 [26]),
    .i1(freqF[26]),
    .sel(\PWMF/n0 ),
    .o(\PWMF/n13 [26]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMF/mux0_b3  (
    .i0(\PWMF/n12 [3]),
    .i1(freqF[3]),
    .sel(\PWMF/n0 ),
    .o(\PWMF/n13 [3]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMF/mux0_b4  (
    .i0(\PWMF/n12 [4]),
    .i1(freqF[4]),
    .sel(\PWMF/n0 ),
    .o(\PWMF/n13 [4]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMF/mux0_b5  (
    .i0(\PWMF/n12 [5]),
    .i1(freqF[5]),
    .sel(\PWMF/n0 ),
    .o(\PWMF/n13 [5]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMF/mux0_b6  (
    .i0(\PWMF/n12 [6]),
    .i1(freqF[6]),
    .sel(\PWMF/n0 ),
    .o(\PWMF/n13 [6]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMF/mux0_b7  (
    .i0(\PWMF/n12 [7]),
    .i1(freqF[7]),
    .sel(\PWMF/n0 ),
    .o(\PWMF/n13 [7]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMF/mux0_b8  (
    .i0(\PWMF/n12 [8]),
    .i1(freqF[8]),
    .sel(\PWMF/n0 ),
    .o(\PWMF/n13 [8]));  // src/OnePWM.v(32)
  binary_mux_s1_w1 \PWMF/mux0_b9  (
    .i0(\PWMF/n12 [9]),
    .i1(freqF[9]),
    .sel(\PWMF/n0 ),
    .o(\PWMF/n13 [9]));  // src/OnePWM.v(32)
  and \PWMF/mux3_b0_sel_is_3  (\PWMF/mux3_b0_sel_is_3_o , \PWMF/n11 , \PWMF/n0 );
  binary_mux_s1_w1 \PWMF/mux4_b0  (
    .i0(\PWMF/pnumr [0]),
    .i1(1'b0),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n22 [0]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux4_b1  (
    .i0(\PWMF/pnumr [1]),
    .i1(1'b0),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n22 [1]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux4_b10  (
    .i0(\PWMF/pnumr [10]),
    .i1(1'b0),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n22 [10]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux4_b11  (
    .i0(\PWMF/pnumr [11]),
    .i1(1'b0),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n22 [11]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux4_b12  (
    .i0(\PWMF/pnumr [12]),
    .i1(1'b0),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n22 [12]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux4_b13  (
    .i0(\PWMF/pnumr [13]),
    .i1(1'b0),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n22 [13]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux4_b14  (
    .i0(\PWMF/pnumr [14]),
    .i1(1'b0),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n22 [14]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux4_b15  (
    .i0(\PWMF/pnumr [15]),
    .i1(1'b0),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n22 [15]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux4_b16  (
    .i0(\PWMF/pnumr [16]),
    .i1(1'b0),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n22 [16]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux4_b17  (
    .i0(\PWMF/pnumr [17]),
    .i1(1'b0),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n22 [17]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux4_b18  (
    .i0(\PWMF/pnumr [18]),
    .i1(1'b0),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n22 [18]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux4_b19  (
    .i0(\PWMF/pnumr [19]),
    .i1(1'b0),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n22 [19]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux4_b2  (
    .i0(\PWMF/pnumr [2]),
    .i1(1'b0),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n22 [2]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux4_b20  (
    .i0(\PWMF/pnumr [20]),
    .i1(1'b0),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n22 [20]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux4_b21  (
    .i0(\PWMF/pnumr [21]),
    .i1(1'b0),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n22 [21]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux4_b22  (
    .i0(\PWMF/pnumr [22]),
    .i1(1'b0),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n22 [22]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux4_b23  (
    .i0(\PWMF/pnumr [23]),
    .i1(1'b0),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n22 [23]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux4_b24  (
    .i0(\PWMF/pnumr [24]),
    .i1(1'b0),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n22 [24]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux4_b25  (
    .i0(\PWMF/pnumr [25]),
    .i1(1'b0),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n22 [25]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux4_b26  (
    .i0(\PWMF/pnumr [26]),
    .i1(1'b0),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n22 [26]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux4_b27  (
    .i0(\PWMF/pnumr [27]),
    .i1(1'b0),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n22 [27]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux4_b28  (
    .i0(\PWMF/pnumr [28]),
    .i1(1'b0),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n22 [28]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux4_b29  (
    .i0(\PWMF/pnumr [29]),
    .i1(1'b0),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n22 [29]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux4_b3  (
    .i0(\PWMF/pnumr [3]),
    .i1(1'b0),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n22 [3]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux4_b30  (
    .i0(\PWMF/pnumr [30]),
    .i1(1'b0),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n22 [30]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux4_b31  (
    .i0(\PWMF/pnumr [31]),
    .i1(1'b0),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n22 [31]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux4_b4  (
    .i0(\PWMF/pnumr [4]),
    .i1(1'b0),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n22 [4]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux4_b5  (
    .i0(\PWMF/pnumr [5]),
    .i1(1'b0),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n22 [5]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux4_b6  (
    .i0(\PWMF/pnumr [6]),
    .i1(1'b0),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n22 [6]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux4_b7  (
    .i0(\PWMF/pnumr [7]),
    .i1(1'b0),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n22 [7]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux4_b8  (
    .i0(\PWMF/pnumr [8]),
    .i1(1'b0),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n22 [8]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux4_b9  (
    .i0(\PWMF/pnumr [9]),
    .i1(1'b0),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n22 [9]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux5_b0  (
    .i0(\PWMF/n22 [0]),
    .i1(pnumF[0]),
    .sel(pnumF[32]),
    .o(\PWMF/n23 [0]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux5_b1  (
    .i0(\PWMF/n22 [1]),
    .i1(pnumF[1]),
    .sel(pnumF[32]),
    .o(\PWMF/n23 [1]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux5_b10  (
    .i0(\PWMF/n22 [10]),
    .i1(pnumF[10]),
    .sel(pnumF[32]),
    .o(\PWMF/n23 [10]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux5_b11  (
    .i0(\PWMF/n22 [11]),
    .i1(pnumF[11]),
    .sel(pnumF[32]),
    .o(\PWMF/n23 [11]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux5_b12  (
    .i0(\PWMF/n22 [12]),
    .i1(pnumF[12]),
    .sel(pnumF[32]),
    .o(\PWMF/n23 [12]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux5_b13  (
    .i0(\PWMF/n22 [13]),
    .i1(pnumF[13]),
    .sel(pnumF[32]),
    .o(\PWMF/n23 [13]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux5_b14  (
    .i0(\PWMF/n22 [14]),
    .i1(pnumF[14]),
    .sel(pnumF[32]),
    .o(\PWMF/n23 [14]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux5_b15  (
    .i0(\PWMF/n22 [15]),
    .i1(pnumF[15]),
    .sel(pnumF[32]),
    .o(\PWMF/n23 [15]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux5_b16  (
    .i0(\PWMF/n22 [16]),
    .i1(pnumF[16]),
    .sel(pnumF[32]),
    .o(\PWMF/n23 [16]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux5_b17  (
    .i0(\PWMF/n22 [17]),
    .i1(pnumF[17]),
    .sel(pnumF[32]),
    .o(\PWMF/n23 [17]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux5_b18  (
    .i0(\PWMF/n22 [18]),
    .i1(pnumF[18]),
    .sel(pnumF[32]),
    .o(\PWMF/n23 [18]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux5_b19  (
    .i0(\PWMF/n22 [19]),
    .i1(pnumF[19]),
    .sel(pnumF[32]),
    .o(\PWMF/n23 [19]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux5_b2  (
    .i0(\PWMF/n22 [2]),
    .i1(pnumF[2]),
    .sel(pnumF[32]),
    .o(\PWMF/n23 [2]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux5_b20  (
    .i0(\PWMF/n22 [20]),
    .i1(pnumF[20]),
    .sel(pnumF[32]),
    .o(\PWMF/n23 [20]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux5_b21  (
    .i0(\PWMF/n22 [21]),
    .i1(pnumF[21]),
    .sel(pnumF[32]),
    .o(\PWMF/n23 [21]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux5_b22  (
    .i0(\PWMF/n22 [22]),
    .i1(pnumF[22]),
    .sel(pnumF[32]),
    .o(\PWMF/n23 [22]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux5_b23  (
    .i0(\PWMF/n22 [23]),
    .i1(pnumF[23]),
    .sel(pnumF[32]),
    .o(\PWMF/n23 [23]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux5_b24  (
    .i0(\PWMF/n22 [24]),
    .i1(pnumF[24]),
    .sel(pnumF[32]),
    .o(\PWMF/n23 [24]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux5_b25  (
    .i0(\PWMF/n22 [25]),
    .i1(pnumF[25]),
    .sel(pnumF[32]),
    .o(\PWMF/n23 [25]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux5_b26  (
    .i0(\PWMF/n22 [26]),
    .i1(pnumF[26]),
    .sel(pnumF[32]),
    .o(\PWMF/n23 [26]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux5_b27  (
    .i0(\PWMF/n22 [27]),
    .i1(pnumF[27]),
    .sel(pnumF[32]),
    .o(\PWMF/n23 [27]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux5_b28  (
    .i0(\PWMF/n22 [28]),
    .i1(pnumF[28]),
    .sel(pnumF[32]),
    .o(\PWMF/n23 [28]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux5_b29  (
    .i0(\PWMF/n22 [29]),
    .i1(pnumF[29]),
    .sel(pnumF[32]),
    .o(\PWMF/n23 [29]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux5_b3  (
    .i0(\PWMF/n22 [3]),
    .i1(pnumF[3]),
    .sel(pnumF[32]),
    .o(\PWMF/n23 [3]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux5_b30  (
    .i0(\PWMF/n22 [30]),
    .i1(pnumF[30]),
    .sel(pnumF[32]),
    .o(\PWMF/n23 [30]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux5_b31  (
    .i0(\PWMF/n22 [31]),
    .i1(pnumF[31]),
    .sel(pnumF[32]),
    .o(\PWMF/n23 [31]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux5_b4  (
    .i0(\PWMF/n22 [4]),
    .i1(pnumF[4]),
    .sel(pnumF[32]),
    .o(\PWMF/n23 [4]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux5_b5  (
    .i0(\PWMF/n22 [5]),
    .i1(pnumF[5]),
    .sel(pnumF[32]),
    .o(\PWMF/n23 [5]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux5_b6  (
    .i0(\PWMF/n22 [6]),
    .i1(pnumF[6]),
    .sel(pnumF[32]),
    .o(\PWMF/n23 [6]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux5_b7  (
    .i0(\PWMF/n22 [7]),
    .i1(pnumF[7]),
    .sel(pnumF[32]),
    .o(\PWMF/n23 [7]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux5_b8  (
    .i0(\PWMF/n22 [8]),
    .i1(pnumF[8]),
    .sel(pnumF[32]),
    .o(\PWMF/n23 [8]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux5_b9  (
    .i0(\PWMF/n22 [9]),
    .i1(pnumF[9]),
    .sel(pnumF[32]),
    .o(\PWMF/n23 [9]));  // src/OnePWM.v(48)
  binary_mux_s1_w1 \PWMF/mux6_b0  (
    .i0(\PWMF/pnumr [0]),
    .i1(\PWMF/n26 [0]),
    .sel(\PWMF/n25 ),
    .o(\PWMF/n27 [0]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMF/mux6_b1  (
    .i0(\PWMF/pnumr [1]),
    .i1(\PWMF/n26 [1]),
    .sel(\PWMF/n25 ),
    .o(\PWMF/n27 [1]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMF/mux6_b10  (
    .i0(\PWMF/pnumr [10]),
    .i1(\PWMF/n26 [10]),
    .sel(\PWMF/n25 ),
    .o(\PWMF/n27 [10]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMF/mux6_b11  (
    .i0(\PWMF/pnumr [11]),
    .i1(\PWMF/n26 [11]),
    .sel(\PWMF/n25 ),
    .o(\PWMF/n27 [11]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMF/mux6_b12  (
    .i0(\PWMF/pnumr [12]),
    .i1(\PWMF/n26 [12]),
    .sel(\PWMF/n25 ),
    .o(\PWMF/n27 [12]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMF/mux6_b13  (
    .i0(\PWMF/pnumr [13]),
    .i1(\PWMF/n26 [13]),
    .sel(\PWMF/n25 ),
    .o(\PWMF/n27 [13]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMF/mux6_b14  (
    .i0(\PWMF/pnumr [14]),
    .i1(\PWMF/n26 [14]),
    .sel(\PWMF/n25 ),
    .o(\PWMF/n27 [14]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMF/mux6_b15  (
    .i0(\PWMF/pnumr [15]),
    .i1(\PWMF/n26 [15]),
    .sel(\PWMF/n25 ),
    .o(\PWMF/n27 [15]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMF/mux6_b16  (
    .i0(\PWMF/pnumr [16]),
    .i1(\PWMF/n26 [16]),
    .sel(\PWMF/n25 ),
    .o(\PWMF/n27 [16]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMF/mux6_b17  (
    .i0(\PWMF/pnumr [17]),
    .i1(\PWMF/n26 [17]),
    .sel(\PWMF/n25 ),
    .o(\PWMF/n27 [17]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMF/mux6_b18  (
    .i0(\PWMF/pnumr [18]),
    .i1(\PWMF/n26 [18]),
    .sel(\PWMF/n25 ),
    .o(\PWMF/n27 [18]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMF/mux6_b19  (
    .i0(\PWMF/pnumr [19]),
    .i1(\PWMF/n26 [19]),
    .sel(\PWMF/n25 ),
    .o(\PWMF/n27 [19]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMF/mux6_b2  (
    .i0(\PWMF/pnumr [2]),
    .i1(\PWMF/n26 [2]),
    .sel(\PWMF/n25 ),
    .o(\PWMF/n27 [2]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMF/mux6_b20  (
    .i0(\PWMF/pnumr [20]),
    .i1(\PWMF/n26 [20]),
    .sel(\PWMF/n25 ),
    .o(\PWMF/n27 [20]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMF/mux6_b21  (
    .i0(\PWMF/pnumr [21]),
    .i1(\PWMF/n26 [21]),
    .sel(\PWMF/n25 ),
    .o(\PWMF/n27 [21]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMF/mux6_b22  (
    .i0(\PWMF/pnumr [22]),
    .i1(\PWMF/n26 [22]),
    .sel(\PWMF/n25 ),
    .o(\PWMF/n27 [22]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMF/mux6_b23  (
    .i0(\PWMF/pnumr [23]),
    .i1(\PWMF/n26 [23]),
    .sel(\PWMF/n25 ),
    .o(\PWMF/n27 [23]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMF/mux6_b3  (
    .i0(\PWMF/pnumr [3]),
    .i1(\PWMF/n26 [3]),
    .sel(\PWMF/n25 ),
    .o(\PWMF/n27 [3]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMF/mux6_b4  (
    .i0(\PWMF/pnumr [4]),
    .i1(\PWMF/n26 [4]),
    .sel(\PWMF/n25 ),
    .o(\PWMF/n27 [4]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMF/mux6_b5  (
    .i0(\PWMF/pnumr [5]),
    .i1(\PWMF/n26 [5]),
    .sel(\PWMF/n25 ),
    .o(\PWMF/n27 [5]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMF/mux6_b6  (
    .i0(\PWMF/pnumr [6]),
    .i1(\PWMF/n26 [6]),
    .sel(\PWMF/n25 ),
    .o(\PWMF/n27 [6]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMF/mux6_b7  (
    .i0(\PWMF/pnumr [7]),
    .i1(\PWMF/n26 [7]),
    .sel(\PWMF/n25 ),
    .o(\PWMF/n27 [7]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMF/mux6_b8  (
    .i0(\PWMF/pnumr [8]),
    .i1(\PWMF/n26 [8]),
    .sel(\PWMF/n25 ),
    .o(\PWMF/n27 [8]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMF/mux6_b9  (
    .i0(\PWMF/pnumr [9]),
    .i1(\PWMF/n26 [9]),
    .sel(\PWMF/n25 ),
    .o(\PWMF/n27 [9]));  // src/OnePWM.v(56)
  binary_mux_s1_w1 \PWMF/mux7_b0  (
    .i0(pnumcntF[0]),
    .i1(\PWMF/n27 [0]),
    .sel(\PWMF/n24 ),
    .o(\PWMF/n29 [0]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux7_b1  (
    .i0(pnumcntF[1]),
    .i1(\PWMF/n27 [1]),
    .sel(\PWMF/n24 ),
    .o(\PWMF/n29 [1]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux7_b10  (
    .i0(pnumcntF[10]),
    .i1(\PWMF/n27 [10]),
    .sel(\PWMF/n24 ),
    .o(\PWMF/n29 [10]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux7_b11  (
    .i0(pnumcntF[11]),
    .i1(\PWMF/n27 [11]),
    .sel(\PWMF/n24 ),
    .o(\PWMF/n29 [11]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux7_b12  (
    .i0(pnumcntF[12]),
    .i1(\PWMF/n27 [12]),
    .sel(\PWMF/n24 ),
    .o(\PWMF/n29 [12]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux7_b13  (
    .i0(pnumcntF[13]),
    .i1(\PWMF/n27 [13]),
    .sel(\PWMF/n24 ),
    .o(\PWMF/n29 [13]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux7_b14  (
    .i0(pnumcntF[14]),
    .i1(\PWMF/n27 [14]),
    .sel(\PWMF/n24 ),
    .o(\PWMF/n29 [14]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux7_b15  (
    .i0(pnumcntF[15]),
    .i1(\PWMF/n27 [15]),
    .sel(\PWMF/n24 ),
    .o(\PWMF/n29 [15]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux7_b16  (
    .i0(pnumcntF[16]),
    .i1(\PWMF/n27 [16]),
    .sel(\PWMF/n24 ),
    .o(\PWMF/n29 [16]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux7_b17  (
    .i0(pnumcntF[17]),
    .i1(\PWMF/n27 [17]),
    .sel(\PWMF/n24 ),
    .o(\PWMF/n29 [17]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux7_b18  (
    .i0(pnumcntF[18]),
    .i1(\PWMF/n27 [18]),
    .sel(\PWMF/n24 ),
    .o(\PWMF/n29 [18]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux7_b19  (
    .i0(pnumcntF[19]),
    .i1(\PWMF/n27 [19]),
    .sel(\PWMF/n24 ),
    .o(\PWMF/n29 [19]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux7_b2  (
    .i0(pnumcntF[2]),
    .i1(\PWMF/n27 [2]),
    .sel(\PWMF/n24 ),
    .o(\PWMF/n29 [2]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux7_b20  (
    .i0(pnumcntF[20]),
    .i1(\PWMF/n27 [20]),
    .sel(\PWMF/n24 ),
    .o(\PWMF/n29 [20]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux7_b21  (
    .i0(pnumcntF[21]),
    .i1(\PWMF/n27 [21]),
    .sel(\PWMF/n24 ),
    .o(\PWMF/n29 [21]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux7_b22  (
    .i0(pnumcntF[22]),
    .i1(\PWMF/n27 [22]),
    .sel(\PWMF/n24 ),
    .o(\PWMF/n29 [22]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux7_b23  (
    .i0(pnumcntF[23]),
    .i1(\PWMF/n27 [23]),
    .sel(\PWMF/n24 ),
    .o(\PWMF/n29 [23]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux7_b3  (
    .i0(pnumcntF[3]),
    .i1(\PWMF/n27 [3]),
    .sel(\PWMF/n24 ),
    .o(\PWMF/n29 [3]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux7_b4  (
    .i0(pnumcntF[4]),
    .i1(\PWMF/n27 [4]),
    .sel(\PWMF/n24 ),
    .o(\PWMF/n29 [4]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux7_b5  (
    .i0(pnumcntF[5]),
    .i1(\PWMF/n27 [5]),
    .sel(\PWMF/n24 ),
    .o(\PWMF/n29 [5]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux7_b6  (
    .i0(pnumcntF[6]),
    .i1(\PWMF/n27 [6]),
    .sel(\PWMF/n24 ),
    .o(\PWMF/n29 [6]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux7_b7  (
    .i0(pnumcntF[7]),
    .i1(\PWMF/n27 [7]),
    .sel(\PWMF/n24 ),
    .o(\PWMF/n29 [7]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux7_b8  (
    .i0(pnumcntF[8]),
    .i1(\PWMF/n27 [8]),
    .sel(\PWMF/n24 ),
    .o(\PWMF/n29 [8]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux7_b9  (
    .i0(pnumcntF[9]),
    .i1(\PWMF/n27 [9]),
    .sel(\PWMF/n24 ),
    .o(\PWMF/n29 [9]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux8_b0  (
    .i0(\PWMF/n29 [0]),
    .i1(\PWMF/pnumr [0]),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n31 [0]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux8_b1  (
    .i0(\PWMF/n29 [1]),
    .i1(\PWMF/pnumr [1]),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n31 [1]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux8_b10  (
    .i0(\PWMF/n29 [10]),
    .i1(\PWMF/pnumr [10]),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n31 [10]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux8_b11  (
    .i0(\PWMF/n29 [11]),
    .i1(\PWMF/pnumr [11]),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n31 [11]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux8_b12  (
    .i0(\PWMF/n29 [12]),
    .i1(\PWMF/pnumr [12]),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n31 [12]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux8_b13  (
    .i0(\PWMF/n29 [13]),
    .i1(\PWMF/pnumr [13]),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n31 [13]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux8_b14  (
    .i0(\PWMF/n29 [14]),
    .i1(\PWMF/pnumr [14]),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n31 [14]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux8_b15  (
    .i0(\PWMF/n29 [15]),
    .i1(\PWMF/pnumr [15]),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n31 [15]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux8_b16  (
    .i0(\PWMF/n29 [16]),
    .i1(\PWMF/pnumr [16]),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n31 [16]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux8_b17  (
    .i0(\PWMF/n29 [17]),
    .i1(\PWMF/pnumr [17]),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n31 [17]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux8_b18  (
    .i0(\PWMF/n29 [18]),
    .i1(\PWMF/pnumr [18]),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n31 [18]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux8_b19  (
    .i0(\PWMF/n29 [19]),
    .i1(\PWMF/pnumr [19]),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n31 [19]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux8_b2  (
    .i0(\PWMF/n29 [2]),
    .i1(\PWMF/pnumr [2]),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n31 [2]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux8_b20  (
    .i0(\PWMF/n29 [20]),
    .i1(\PWMF/pnumr [20]),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n31 [20]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux8_b21  (
    .i0(\PWMF/n29 [21]),
    .i1(\PWMF/pnumr [21]),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n31 [21]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux8_b22  (
    .i0(\PWMF/n29 [22]),
    .i1(\PWMF/pnumr [22]),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n31 [22]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux8_b23  (
    .i0(\PWMF/n29 [23]),
    .i1(\PWMF/pnumr [23]),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n31 [23]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux8_b3  (
    .i0(\PWMF/n29 [3]),
    .i1(\PWMF/pnumr [3]),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n31 [3]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux8_b4  (
    .i0(\PWMF/n29 [4]),
    .i1(\PWMF/pnumr [4]),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n31 [4]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux8_b5  (
    .i0(\PWMF/n29 [5]),
    .i1(\PWMF/pnumr [5]),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n31 [5]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux8_b6  (
    .i0(\PWMF/n29 [6]),
    .i1(\PWMF/pnumr [6]),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n31 [6]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux8_b7  (
    .i0(\PWMF/n29 [7]),
    .i1(\PWMF/pnumr [7]),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n31 [7]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux8_b8  (
    .i0(\PWMF/n29 [8]),
    .i1(\PWMF/pnumr [8]),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n31 [8]));  // src/OnePWM.v(57)
  binary_mux_s1_w1 \PWMF/mux8_b9  (
    .i0(\PWMF/n29 [9]),
    .i1(\PWMF/pnumr [9]),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n31 [9]));  // src/OnePWM.v(57)
  not \PWMF/n17_inv  (\PWMF/n17_neg , \PWMF/n17 );
  not \PWMF/n25_inv  (\PWMF/n25_neg , \PWMF/n25 );
  not \PWMF/n4_inv  (\PWMF/n4_neg , \PWMF/n4 );
  not \PWMF/n6_inv  (\PWMF/n6_neg , \PWMF/n6 );
  ne_w24 \PWMF/neq0  (
    .i0(pnumcntF),
    .i1(24'b000000000000000000000000),
    .o(\PWMF/n25 ));  // src/OnePWM.v(55)
  reg_sr_ss_w1 \PWMF/pwm_reg  (
    .clk(clk100m),
    .d(pwm[15]),
    .en(1'b1),
    .reset(~\PWMF/u14_sel_is_1_o ),
    .set(\PWMF/n18 ),
    .q(\PWMF/pwm_keep ));  // src/OnePWM.v(45)
  reg_sr_as_w1 \PWMF/reg0_b0  (
    .clk(clk100m),
    .d(\PWMF/n13 [0]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [0]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b1  (
    .clk(clk100m),
    .d(\PWMF/n13 [1]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [1]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b10  (
    .clk(clk100m),
    .d(\PWMF/n13 [10]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [10]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b11  (
    .clk(clk100m),
    .d(\PWMF/n13 [11]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [11]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b12  (
    .clk(clk100m),
    .d(\PWMF/n13 [12]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [12]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b13  (
    .clk(clk100m),
    .d(\PWMF/n13 [13]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [13]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b14  (
    .clk(clk100m),
    .d(\PWMF/n13 [14]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [14]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b15  (
    .clk(clk100m),
    .d(\PWMF/n13 [15]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [15]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b16  (
    .clk(clk100m),
    .d(\PWMF/n13 [16]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [16]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b17  (
    .clk(clk100m),
    .d(\PWMF/n13 [17]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [17]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b18  (
    .clk(clk100m),
    .d(\PWMF/n13 [18]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [18]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b19  (
    .clk(clk100m),
    .d(\PWMF/n13 [19]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [19]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b2  (
    .clk(clk100m),
    .d(\PWMF/n13 [2]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [2]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b20  (
    .clk(clk100m),
    .d(\PWMF/n13 [20]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [20]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b21  (
    .clk(clk100m),
    .d(\PWMF/n13 [21]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [21]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b22  (
    .clk(clk100m),
    .d(\PWMF/n13 [22]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [22]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b23  (
    .clk(clk100m),
    .d(\PWMF/n13 [23]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [23]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b24  (
    .clk(clk100m),
    .d(\PWMF/n13 [24]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [24]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b25  (
    .clk(clk100m),
    .d(\PWMF/n13 [25]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [25]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b26  (
    .clk(clk100m),
    .d(\PWMF/n13 [26]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [26]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b3  (
    .clk(clk100m),
    .d(\PWMF/n13 [3]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [3]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b4  (
    .clk(clk100m),
    .d(\PWMF/n13 [4]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [4]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b5  (
    .clk(clk100m),
    .d(\PWMF/n13 [5]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [5]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b6  (
    .clk(clk100m),
    .d(\PWMF/n13 [6]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [6]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b7  (
    .clk(clk100m),
    .d(\PWMF/n13 [7]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [7]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b8  (
    .clk(clk100m),
    .d(\PWMF/n13 [8]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [8]));  // src/OnePWM.v(37)
  reg_sr_as_w1 \PWMF/reg0_b9  (
    .clk(clk100m),
    .d(\PWMF/n13 [9]),
    .en(1'b1),
    .reset(~\PWMF/n11 ),
    .set(1'b0),
    .q(\PWMF/FreCnt [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b0  (
    .clk(clk100m),
    .d(freqF[0]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [0]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b1  (
    .clk(clk100m),
    .d(freqF[1]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [1]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b10  (
    .clk(clk100m),
    .d(freqF[10]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [10]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b11  (
    .clk(clk100m),
    .d(freqF[11]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [11]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b12  (
    .clk(clk100m),
    .d(freqF[12]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [12]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b13  (
    .clk(clk100m),
    .d(freqF[13]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [13]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b14  (
    .clk(clk100m),
    .d(freqF[14]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [14]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b15  (
    .clk(clk100m),
    .d(freqF[15]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [15]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b16  (
    .clk(clk100m),
    .d(freqF[16]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [16]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b17  (
    .clk(clk100m),
    .d(freqF[17]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [17]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b18  (
    .clk(clk100m),
    .d(freqF[18]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [18]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b19  (
    .clk(clk100m),
    .d(freqF[19]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [19]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b2  (
    .clk(clk100m),
    .d(freqF[2]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [2]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b20  (
    .clk(clk100m),
    .d(freqF[20]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [20]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b21  (
    .clk(clk100m),
    .d(freqF[21]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [21]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b22  (
    .clk(clk100m),
    .d(freqF[22]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [22]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b23  (
    .clk(clk100m),
    .d(freqF[23]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [23]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b24  (
    .clk(clk100m),
    .d(freqF[24]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [24]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b25  (
    .clk(clk100m),
    .d(freqF[25]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [25]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b26  (
    .clk(clk100m),
    .d(freqF[26]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [26]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b3  (
    .clk(clk100m),
    .d(freqF[3]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [3]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b4  (
    .clk(clk100m),
    .d(freqF[4]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [4]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b5  (
    .clk(clk100m),
    .d(freqF[5]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [5]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b6  (
    .clk(clk100m),
    .d(freqF[6]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [6]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b7  (
    .clk(clk100m),
    .d(freqF[7]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [7]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b8  (
    .clk(clk100m),
    .d(freqF[8]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [8]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg1_b9  (
    .clk(clk100m),
    .d(freqF[9]),
    .en(\PWMF/mux3_b0_sel_is_3_o ),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/FreCntr [9]));  // src/OnePWM.v(37)
  reg_ar_as_w1 \PWMF/reg2_b0  (
    .clk(clk100m),
    .d(\PWMF/n23 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[0]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b1  (
    .clk(clk100m),
    .d(\PWMF/n23 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[1]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b10  (
    .clk(clk100m),
    .d(\PWMF/n23 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[10]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b11  (
    .clk(clk100m),
    .d(\PWMF/n23 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[11]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b12  (
    .clk(clk100m),
    .d(\PWMF/n23 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[12]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b13  (
    .clk(clk100m),
    .d(\PWMF/n23 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[13]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b14  (
    .clk(clk100m),
    .d(\PWMF/n23 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[14]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b15  (
    .clk(clk100m),
    .d(\PWMF/n23 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[15]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b16  (
    .clk(clk100m),
    .d(\PWMF/n23 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[16]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b17  (
    .clk(clk100m),
    .d(\PWMF/n23 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[17]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b18  (
    .clk(clk100m),
    .d(\PWMF/n23 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[18]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b19  (
    .clk(clk100m),
    .d(\PWMF/n23 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[19]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b2  (
    .clk(clk100m),
    .d(\PWMF/n23 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[2]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b20  (
    .clk(clk100m),
    .d(\PWMF/n23 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[20]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b21  (
    .clk(clk100m),
    .d(\PWMF/n23 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[21]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b22  (
    .clk(clk100m),
    .d(\PWMF/n23 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[22]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b23  (
    .clk(clk100m),
    .d(\PWMF/n23 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[23]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b24  (
    .clk(clk100m),
    .d(\PWMF/n23 [24]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[24]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b25  (
    .clk(clk100m),
    .d(\PWMF/n23 [25]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[25]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b26  (
    .clk(clk100m),
    .d(\PWMF/n23 [26]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[26]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b27  (
    .clk(clk100m),
    .d(\PWMF/n23 [27]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[27]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b28  (
    .clk(clk100m),
    .d(\PWMF/n23 [28]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[28]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b29  (
    .clk(clk100m),
    .d(\PWMF/n23 [29]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[29]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b3  (
    .clk(clk100m),
    .d(\PWMF/n23 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[3]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b30  (
    .clk(clk100m),
    .d(\PWMF/n23 [30]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[30]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b31  (
    .clk(clk100m),
    .d(\PWMF/n23 [31]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[31]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b4  (
    .clk(clk100m),
    .d(\PWMF/n23 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[4]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b5  (
    .clk(clk100m),
    .d(\PWMF/n23 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[5]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b6  (
    .clk(clk100m),
    .d(\PWMF/n23 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[6]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b7  (
    .clk(clk100m),
    .d(\PWMF/n23 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[7]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b8  (
    .clk(clk100m),
    .d(\PWMF/n23 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[8]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg2_b9  (
    .clk(clk100m),
    .d(\PWMF/n23 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/pnumr[9]_keep ));  // src/OnePWM.v(48)
  reg_ar_as_w1 \PWMF/reg3_b0  (
    .clk(clk100m),
    .d(\PWMF/n31 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[0]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b1  (
    .clk(clk100m),
    .d(\PWMF/n31 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[1]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b10  (
    .clk(clk100m),
    .d(\PWMF/n31 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[10]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b11  (
    .clk(clk100m),
    .d(\PWMF/n31 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[11]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b12  (
    .clk(clk100m),
    .d(\PWMF/n31 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[12]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b13  (
    .clk(clk100m),
    .d(\PWMF/n31 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[13]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b14  (
    .clk(clk100m),
    .d(\PWMF/n31 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[14]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b15  (
    .clk(clk100m),
    .d(\PWMF/n31 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[15]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b16  (
    .clk(clk100m),
    .d(\PWMF/n31 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[16]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b17  (
    .clk(clk100m),
    .d(\PWMF/n31 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[17]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b18  (
    .clk(clk100m),
    .d(\PWMF/n31 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[18]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b19  (
    .clk(clk100m),
    .d(\PWMF/n31 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[19]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b2  (
    .clk(clk100m),
    .d(\PWMF/n31 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[2]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b20  (
    .clk(clk100m),
    .d(\PWMF/n31 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[20]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b21  (
    .clk(clk100m),
    .d(\PWMF/n31 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[21]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b22  (
    .clk(clk100m),
    .d(\PWMF/n31 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[22]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b23  (
    .clk(clk100m),
    .d(\PWMF/n31 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[23]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b3  (
    .clk(clk100m),
    .d(\PWMF/n31 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[3]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b4  (
    .clk(clk100m),
    .d(\PWMF/n31 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[4]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b5  (
    .clk(clk100m),
    .d(\PWMF/n31 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[5]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b6  (
    .clk(clk100m),
    .d(\PWMF/n31 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[6]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b7  (
    .clk(clk100m),
    .d(\PWMF/n31 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[7]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b8  (
    .clk(clk100m),
    .d(\PWMF/n31 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[8]_keep ));  // src/OnePWM.v(58)
  reg_ar_as_w1 \PWMF/reg3_b9  (
    .clk(clk100m),
    .d(\PWMF/n31 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\PWMF/RemaTxNum[9]_keep ));  // src/OnePWM.v(58)
  reg_ar_ss_w1 \PWMF/stopreq_reg  (
    .clk(clk100m),
    .d(\PWMF/n1 ),
    .en(1'b1),
    .reset(1'b0),
    .set(pwm_start_stop[15]),
    .q(\PWMF/stopreq_keep ));  // src/OnePWM.v(15)
  add_pu27_mu27_o27 \PWMF/sub0  (
    .i0(\PWMF/FreCnt ),
    .i1(27'b000000000000000000000000001),
    .o(\PWMF/n12 [26:0]));  // src/OnePWM.v(32)
  add_pu24_mu24_o24 \PWMF/sub1  (
    .i0(pnumcntF),
    .i1(24'b000000000000000000000001),
    .o(\PWMF/n26 [23:0]));  // src/OnePWM.v(55)
  AL_MUX \PWMF/u10  (
    .i0(1'b0),
    .i1(\PWMF/n9 ),
    .sel(n26),
    .o(\PWMF/n10 ));  // src/OnePWM.v(26)
  or \PWMF/u11  (\PWMF/n11 , pwm_state_read[15], pwm_start_stop[31]);  // src/OnePWM.v(30)
  and \PWMF/u14_sel_is_1  (\PWMF/u14_sel_is_1_o , pwm_state_read[15], \PWMF/n17_neg );
  and \PWMF/u15  (\PWMF/n24 , \PWMF/n0 , pwm_state_read[15]);  // src/OnePWM.v(54)
  and \PWMF/u17_sel_is_1  (\PWMF/u17_sel_is_1_o , \PWMF/n24 , \PWMF/n25_neg );
  not \PWMF/u17_sel_is_1_o_inv  (\PWMF/u17_sel_is_1_o_neg , \PWMF/u17_sel_is_1_o );
  AL_MUX \PWMF/u18  (
    .i0(\PWMF/pnumr [31]),
    .i1(dir[15]),
    .sel(\PWMF/u18_sel_is_0_o ),
    .o(\PWMF/n32 ));
  and \PWMF/u18_sel_is_0  (\PWMF/u18_sel_is_0_o , \pwm_start_stop[31]_neg , \PWMF/u17_sel_is_1_o_neg );
  AL_MUX \PWMF/u2  (
    .i0(\PWMF/stopreq ),
    .i1(1'b0),
    .sel(\PWMF/n0 ),
    .o(\PWMF/n1 ));  // src/OnePWM.v(15)
  and \PWMF/u5  (\PWMF/n4 , \PWMF/stopreq , \PWMF/n0 );  // src/OnePWM.v(23)
  and \PWMF/u6  (\PWMF/n6 , \PWMF/n5 , \PWMF/n0 );  // src/OnePWM.v(25)
  AL_MUX \PWMF/u8  (
    .i0(1'b0),
    .i1(pwm_state_read[15]),
    .sel(\PWMF/u8_sel_is_0_o ),
    .o(\PWMF/n8 ));
  and \PWMF/u8_sel_is_0  (\PWMF/u8_sel_is_0_o , \PWMF/n4_neg , \PWMF/n6_neg );
  AL_MUX \PWMF/u9  (
    .i0(\PWMF/n8 ),
    .i1(1'b1),
    .sel(pwm_start_stop[31]),
    .o(\PWMF/n9 ));  // src/OnePWM.v(26)
  EF2_PHY_MCU #(
    .GPIO_L0("ENABLE"),
    .GPIO_L1("ENABLE"),
    .GPIO_L10("DISABLE"),
    .GPIO_L11("DISABLE"),
    .GPIO_L12("DISABLE"),
    .GPIO_L13("DISABLE"),
    .GPIO_L14("DISABLE"),
    .GPIO_L15("DISABLE"),
    .GPIO_L2("DISABLE"),
    .GPIO_L3("DISABLE"),
    .GPIO_L4("DISABLE"),
    .GPIO_L5("DISABLE"),
    .GPIO_L6("DISABLE"),
    .GPIO_L7("DISABLE"),
    .GPIO_L8("ENABLE"),
    .GPIO_L9("ENABLE"))
    \U_AHB/M3WithAHB/mcu_inst  (
    .gpio_h_in(16'b0000000000000000),
    .h2h_hrdata(\U_AHB/h2h_hrdata ),
    .h2h_hreadyout(1'b1),
    .h2h_hresp(2'b00),
    .h2h_mclk(clk100m),
    .h2h_rstn(rstn),
    .ppm_clk(clk25m),
    .h2h_haddr({open_n43,open_n44,open_n45,open_n46,open_n47,open_n48,open_n49,open_n50,open_n51,open_n52,open_n53,open_n54,open_n55,open_n56,open_n57,open_n58,open_n59,\U_AHB/h2h_haddrw [14:2],open_n60,open_n61}),
    .h2h_hwdata(\U_AHB/h2h_hwdata ),
    .h2h_hwrite(\U_AHB/h2h_hwritew ));  // al_ip/M3WithAHB.v(46)
  eq_w2 \U_AHB/eq0  (
    .i0(\U_AHB/h2h_haddr [14:13]),
    .i1(2'b01),
    .o(\U_AHB/n0 ));  // src/AHB.v(46)
  eq_w2 \U_AHB/eq1  (
    .i0(\U_AHB/h2h_haddr [14:13]),
    .i1(2'b00),
    .o(\U_AHB/n6 ));  // src/AHB.v(48)
  eq_w2 \U_AHB/eq2  (
    .i0(\U_AHB/h2h_haddr [14:13]),
    .i1(2'b11),
    .o(\U_AHB/n43 ));  // src/AHB.v(67)
  eq_w2 \U_AHB/eq3  (
    .i0(\U_AHB/h2h_haddr [14:13]),
    .i1(2'b10),
    .o(\U_AHB/n49 ));  // src/AHB.v(69)
  reg_ar_as_w1 \U_AHB/h2h_hwrite_reg  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwritew ),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hwrite ));  // src/AHB.v(24)
  binary_mux_s1_w1 \U_AHB/mux16_b0  (
    .i0(gpio_out[0]),
    .i1(\U_AHB/n40 [0]),
    .sel(\U_AHB/n38 ),
    .o(\U_AHB/n41 [0]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux16_b1  (
    .i0(gpio_out[1]),
    .i1(\U_AHB/n40 [1]),
    .sel(\U_AHB/n38 ),
    .o(\U_AHB/n41 [1]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux16_b10  (
    .i0(gpio_out[10]),
    .i1(\U_AHB/n40 [10]),
    .sel(\U_AHB/n38 ),
    .o(\U_AHB/n41 [10]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux16_b11  (
    .i0(gpio_out[11]),
    .i1(\U_AHB/n40 [11]),
    .sel(\U_AHB/n38 ),
    .o(\U_AHB/n41 [11]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux16_b12  (
    .i0(gpio_out[12]),
    .i1(\U_AHB/n40 [12]),
    .sel(\U_AHB/n38 ),
    .o(\U_AHB/n41 [12]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux16_b13  (
    .i0(gpio_out[13]),
    .i1(\U_AHB/n40 [13]),
    .sel(\U_AHB/n38 ),
    .o(\U_AHB/n41 [13]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux16_b14  (
    .i0(gpio_out[14]),
    .i1(\U_AHB/n40 [14]),
    .sel(\U_AHB/n38 ),
    .o(\U_AHB/n41 [14]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux16_b15  (
    .i0(gpio_out[15]),
    .i1(\U_AHB/n40 [15]),
    .sel(\U_AHB/n38 ),
    .o(\U_AHB/n41 [15]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux16_b16  (
    .i0(gpio_out[16]),
    .i1(\U_AHB/n40 [16]),
    .sel(\U_AHB/n38 ),
    .o(\U_AHB/n41 [16]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux16_b17  (
    .i0(gpio_out[17]),
    .i1(\U_AHB/n40 [17]),
    .sel(\U_AHB/n38 ),
    .o(\U_AHB/n41 [17]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux16_b18  (
    .i0(gpio_out[18]),
    .i1(\U_AHB/n40 [18]),
    .sel(\U_AHB/n38 ),
    .o(\U_AHB/n41 [18]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux16_b19  (
    .i0(gpio_out[19]),
    .i1(\U_AHB/n40 [19]),
    .sel(\U_AHB/n38 ),
    .o(\U_AHB/n41 [19]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux16_b2  (
    .i0(gpio_out[2]),
    .i1(\U_AHB/n40 [2]),
    .sel(\U_AHB/n38 ),
    .o(\U_AHB/n41 [2]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux16_b20  (
    .i0(gpio_out[20]),
    .i1(\U_AHB/n40 [20]),
    .sel(\U_AHB/n38 ),
    .o(\U_AHB/n41 [20]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux16_b21  (
    .i0(gpio_out[21]),
    .i1(\U_AHB/n40 [21]),
    .sel(\U_AHB/n38 ),
    .o(\U_AHB/n41 [21]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux16_b22  (
    .i0(gpio_out[22]),
    .i1(\U_AHB/n40 [22]),
    .sel(\U_AHB/n38 ),
    .o(\U_AHB/n41 [22]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux16_b23  (
    .i0(gpio_out[23]),
    .i1(\U_AHB/n40 [23]),
    .sel(\U_AHB/n38 ),
    .o(\U_AHB/n41 [23]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux16_b24  (
    .i0(gpio_out[24]),
    .i1(\U_AHB/n40 [24]),
    .sel(\U_AHB/n38 ),
    .o(\U_AHB/n41 [24]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux16_b25  (
    .i0(gpio_out[25]),
    .i1(\U_AHB/n40 [25]),
    .sel(\U_AHB/n38 ),
    .o(\U_AHB/n41 [25]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux16_b26  (
    .i0(gpio_out[26]),
    .i1(\U_AHB/n40 [26]),
    .sel(\U_AHB/n38 ),
    .o(\U_AHB/n41 [26]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux16_b27  (
    .i0(gpio_out[27]),
    .i1(\U_AHB/n40 [27]),
    .sel(\U_AHB/n38 ),
    .o(\U_AHB/n41 [27]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux16_b28  (
    .i0(gpio_out[28]),
    .i1(\U_AHB/n40 [28]),
    .sel(\U_AHB/n38 ),
    .o(\U_AHB/n41 [28]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux16_b29  (
    .i0(gpio_out[29]),
    .i1(\U_AHB/n40 [29]),
    .sel(\U_AHB/n38 ),
    .o(\U_AHB/n41 [29]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux16_b3  (
    .i0(gpio_out[3]),
    .i1(\U_AHB/n40 [3]),
    .sel(\U_AHB/n38 ),
    .o(\U_AHB/n41 [3]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux16_b30  (
    .i0(gpio_out[30]),
    .i1(\U_AHB/n40 [30]),
    .sel(\U_AHB/n38 ),
    .o(\U_AHB/n41 [30]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux16_b31  (
    .i0(gpio_out[31]),
    .i1(\U_AHB/n40 [31]),
    .sel(\U_AHB/n38 ),
    .o(\U_AHB/n41 [31]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux16_b4  (
    .i0(gpio_out[4]),
    .i1(\U_AHB/n40 [4]),
    .sel(\U_AHB/n38 ),
    .o(\U_AHB/n41 [4]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux16_b5  (
    .i0(gpio_out[5]),
    .i1(\U_AHB/n40 [5]),
    .sel(\U_AHB/n38 ),
    .o(\U_AHB/n41 [5]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux16_b6  (
    .i0(gpio_out[6]),
    .i1(\U_AHB/n40 [6]),
    .sel(\U_AHB/n38 ),
    .o(\U_AHB/n41 [6]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux16_b7  (
    .i0(gpio_out[7]),
    .i1(\U_AHB/n40 [7]),
    .sel(\U_AHB/n38 ),
    .o(\U_AHB/n41 [7]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux16_b8  (
    .i0(gpio_out[8]),
    .i1(\U_AHB/n40 [8]),
    .sel(\U_AHB/n38 ),
    .o(\U_AHB/n41 [8]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux16_b9  (
    .i0(gpio_out[9]),
    .i1(\U_AHB/n40 [9]),
    .sel(\U_AHB/n38 ),
    .o(\U_AHB/n41 [9]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux17_b0  (
    .i0(\U_AHB/n41 [0]),
    .i1(\U_AHB/n37 [0]),
    .sel(\U_AHB/n36 ),
    .o(\U_AHB/n42 [0]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux17_b1  (
    .i0(\U_AHB/n41 [1]),
    .i1(\U_AHB/n37 [1]),
    .sel(\U_AHB/n36 ),
    .o(\U_AHB/n42 [1]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux17_b10  (
    .i0(\U_AHB/n41 [10]),
    .i1(\U_AHB/n37 [10]),
    .sel(\U_AHB/n36 ),
    .o(\U_AHB/n42 [10]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux17_b11  (
    .i0(\U_AHB/n41 [11]),
    .i1(\U_AHB/n37 [11]),
    .sel(\U_AHB/n36 ),
    .o(\U_AHB/n42 [11]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux17_b12  (
    .i0(\U_AHB/n41 [12]),
    .i1(\U_AHB/n37 [12]),
    .sel(\U_AHB/n36 ),
    .o(\U_AHB/n42 [12]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux17_b13  (
    .i0(\U_AHB/n41 [13]),
    .i1(\U_AHB/n37 [13]),
    .sel(\U_AHB/n36 ),
    .o(\U_AHB/n42 [13]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux17_b14  (
    .i0(\U_AHB/n41 [14]),
    .i1(\U_AHB/n37 [14]),
    .sel(\U_AHB/n36 ),
    .o(\U_AHB/n42 [14]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux17_b15  (
    .i0(\U_AHB/n41 [15]),
    .i1(\U_AHB/n37 [15]),
    .sel(\U_AHB/n36 ),
    .o(\U_AHB/n42 [15]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux17_b16  (
    .i0(\U_AHB/n41 [16]),
    .i1(\U_AHB/n37 [16]),
    .sel(\U_AHB/n36 ),
    .o(\U_AHB/n42 [16]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux17_b17  (
    .i0(\U_AHB/n41 [17]),
    .i1(\U_AHB/n37 [17]),
    .sel(\U_AHB/n36 ),
    .o(\U_AHB/n42 [17]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux17_b18  (
    .i0(\U_AHB/n41 [18]),
    .i1(\U_AHB/n37 [18]),
    .sel(\U_AHB/n36 ),
    .o(\U_AHB/n42 [18]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux17_b19  (
    .i0(\U_AHB/n41 [19]),
    .i1(\U_AHB/n37 [19]),
    .sel(\U_AHB/n36 ),
    .o(\U_AHB/n42 [19]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux17_b2  (
    .i0(\U_AHB/n41 [2]),
    .i1(\U_AHB/n37 [2]),
    .sel(\U_AHB/n36 ),
    .o(\U_AHB/n42 [2]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux17_b20  (
    .i0(\U_AHB/n41 [20]),
    .i1(\U_AHB/n37 [20]),
    .sel(\U_AHB/n36 ),
    .o(\U_AHB/n42 [20]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux17_b21  (
    .i0(\U_AHB/n41 [21]),
    .i1(\U_AHB/n37 [21]),
    .sel(\U_AHB/n36 ),
    .o(\U_AHB/n42 [21]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux17_b22  (
    .i0(\U_AHB/n41 [22]),
    .i1(\U_AHB/n37 [22]),
    .sel(\U_AHB/n36 ),
    .o(\U_AHB/n42 [22]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux17_b23  (
    .i0(\U_AHB/n41 [23]),
    .i1(\U_AHB/n37 [23]),
    .sel(\U_AHB/n36 ),
    .o(\U_AHB/n42 [23]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux17_b24  (
    .i0(\U_AHB/n41 [24]),
    .i1(\U_AHB/n37 [24]),
    .sel(\U_AHB/n36 ),
    .o(\U_AHB/n42 [24]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux17_b25  (
    .i0(\U_AHB/n41 [25]),
    .i1(\U_AHB/n37 [25]),
    .sel(\U_AHB/n36 ),
    .o(\U_AHB/n42 [25]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux17_b26  (
    .i0(\U_AHB/n41 [26]),
    .i1(\U_AHB/n37 [26]),
    .sel(\U_AHB/n36 ),
    .o(\U_AHB/n42 [26]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux17_b27  (
    .i0(\U_AHB/n41 [27]),
    .i1(\U_AHB/n37 [27]),
    .sel(\U_AHB/n36 ),
    .o(\U_AHB/n42 [27]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux17_b28  (
    .i0(\U_AHB/n41 [28]),
    .i1(\U_AHB/n37 [28]),
    .sel(\U_AHB/n36 ),
    .o(\U_AHB/n42 [28]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux17_b29  (
    .i0(\U_AHB/n41 [29]),
    .i1(\U_AHB/n37 [29]),
    .sel(\U_AHB/n36 ),
    .o(\U_AHB/n42 [29]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux17_b3  (
    .i0(\U_AHB/n41 [3]),
    .i1(\U_AHB/n37 [3]),
    .sel(\U_AHB/n36 ),
    .o(\U_AHB/n42 [3]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux17_b30  (
    .i0(\U_AHB/n41 [30]),
    .i1(\U_AHB/n37 [30]),
    .sel(\U_AHB/n36 ),
    .o(\U_AHB/n42 [30]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux17_b31  (
    .i0(\U_AHB/n41 [31]),
    .i1(\U_AHB/n37 [31]),
    .sel(\U_AHB/n36 ),
    .o(\U_AHB/n42 [31]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux17_b4  (
    .i0(\U_AHB/n41 [4]),
    .i1(\U_AHB/n37 [4]),
    .sel(\U_AHB/n36 ),
    .o(\U_AHB/n42 [4]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux17_b5  (
    .i0(\U_AHB/n41 [5]),
    .i1(\U_AHB/n37 [5]),
    .sel(\U_AHB/n36 ),
    .o(\U_AHB/n42 [5]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux17_b6  (
    .i0(\U_AHB/n41 [6]),
    .i1(\U_AHB/n37 [6]),
    .sel(\U_AHB/n36 ),
    .o(\U_AHB/n42 [6]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux17_b7  (
    .i0(\U_AHB/n41 [7]),
    .i1(\U_AHB/n37 [7]),
    .sel(\U_AHB/n36 ),
    .o(\U_AHB/n42 [7]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux17_b8  (
    .i0(\U_AHB/n41 [8]),
    .i1(\U_AHB/n37 [8]),
    .sel(\U_AHB/n36 ),
    .o(\U_AHB/n42 [8]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux17_b9  (
    .i0(\U_AHB/n41 [9]),
    .i1(\U_AHB/n37 [9]),
    .sel(\U_AHB/n36 ),
    .o(\U_AHB/n42 [9]));  // src/AHB.v(64)
  binary_mux_s1_w1 \U_AHB/mux35_b0  (
    .i0(\U_AHB/h2h_hrdata [0]),
    .i1(\U_AHB/n116 [0]),
    .sel(\U_AHB/n115 ),
    .o(\U_AHB/n117 [0]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux35_b1  (
    .i0(\U_AHB/h2h_hrdata [1]),
    .i1(\U_AHB/n116 [1]),
    .sel(\U_AHB/n115 ),
    .o(\U_AHB/n117 [1]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux35_b10  (
    .i0(\U_AHB/h2h_hrdata [10]),
    .i1(\U_AHB/n116 [10]),
    .sel(\U_AHB/n115 ),
    .o(\U_AHB/n117 [10]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux35_b11  (
    .i0(\U_AHB/h2h_hrdata [11]),
    .i1(\U_AHB/n116 [11]),
    .sel(\U_AHB/n115 ),
    .o(\U_AHB/n117 [11]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux35_b12  (
    .i0(\U_AHB/h2h_hrdata [12]),
    .i1(\U_AHB/n116 [12]),
    .sel(\U_AHB/n115 ),
    .o(\U_AHB/n117 [12]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux35_b13  (
    .i0(\U_AHB/h2h_hrdata [13]),
    .i1(\U_AHB/n116 [13]),
    .sel(\U_AHB/n115 ),
    .o(\U_AHB/n117 [13]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux35_b14  (
    .i0(\U_AHB/h2h_hrdata [14]),
    .i1(\U_AHB/n116 [14]),
    .sel(\U_AHB/n115 ),
    .o(\U_AHB/n117 [14]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux35_b15  (
    .i0(\U_AHB/h2h_hrdata [15]),
    .i1(\U_AHB/n116 [15]),
    .sel(\U_AHB/n115 ),
    .o(\U_AHB/n117 [15]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux35_b16  (
    .i0(\U_AHB/h2h_hrdata [16]),
    .i1(\U_AHB/n116 [16]),
    .sel(\U_AHB/n115 ),
    .o(\U_AHB/n117 [16]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux35_b17  (
    .i0(\U_AHB/h2h_hrdata [17]),
    .i1(\U_AHB/n116 [17]),
    .sel(\U_AHB/n115 ),
    .o(\U_AHB/n117 [17]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux35_b18  (
    .i0(\U_AHB/h2h_hrdata [18]),
    .i1(\U_AHB/n116 [18]),
    .sel(\U_AHB/n115 ),
    .o(\U_AHB/n117 [18]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux35_b19  (
    .i0(\U_AHB/h2h_hrdata [19]),
    .i1(\U_AHB/n116 [19]),
    .sel(\U_AHB/n115 ),
    .o(\U_AHB/n117 [19]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux35_b2  (
    .i0(\U_AHB/h2h_hrdata [2]),
    .i1(\U_AHB/n116 [2]),
    .sel(\U_AHB/n115 ),
    .o(\U_AHB/n117 [2]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux35_b20  (
    .i0(\U_AHB/h2h_hrdata [20]),
    .i1(\U_AHB/n116 [20]),
    .sel(\U_AHB/n115 ),
    .o(\U_AHB/n117 [20]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux35_b21  (
    .i0(\U_AHB/h2h_hrdata [21]),
    .i1(\U_AHB/n116 [21]),
    .sel(\U_AHB/n115 ),
    .o(\U_AHB/n117 [21]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux35_b22  (
    .i0(\U_AHB/h2h_hrdata [22]),
    .i1(\U_AHB/n116 [22]),
    .sel(\U_AHB/n115 ),
    .o(\U_AHB/n117 [22]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux35_b23  (
    .i0(\U_AHB/h2h_hrdata [23]),
    .i1(\U_AHB/n116 [23]),
    .sel(\U_AHB/n115 ),
    .o(\U_AHB/n117 [23]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux35_b24  (
    .i0(\U_AHB/h2h_hrdata [24]),
    .i1(\U_AHB/sel1_b24/or_or_B0_B1_o_or_B2__o ),
    .sel(\U_AHB/n115 ),
    .o(\U_AHB/n117 [24]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux35_b25  (
    .i0(\U_AHB/h2h_hrdata [25]),
    .i1(\U_AHB/sel1_b25/or_or_B0_B1_o_or_B2__o ),
    .sel(\U_AHB/n115 ),
    .o(\U_AHB/n117 [25]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux35_b26  (
    .i0(\U_AHB/h2h_hrdata [26]),
    .i1(\U_AHB/sel1_b26/or_or_B0_B1_o_or_B2__o ),
    .sel(\U_AHB/n115 ),
    .o(\U_AHB/n117 [26]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux35_b27  (
    .i0(\U_AHB/h2h_hrdata [27]),
    .i1(\U_AHB/sel1_b27/or_or_B0_B1_o_or_B2__o ),
    .sel(\U_AHB/n115 ),
    .o(\U_AHB/n117 [27]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux35_b28  (
    .i0(\U_AHB/h2h_hrdata [28]),
    .i1(\U_AHB/sel1_b28/or_or_B0_B1_o_or_B2__o ),
    .sel(\U_AHB/n115 ),
    .o(\U_AHB/n117 [28]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux35_b29  (
    .i0(\U_AHB/h2h_hrdata [29]),
    .i1(\U_AHB/sel1_b29/or_or_B0_B1_o_or_B2__o ),
    .sel(\U_AHB/n115 ),
    .o(\U_AHB/n117 [29]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux35_b3  (
    .i0(\U_AHB/h2h_hrdata [3]),
    .i1(\U_AHB/n116 [3]),
    .sel(\U_AHB/n115 ),
    .o(\U_AHB/n117 [3]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux35_b30  (
    .i0(\U_AHB/h2h_hrdata [30]),
    .i1(\U_AHB/sel1_b30/or_or_B0_B1_o_or_B2__o ),
    .sel(\U_AHB/n115 ),
    .o(\U_AHB/n117 [30]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux35_b31  (
    .i0(\U_AHB/h2h_hrdata [31]),
    .i1(\U_AHB/sel1_b31/or_or_B0_B1_o_or_B2__o ),
    .sel(\U_AHB/n115 ),
    .o(\U_AHB/n117 [31]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux35_b4  (
    .i0(\U_AHB/h2h_hrdata [4]),
    .i1(\U_AHB/n116 [4]),
    .sel(\U_AHB/n115 ),
    .o(\U_AHB/n117 [4]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux35_b5  (
    .i0(\U_AHB/h2h_hrdata [5]),
    .i1(\U_AHB/n116 [5]),
    .sel(\U_AHB/n115 ),
    .o(\U_AHB/n117 [5]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux35_b6  (
    .i0(\U_AHB/h2h_hrdata [6]),
    .i1(\U_AHB/n116 [6]),
    .sel(\U_AHB/n115 ),
    .o(\U_AHB/n117 [6]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux35_b7  (
    .i0(\U_AHB/h2h_hrdata [7]),
    .i1(\U_AHB/n116 [7]),
    .sel(\U_AHB/n115 ),
    .o(\U_AHB/n117 [7]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux35_b8  (
    .i0(\U_AHB/h2h_hrdata [8]),
    .i1(\U_AHB/n116 [8]),
    .sel(\U_AHB/n115 ),
    .o(\U_AHB/n117 [8]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux35_b9  (
    .i0(\U_AHB/h2h_hrdata [9]),
    .i1(\U_AHB/n116 [9]),
    .sel(\U_AHB/n115 ),
    .o(\U_AHB/n117 [9]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux36_b0  (
    .i0(\U_AHB/n117 [0]),
    .i1(\U_AHB/n114 [0]),
    .sel(\U_AHB/n82 ),
    .o(\U_AHB/n118 [0]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux36_b1  (
    .i0(\U_AHB/n117 [1]),
    .i1(\U_AHB/n114 [1]),
    .sel(\U_AHB/n82 ),
    .o(\U_AHB/n118 [1]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux36_b10  (
    .i0(\U_AHB/n117 [10]),
    .i1(\U_AHB/n114 [10]),
    .sel(\U_AHB/n82 ),
    .o(\U_AHB/n118 [10]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux36_b11  (
    .i0(\U_AHB/n117 [11]),
    .i1(\U_AHB/n114 [11]),
    .sel(\U_AHB/n82 ),
    .o(\U_AHB/n118 [11]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux36_b12  (
    .i0(\U_AHB/n117 [12]),
    .i1(\U_AHB/n114 [12]),
    .sel(\U_AHB/n82 ),
    .o(\U_AHB/n118 [12]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux36_b13  (
    .i0(\U_AHB/n117 [13]),
    .i1(\U_AHB/n114 [13]),
    .sel(\U_AHB/n82 ),
    .o(\U_AHB/n118 [13]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux36_b14  (
    .i0(\U_AHB/n117 [14]),
    .i1(\U_AHB/n114 [14]),
    .sel(\U_AHB/n82 ),
    .o(\U_AHB/n118 [14]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux36_b15  (
    .i0(\U_AHB/n117 [15]),
    .i1(\U_AHB/n114 [15]),
    .sel(\U_AHB/n82 ),
    .o(\U_AHB/n118 [15]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux36_b16  (
    .i0(\U_AHB/n117 [16]),
    .i1(\U_AHB/n114 [16]),
    .sel(\U_AHB/n82 ),
    .o(\U_AHB/n118 [16]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux36_b17  (
    .i0(\U_AHB/n117 [17]),
    .i1(\U_AHB/n114 [17]),
    .sel(\U_AHB/n82 ),
    .o(\U_AHB/n118 [17]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux36_b18  (
    .i0(\U_AHB/n117 [18]),
    .i1(\U_AHB/n114 [18]),
    .sel(\U_AHB/n82 ),
    .o(\U_AHB/n118 [18]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux36_b19  (
    .i0(\U_AHB/n117 [19]),
    .i1(\U_AHB/n114 [19]),
    .sel(\U_AHB/n82 ),
    .o(\U_AHB/n118 [19]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux36_b2  (
    .i0(\U_AHB/n117 [2]),
    .i1(\U_AHB/n114 [2]),
    .sel(\U_AHB/n82 ),
    .o(\U_AHB/n118 [2]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux36_b20  (
    .i0(\U_AHB/n117 [20]),
    .i1(\U_AHB/n114 [20]),
    .sel(\U_AHB/n82 ),
    .o(\U_AHB/n118 [20]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux36_b21  (
    .i0(\U_AHB/n117 [21]),
    .i1(\U_AHB/n114 [21]),
    .sel(\U_AHB/n82 ),
    .o(\U_AHB/n118 [21]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux36_b22  (
    .i0(\U_AHB/n117 [22]),
    .i1(\U_AHB/n114 [22]),
    .sel(\U_AHB/n82 ),
    .o(\U_AHB/n118 [22]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux36_b23  (
    .i0(\U_AHB/n117 [23]),
    .i1(\U_AHB/n114 [23]),
    .sel(\U_AHB/n82 ),
    .o(\U_AHB/n118 [23]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux36_b24  (
    .i0(\U_AHB/n117 [24]),
    .i1(\U_AHB/n114 [24]),
    .sel(\U_AHB/n82 ),
    .o(\U_AHB/n118 [24]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux36_b25  (
    .i0(\U_AHB/n117 [25]),
    .i1(\U_AHB/n114 [25]),
    .sel(\U_AHB/n82 ),
    .o(\U_AHB/n118 [25]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux36_b26  (
    .i0(\U_AHB/n117 [26]),
    .i1(\U_AHB/n114 [26]),
    .sel(\U_AHB/n82 ),
    .o(\U_AHB/n118 [26]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux36_b27  (
    .i0(\U_AHB/n117 [27]),
    .i1(\U_AHB/n114 [27]),
    .sel(\U_AHB/n82 ),
    .o(\U_AHB/n118 [27]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux36_b28  (
    .i0(\U_AHB/n117 [28]),
    .i1(\U_AHB/n114 [28]),
    .sel(\U_AHB/n82 ),
    .o(\U_AHB/n118 [28]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux36_b29  (
    .i0(\U_AHB/n117 [29]),
    .i1(\U_AHB/n114 [29]),
    .sel(\U_AHB/n82 ),
    .o(\U_AHB/n118 [29]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux36_b3  (
    .i0(\U_AHB/n117 [3]),
    .i1(\U_AHB/n114 [3]),
    .sel(\U_AHB/n82 ),
    .o(\U_AHB/n118 [3]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux36_b30  (
    .i0(\U_AHB/n117 [30]),
    .i1(\U_AHB/n114 [30]),
    .sel(\U_AHB/n82 ),
    .o(\U_AHB/n118 [30]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux36_b31  (
    .i0(\U_AHB/n117 [31]),
    .i1(\U_AHB/n114 [31]),
    .sel(\U_AHB/n82 ),
    .o(\U_AHB/n118 [31]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux36_b4  (
    .i0(\U_AHB/n117 [4]),
    .i1(\U_AHB/n114 [4]),
    .sel(\U_AHB/n82 ),
    .o(\U_AHB/n118 [4]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux36_b5  (
    .i0(\U_AHB/n117 [5]),
    .i1(\U_AHB/n114 [5]),
    .sel(\U_AHB/n82 ),
    .o(\U_AHB/n118 [5]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux36_b6  (
    .i0(\U_AHB/n117 [6]),
    .i1(\U_AHB/n114 [6]),
    .sel(\U_AHB/n82 ),
    .o(\U_AHB/n118 [6]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux36_b7  (
    .i0(\U_AHB/n117 [7]),
    .i1(\U_AHB/n114 [7]),
    .sel(\U_AHB/n82 ),
    .o(\U_AHB/n118 [7]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux36_b8  (
    .i0(\U_AHB/n117 [8]),
    .i1(\U_AHB/n114 [8]),
    .sel(\U_AHB/n82 ),
    .o(\U_AHB/n118 [8]));  // src/AHB.v(114)
  binary_mux_s1_w1 \U_AHB/mux36_b9  (
    .i0(\U_AHB/n117 [9]),
    .i1(\U_AHB/n114 [9]),
    .sel(\U_AHB/n82 ),
    .o(\U_AHB/n118 [9]));  // src/AHB.v(114)
  reg_ar_as_w1 \U_AHB/reg0_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_haddrw [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_haddr [2]));  // src/AHB.v(25)
  reg_ar_as_w1 \U_AHB/reg0_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_haddrw [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_haddr [3]));  // src/AHB.v(25)
  reg_ar_as_w1 \U_AHB/reg0_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_haddrw [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_haddr [12]));  // src/AHB.v(25)
  reg_ar_as_w1 \U_AHB/reg0_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_haddrw [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_haddr [13]));  // src/AHB.v(25)
  reg_ar_as_w1 \U_AHB/reg0_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_haddrw [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_haddr [14]));  // src/AHB.v(25)
  reg_ar_as_w1 \U_AHB/reg0_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_haddrw [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_haddr [4]));  // src/AHB.v(25)
  reg_ar_as_w1 \U_AHB/reg0_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_haddrw [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_haddr [5]));  // src/AHB.v(25)
  reg_ar_as_w1 \U_AHB/reg0_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_haddrw [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_haddr [6]));  // src/AHB.v(25)
  reg_ar_as_w1 \U_AHB/reg0_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_haddrw [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_haddr [7]));  // src/AHB.v(25)
  reg_ar_as_w1 \U_AHB/reg0_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_haddrw [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_haddr [8]));  // src/AHB.v(25)
  reg_ar_as_w1 \U_AHB/reg0_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_haddrw [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_haddr [9]));  // src/AHB.v(25)
  reg_ar_as_w1 \U_AHB/reg0_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_haddrw [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_haddr [10]));  // src/AHB.v(25)
  reg_ar_as_w1 \U_AHB/reg0_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_haddrw [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_haddr [11]));  // src/AHB.v(25)
  reg_ar_as_w1 \U_AHB/reg10_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[0]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[1]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[10]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[11]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[12]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[13]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[14]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[15]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[16]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[17]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[18]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[19]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[2]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[20]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[21]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[22]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[23]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[24]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[25]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[26]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[3]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[4]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[5]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[6]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[7]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[8]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg10_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(\U_AHB/n22 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq9[9]));  // src/AHB.v(55)
  reg_ar_as_w1 \U_AHB/reg11_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[0]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[1]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[10]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[11]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[12]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[13]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[14]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[15]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[16]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[17]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[18]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[19]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[2]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[20]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[21]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[22]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[23]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[24]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[25]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[26]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[3]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[4]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[5]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[6]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[7]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[8]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg11_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(\U_AHB/n24 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqA[9]));  // src/AHB.v(56)
  reg_ar_as_w1 \U_AHB/reg12_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[0]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[1]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[10]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[11]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[12]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[13]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[14]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[15]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[16]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[17]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[18]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[19]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[2]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[20]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[21]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[22]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[23]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[24]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[25]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[26]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[3]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[4]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[5]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[6]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[7]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[8]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg12_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(\U_AHB/n26 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqB[9]));  // src/AHB.v(57)
  reg_ar_as_w1 \U_AHB/reg13_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[0]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[1]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[10]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[11]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[12]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[13]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[14]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[15]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[16]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[17]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[18]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[19]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[2]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[20]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[21]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[22]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[23]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[24]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[25]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[26]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[3]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[4]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[5]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[6]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[7]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[8]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg13_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(\U_AHB/n28 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqC[9]));  // src/AHB.v(58)
  reg_ar_as_w1 \U_AHB/reg14_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[0]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[1]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[10]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[11]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[12]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[13]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[14]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[15]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[16]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[17]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[18]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[19]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[2]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[20]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[21]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[22]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[23]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[24]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[25]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[26]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[3]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[4]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[5]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[6]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[7]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[8]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg14_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(\U_AHB/n30 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqD[9]));  // src/AHB.v(60)
  reg_ar_as_w1 \U_AHB/reg15_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[0]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[1]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[10]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[11]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[12]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[13]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[14]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[15]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[16]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[17]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[18]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[19]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[2]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[20]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[21]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[22]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[23]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[24]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[25]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[26]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[3]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[4]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[5]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[6]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[7]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[8]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg15_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(\U_AHB/n32 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqE[9]));  // src/AHB.v(61)
  reg_ar_as_w1 \U_AHB/reg16_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[0]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[1]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[10]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[11]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[12]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[13]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[14]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[15]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[16]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[17]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[18]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[19]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[2]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[20]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[21]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[22]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[23]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[24]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[25]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[26]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[3]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[4]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[5]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[6]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[7]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[8]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg16_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(\U_AHB/n34 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freqF[9]));  // src/AHB.v(62)
  reg_ar_as_w1 \U_AHB/reg17_b0  (
    .clk(clk100m),
    .d(\U_AHB/n42 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out[0]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b1  (
    .clk(clk100m),
    .d(\U_AHB/n42 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out[1]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b10  (
    .clk(clk100m),
    .d(\U_AHB/n42 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out[10]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b11  (
    .clk(clk100m),
    .d(\U_AHB/n42 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out[11]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b12  (
    .clk(clk100m),
    .d(\U_AHB/n42 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out[12]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b13  (
    .clk(clk100m),
    .d(\U_AHB/n42 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out[13]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b14  (
    .clk(clk100m),
    .d(\U_AHB/n42 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out[14]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b15  (
    .clk(clk100m),
    .d(\U_AHB/n42 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out[15]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b16  (
    .clk(clk100m),
    .d(\U_AHB/n42 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out[16]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b17  (
    .clk(clk100m),
    .d(\U_AHB/n42 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out[17]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b18  (
    .clk(clk100m),
    .d(\U_AHB/n42 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out[18]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b19  (
    .clk(clk100m),
    .d(\U_AHB/n42 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out[19]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b2  (
    .clk(clk100m),
    .d(\U_AHB/n42 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out[2]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b20  (
    .clk(clk100m),
    .d(\U_AHB/n42 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out[20]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b21  (
    .clk(clk100m),
    .d(\U_AHB/n42 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out[21]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b22  (
    .clk(clk100m),
    .d(\U_AHB/n42 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out[22]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b23  (
    .clk(clk100m),
    .d(\U_AHB/n42 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out[23]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b24  (
    .clk(clk100m),
    .d(\U_AHB/n42 [24]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out[24]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b25  (
    .clk(clk100m),
    .d(\U_AHB/n42 [25]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out[25]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b26  (
    .clk(clk100m),
    .d(\U_AHB/n42 [26]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out[26]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b27  (
    .clk(clk100m),
    .d(\U_AHB/n42 [27]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out[27]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b28  (
    .clk(clk100m),
    .d(\U_AHB/n42 [28]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out[28]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b29  (
    .clk(clk100m),
    .d(\U_AHB/n42 [29]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out[29]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b3  (
    .clk(clk100m),
    .d(\U_AHB/n42 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out[3]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b30  (
    .clk(clk100m),
    .d(\U_AHB/n42 [30]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out[30]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b31  (
    .clk(clk100m),
    .d(\U_AHB/n42 [31]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out[31]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b4  (
    .clk(clk100m),
    .d(\U_AHB/n42 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out[4]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b5  (
    .clk(clk100m),
    .d(\U_AHB/n42 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out[5]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b6  (
    .clk(clk100m),
    .d(\U_AHB/n42 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out[6]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b7  (
    .clk(clk100m),
    .d(\U_AHB/n42 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out[7]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b8  (
    .clk(clk100m),
    .d(\U_AHB/n42 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out[8]));  // src/AHB.v(64)
  reg_ar_as_w1 \U_AHB/reg17_b9  (
    .clk(clk100m),
    .d(\U_AHB/n42 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(gpio_out[9]));  // src/AHB.v(64)
  reg_sr_as_w1 \U_AHB/reg18_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[0]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[1]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[10]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[11]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[12]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[13]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[14]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[15]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[16]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[17]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[18]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[19]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[2]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[20]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[21]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[22]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[23]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[24]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[25]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[26]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b27  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [27]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[27]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b28  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [28]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[28]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b29  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [29]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[29]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[3]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b30  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [30]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[30]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b31  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [31]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[31]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b32  (
    .clk(clk100m),
    .d(1'b1),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[32]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[4]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[5]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[6]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[7]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[8]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg18_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(1'b1),
    .reset(~\U_AHB/n45 ),
    .set(1'b0),
    .q(pnum0[9]));  // src/AHB.v(67)
  reg_sr_as_w1 \U_AHB/reg19_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[0]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[1]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[10]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[11]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[12]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[13]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[14]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[15]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[16]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[17]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[18]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[19]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[2]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[20]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[21]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[22]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[23]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[24]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[25]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[26]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b27  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [27]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[27]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b28  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [28]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[28]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b29  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [29]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[29]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[3]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b30  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [30]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[30]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b31  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [31]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[31]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b32  (
    .clk(clk100m),
    .d(1'b1),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[32]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[4]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[5]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[6]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[7]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[8]));  // src/AHB.v(68)
  reg_sr_as_w1 \U_AHB/reg19_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(1'b1),
    .reset(~\U_AHB/n47 ),
    .set(1'b0),
    .q(pnum1[9]));  // src/AHB.v(68)
  reg_ar_as_w1 \U_AHB/reg1_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[0]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[1]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[10]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[11]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[12]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[13]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[14]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[15]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[16]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[17]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[18]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[19]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[2]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[20]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[21]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[22]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[23]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[24]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[25]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[26]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[3]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[4]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[5]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[6]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[7]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[8]));  // src/AHB.v(46)
  reg_ar_as_w1 \U_AHB/reg1_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(\U_AHB/n2 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq0[9]));  // src/AHB.v(46)
  reg_sr_as_w1 \U_AHB/reg20_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[0]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[1]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[10]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[11]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[12]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[13]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[14]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[15]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[16]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[17]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[18]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[19]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[2]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[20]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[21]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[22]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[23]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[24]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[25]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[26]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b27  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [27]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[27]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b28  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [28]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[28]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b29  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [29]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[29]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[3]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b30  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [30]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[30]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b31  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [31]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[31]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b32  (
    .clk(clk100m),
    .d(1'b1),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[32]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[4]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[5]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[6]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[7]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[8]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg20_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(1'b1),
    .reset(~\U_AHB/n51 ),
    .set(1'b0),
    .q(pnum2[9]));  // src/AHB.v(69)
  reg_sr_as_w1 \U_AHB/reg21_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[0]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[1]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[10]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[11]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[12]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[13]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[14]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[15]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[16]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[17]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[18]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[19]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[2]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[20]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[21]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[22]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[23]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[24]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[25]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[26]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b27  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [27]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[27]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b28  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [28]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[28]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b29  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [29]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[29]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[3]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b30  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [30]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[30]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b31  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [31]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[31]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b32  (
    .clk(clk100m),
    .d(1'b1),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[32]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[4]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[5]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[6]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[7]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[8]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg21_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(1'b1),
    .reset(~\U_AHB/n53 ),
    .set(1'b0),
    .q(pnum3[9]));  // src/AHB.v(70)
  reg_sr_as_w1 \U_AHB/reg22_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[0]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[1]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[10]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[11]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[12]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[13]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[14]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[15]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[16]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[17]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[18]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[19]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[2]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[20]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[21]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[22]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[23]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[24]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[25]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[26]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b27  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [27]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[27]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b28  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [28]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[28]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b29  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [29]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[29]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[3]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b30  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [30]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[30]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b31  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [31]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[31]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b32  (
    .clk(clk100m),
    .d(1'b1),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[32]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[4]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[5]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[6]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[7]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[8]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg22_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(1'b1),
    .reset(~\U_AHB/n55 ),
    .set(1'b0),
    .q(pnum4[9]));  // src/AHB.v(71)
  reg_sr_as_w1 \U_AHB/reg23_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[0]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[1]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[10]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[11]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[12]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[13]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[14]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[15]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[16]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[17]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[18]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[19]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[2]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[20]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[21]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[22]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[23]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[24]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[25]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[26]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b27  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [27]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[27]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b28  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [28]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[28]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b29  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [29]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[29]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[3]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b30  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [30]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[30]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b31  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [31]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[31]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b32  (
    .clk(clk100m),
    .d(1'b1),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[32]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[4]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[5]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[6]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[7]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[8]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg23_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(1'b1),
    .reset(~\U_AHB/n57 ),
    .set(1'b0),
    .q(pnum5[9]));  // src/AHB.v(72)
  reg_sr_as_w1 \U_AHB/reg24_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[0]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[1]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[10]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[11]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[12]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[13]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[14]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[15]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[16]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[17]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[18]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[19]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[2]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[20]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[21]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[22]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[23]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[24]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[25]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[26]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b27  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [27]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[27]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b28  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [28]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[28]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b29  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [29]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[29]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[3]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b30  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [30]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[30]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b31  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [31]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[31]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b32  (
    .clk(clk100m),
    .d(1'b1),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[32]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[4]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[5]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[6]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[7]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[8]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg24_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(1'b1),
    .reset(~\U_AHB/n59 ),
    .set(1'b0),
    .q(pnum6[9]));  // src/AHB.v(73)
  reg_sr_as_w1 \U_AHB/reg25_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[0]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[1]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[10]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[11]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[12]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[13]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[14]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[15]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[16]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[17]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[18]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[19]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[2]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[20]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[21]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[22]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[23]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[24]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[25]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[26]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b27  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [27]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[27]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b28  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [28]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[28]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b29  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [29]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[29]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[3]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b30  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [30]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[30]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b31  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [31]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[31]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b32  (
    .clk(clk100m),
    .d(1'b1),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[32]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[4]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[5]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[6]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[7]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[8]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg25_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(1'b1),
    .reset(~\U_AHB/n61 ),
    .set(1'b0),
    .q(pnum7[9]));  // src/AHB.v(74)
  reg_sr_as_w1 \U_AHB/reg26_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[0]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[1]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[10]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[11]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[12]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[13]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[14]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[15]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[16]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[17]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[18]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[19]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[2]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[20]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[21]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[22]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[23]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[24]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[25]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[26]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b27  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [27]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[27]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b28  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [28]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[28]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b29  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [29]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[29]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[3]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b30  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [30]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[30]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b31  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [31]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[31]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b32  (
    .clk(clk100m),
    .d(1'b1),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[32]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[4]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[5]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[6]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[7]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[8]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg26_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(1'b1),
    .reset(~\U_AHB/n63 ),
    .set(1'b0),
    .q(pnum8[9]));  // src/AHB.v(75)
  reg_sr_as_w1 \U_AHB/reg27_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[0]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[1]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[10]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[11]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[12]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[13]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[14]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[15]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[16]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[17]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[18]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[19]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[2]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[20]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[21]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[22]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[23]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[24]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[25]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[26]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b27  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [27]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[27]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b28  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [28]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[28]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b29  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [29]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[29]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[3]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b30  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [30]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[30]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b31  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [31]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[31]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b32  (
    .clk(clk100m),
    .d(1'b1),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[32]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[4]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[5]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[6]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[7]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[8]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg27_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(1'b1),
    .reset(~\U_AHB/n65 ),
    .set(1'b0),
    .q(pnum9[9]));  // src/AHB.v(76)
  reg_sr_as_w1 \U_AHB/reg28_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[0]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[1]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[10]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[11]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[12]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[13]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[14]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[15]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[16]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[17]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[18]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[19]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[2]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[20]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[21]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[22]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[23]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[24]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[25]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[26]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b27  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [27]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[27]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b28  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [28]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[28]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b29  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [29]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[29]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[3]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b30  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [30]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[30]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b31  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [31]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[31]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b32  (
    .clk(clk100m),
    .d(1'b1),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[32]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[4]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[5]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[6]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[7]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[8]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg28_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(1'b1),
    .reset(~\U_AHB/n67 ),
    .set(1'b0),
    .q(pnumA[9]));  // src/AHB.v(77)
  reg_sr_as_w1 \U_AHB/reg29_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[0]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[1]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[10]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[11]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[12]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[13]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[14]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[15]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[16]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[17]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[18]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[19]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[2]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[20]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[21]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[22]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[23]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[24]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[25]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[26]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b27  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [27]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[27]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b28  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [28]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[28]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b29  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [29]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[29]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[3]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b30  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [30]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[30]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b31  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [31]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[31]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b32  (
    .clk(clk100m),
    .d(1'b1),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[32]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[4]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[5]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[6]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[7]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[8]));  // src/AHB.v(78)
  reg_sr_as_w1 \U_AHB/reg29_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(1'b1),
    .reset(~\U_AHB/n69 ),
    .set(1'b0),
    .q(pnumB[9]));  // src/AHB.v(78)
  reg_ar_as_w1 \U_AHB/reg2_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[0]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[1]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[10]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[11]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[12]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[13]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[14]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[15]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[16]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[17]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[18]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[19]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[2]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[20]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[21]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[22]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[23]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[24]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[25]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[26]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[3]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[4]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[5]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[6]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[7]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[8]));  // src/AHB.v(47)
  reg_ar_as_w1 \U_AHB/reg2_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(\U_AHB/n4 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq1[9]));  // src/AHB.v(47)
  reg_sr_as_w1 \U_AHB/reg30_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[0]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[1]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[10]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[11]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[12]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[13]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[14]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[15]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[16]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[17]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[18]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[19]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[2]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[20]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[21]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[22]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[23]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[24]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[25]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[26]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b27  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [27]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[27]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b28  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [28]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[28]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b29  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [29]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[29]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[3]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b30  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [30]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[30]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b31  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [31]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[31]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b32  (
    .clk(clk100m),
    .d(1'b1),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[32]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[4]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[5]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[6]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[7]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[8]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg30_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(1'b1),
    .reset(~\U_AHB/n71 ),
    .set(1'b0),
    .q(pnumC[9]));  // src/AHB.v(79)
  reg_sr_as_w1 \U_AHB/reg31_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[0]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[1]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[10]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[11]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[12]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[13]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[14]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[15]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[16]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[17]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[18]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[19]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[2]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[20]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[21]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[22]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[23]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[24]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[25]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[26]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b27  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [27]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[27]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b28  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [28]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[28]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b29  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [29]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[29]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[3]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b30  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [30]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[30]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b31  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [31]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[31]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b32  (
    .clk(clk100m),
    .d(1'b1),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[32]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[4]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[5]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[6]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[7]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[8]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg31_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(1'b1),
    .reset(~\U_AHB/n73 ),
    .set(1'b0),
    .q(pnumD[9]));  // src/AHB.v(80)
  reg_sr_as_w1 \U_AHB/reg32_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[0]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[1]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[10]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[11]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[12]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[13]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[14]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[15]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[16]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[17]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[18]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[19]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[2]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[20]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[21]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[22]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[23]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[24]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[25]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[26]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b27  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [27]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[27]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b28  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [28]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[28]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b29  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [29]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[29]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[3]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b30  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [30]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[30]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b31  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [31]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[31]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b32  (
    .clk(clk100m),
    .d(1'b1),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[32]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[4]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[5]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[6]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[7]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[8]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg32_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(1'b1),
    .reset(~\U_AHB/n75 ),
    .set(1'b0),
    .q(pnumE[9]));  // src/AHB.v(81)
  reg_sr_as_w1 \U_AHB/reg33_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[0]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[1]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[10]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[11]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[12]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[13]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[14]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[15]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[16]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[17]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[18]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[19]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[2]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[20]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[21]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[22]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[23]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[24]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[25]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[26]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b27  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [27]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[27]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b28  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [28]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[28]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b29  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [29]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[29]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[3]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b30  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [30]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[30]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b31  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [31]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[31]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b32  (
    .clk(clk100m),
    .d(1'b1),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[32]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[4]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[5]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[6]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[7]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[8]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg33_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(1'b1),
    .reset(~\U_AHB/n77 ),
    .set(1'b0),
    .q(pnumF[9]));  // src/AHB.v(82)
  reg_sr_as_w1 \U_AHB/reg34_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[0]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[1]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[10]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[11]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[12]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[13]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[14]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[15]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[16]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[17]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[18]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[19]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[2]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[20]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[21]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[22]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[23]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[24]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[25]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[26]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b27  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [27]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[27]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b28  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [28]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[28]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b29  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [29]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[29]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[3]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b30  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [30]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[30]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b31  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [31]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[31]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[4]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[5]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[6]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[7]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[8]));  // src/AHB.v(84)
  reg_sr_as_w1 \U_AHB/reg34_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(1'b1),
    .reset(~\U_AHB/n79 ),
    .set(1'b0),
    .q(pwm_start_stop[9]));  // src/AHB.v(84)
  reg_ar_as_w1 \U_AHB/reg35_b0  (
    .clk(clk100m),
    .d(\U_AHB/n118 [0]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [0]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b1  (
    .clk(clk100m),
    .d(\U_AHB/n118 [1]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [1]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b10  (
    .clk(clk100m),
    .d(\U_AHB/n118 [10]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [10]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b11  (
    .clk(clk100m),
    .d(\U_AHB/n118 [11]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [11]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b12  (
    .clk(clk100m),
    .d(\U_AHB/n118 [12]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [12]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b13  (
    .clk(clk100m),
    .d(\U_AHB/n118 [13]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [13]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b14  (
    .clk(clk100m),
    .d(\U_AHB/n118 [14]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [14]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b15  (
    .clk(clk100m),
    .d(\U_AHB/n118 [15]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [15]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b16  (
    .clk(clk100m),
    .d(\U_AHB/n118 [16]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [16]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b17  (
    .clk(clk100m),
    .d(\U_AHB/n118 [17]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [17]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b18  (
    .clk(clk100m),
    .d(\U_AHB/n118 [18]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [18]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b19  (
    .clk(clk100m),
    .d(\U_AHB/n118 [19]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [19]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b2  (
    .clk(clk100m),
    .d(\U_AHB/n118 [2]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [2]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b20  (
    .clk(clk100m),
    .d(\U_AHB/n118 [20]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [20]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b21  (
    .clk(clk100m),
    .d(\U_AHB/n118 [21]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [21]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b22  (
    .clk(clk100m),
    .d(\U_AHB/n118 [22]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [22]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b23  (
    .clk(clk100m),
    .d(\U_AHB/n118 [23]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [23]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b24  (
    .clk(clk100m),
    .d(\U_AHB/n118 [24]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [24]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b25  (
    .clk(clk100m),
    .d(\U_AHB/n118 [25]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [25]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b26  (
    .clk(clk100m),
    .d(\U_AHB/n118 [26]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [26]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b27  (
    .clk(clk100m),
    .d(\U_AHB/n118 [27]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [27]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b28  (
    .clk(clk100m),
    .d(\U_AHB/n118 [28]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [28]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b29  (
    .clk(clk100m),
    .d(\U_AHB/n118 [29]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [29]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b3  (
    .clk(clk100m),
    .d(\U_AHB/n118 [3]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [3]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b30  (
    .clk(clk100m),
    .d(\U_AHB/n118 [30]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [30]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b31  (
    .clk(clk100m),
    .d(\U_AHB/n118 [31]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [31]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b4  (
    .clk(clk100m),
    .d(\U_AHB/n118 [4]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [4]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b5  (
    .clk(clk100m),
    .d(\U_AHB/n118 [5]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [5]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b6  (
    .clk(clk100m),
    .d(\U_AHB/n118 [6]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [6]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b7  (
    .clk(clk100m),
    .d(\U_AHB/n118 [7]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [7]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b8  (
    .clk(clk100m),
    .d(\U_AHB/n118 [8]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [8]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg35_b9  (
    .clk(clk100m),
    .d(\U_AHB/n118 [9]),
    .en(1'b1),
    .reset(1'b0),
    .set(1'b0),
    .q(\U_AHB/h2h_hrdata [9]));  // src/AHB.v(115)
  reg_ar_as_w1 \U_AHB/reg3_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[0]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[1]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[10]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[11]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[12]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[13]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[14]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[15]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[16]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[17]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[18]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[19]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[2]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[20]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[21]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[22]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[23]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[24]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[25]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[26]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[3]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[4]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[5]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[6]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[7]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[8]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg3_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(\U_AHB/n8 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq2[9]));  // src/AHB.v(48)
  reg_ar_as_w1 \U_AHB/reg4_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[0]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[1]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[10]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[11]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[12]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[13]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[14]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[15]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[16]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[17]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[18]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[19]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[2]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[20]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[21]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[22]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[23]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[24]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[25]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[26]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[3]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[4]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[5]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[6]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[7]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[8]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg4_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(\U_AHB/n10 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq3[9]));  // src/AHB.v(49)
  reg_ar_as_w1 \U_AHB/reg5_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[0]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[1]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[10]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[11]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[12]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[13]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[14]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[15]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[16]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[17]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[18]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[19]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[2]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[20]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[21]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[22]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[23]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[24]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[25]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[26]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[3]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[4]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[5]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[6]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[7]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[8]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg5_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(\U_AHB/n12 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq4[9]));  // src/AHB.v(50)
  reg_ar_as_w1 \U_AHB/reg6_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[0]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[1]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[10]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[11]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[12]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[13]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[14]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[15]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[16]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[17]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[18]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[19]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[2]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[20]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[21]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[22]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[23]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[24]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[25]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[26]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[3]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[4]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[5]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[6]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[7]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[8]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg6_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(\U_AHB/n14 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq5[9]));  // src/AHB.v(51)
  reg_ar_as_w1 \U_AHB/reg7_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[0]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[1]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[10]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[11]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[12]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[13]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[14]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[15]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[16]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[17]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[18]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[19]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[2]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[20]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[21]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[22]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[23]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[24]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[25]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[26]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[3]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[4]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[5]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[6]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[7]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[8]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg7_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(\U_AHB/n16 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq6[9]));  // src/AHB.v(52)
  reg_ar_as_w1 \U_AHB/reg8_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[0]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[1]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[10]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[11]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[12]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[13]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[14]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[15]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[16]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[17]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[18]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[19]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[2]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[20]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[21]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[22]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[23]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[24]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[25]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[26]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[3]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[4]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[5]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[6]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[7]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[8]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg8_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(\U_AHB/n18 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq7[9]));  // src/AHB.v(53)
  reg_ar_as_w1 \U_AHB/reg9_b0  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [0]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[0]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b1  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [1]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[1]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b10  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [10]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[10]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b11  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [11]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[11]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b12  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [12]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[12]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b13  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [13]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[13]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b14  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [14]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[14]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b15  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [15]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[15]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b16  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [16]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[16]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b17  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [17]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[17]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b18  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [18]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[18]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b19  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [19]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[19]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b2  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [2]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[2]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b20  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [20]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[20]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b21  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [21]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[21]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b22  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [22]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[22]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b23  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [23]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[23]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b24  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [24]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[24]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b25  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [25]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[25]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b26  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [26]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[26]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b3  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [3]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[3]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b4  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [4]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[4]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b5  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [5]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[5]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b6  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [6]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[6]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b7  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [7]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[7]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b8  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [8]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[8]));  // src/AHB.v(54)
  reg_ar_as_w1 \U_AHB/reg9_b9  (
    .clk(clk100m),
    .d(\U_AHB/h2h_hwdata [9]),
    .en(\U_AHB/n20 ),
    .reset(1'b0),
    .set(1'b0),
    .q(freq8[9]));  // src/AHB.v(54)
  and \U_AHB/sel0_b0/and_b0_0  (\U_AHB/sel0_b0/B0 , \U_AHB/h2h_hrdata [0], \U_AHB/n113 );
  and \U_AHB/sel0_b0/and_b0_1  (\U_AHB/sel0_b0/B1 , pnumcntA[0], \U_AHB/n111 );
  and \U_AHB/sel0_b0/and_b0_10  (\U_AHB/sel0_b0/B10 , pnumcnt1[0], \U_AHB/n84 );
  and \U_AHB/sel0_b0/and_b0_11  (\U_AHB/sel0_b0/B11 , pnumcnt0[0], \U_AHB/h2h_haddr [2]);
  and \U_AHB/sel0_b0/and_b0_2  (\U_AHB/sel0_b0/B2 , pnumcnt9[0], \U_AHB/n108 );
  and \U_AHB/sel0_b0/and_b0_3  (\U_AHB/sel0_b0/B3 , pnumcnt8[0], \U_AHB/n105 );
  and \U_AHB/sel0_b0/and_b0_4  (\U_AHB/sel0_b0/B4 , pnumcnt7[0], \U_AHB/n102 );
  and \U_AHB/sel0_b0/and_b0_5  (\U_AHB/sel0_b0/B5 , pnumcnt6[0], \U_AHB/n99 );
  and \U_AHB/sel0_b0/and_b0_6  (\U_AHB/sel0_b0/B6 , pnumcnt5[0], \U_AHB/n96 );
  and \U_AHB/sel0_b0/and_b0_7  (\U_AHB/sel0_b0/B7 , pnumcnt4[0], \U_AHB/n93 );
  and \U_AHB/sel0_b0/and_b0_8  (\U_AHB/sel0_b0/B8 , pnumcnt3[0], \U_AHB/n90 );
  and \U_AHB/sel0_b0/and_b0_9  (\U_AHB/sel0_b0/B9 , pnumcnt2[0], \U_AHB/n87 );
  or \U_AHB/sel0_b0/or_B0_or_B1_B2_o  (\U_AHB/sel0_b0/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b0/B0 , \U_AHB/sel0_b0/or_B1_B2_o );
  or \U_AHB/sel0_b0/or_B10_B11  (\U_AHB/sel0_b0/or_B10_B11_o , \U_AHB/sel0_b0/B10 , \U_AHB/sel0_b0/B11 );
  or \U_AHB/sel0_b0/or_B1_B2  (\U_AHB/sel0_b0/or_B1_B2_o , \U_AHB/sel0_b0/B1 , \U_AHB/sel0_b0/B2 );
  or \U_AHB/sel0_b0/or_B3_or_B4_B5_o  (\U_AHB/sel0_b0/or_B3_or_B4_B5_o_o , \U_AHB/sel0_b0/B3 , \U_AHB/sel0_b0/or_B4_B5_o );
  or \U_AHB/sel0_b0/or_B4_B5  (\U_AHB/sel0_b0/or_B4_B5_o , \U_AHB/sel0_b0/B4 , \U_AHB/sel0_b0/B5 );
  or \U_AHB/sel0_b0/or_B6_or_B7_B8_o  (\U_AHB/sel0_b0/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b0/B6 , \U_AHB/sel0_b0/or_B7_B8_o );
  or \U_AHB/sel0_b0/or_B7_B8  (\U_AHB/sel0_b0/or_B7_B8_o , \U_AHB/sel0_b0/B7 , \U_AHB/sel0_b0/B8 );
  or \U_AHB/sel0_b0/or_B9_or_B10_B11_o  (\U_AHB/sel0_b0/or_B9_or_B10_B11_o_o , \U_AHB/sel0_b0/B9 , \U_AHB/sel0_b0/or_B10_B11_o );
  or \U_AHB/sel0_b0/or_or_B0_or_B1_B2_o_  (\U_AHB/sel0_b0/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b0/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b0/or_B3_or_B4_B5_o_o );
  or \U_AHB/sel0_b0/or_or_B6_or_B7_B8_o_  (\U_AHB/sel0_b0/or_or_B6_or_B7_B8_o__o , \U_AHB/sel0_b0/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b0/or_B9_or_B10_B11_o_o );
  or \U_AHB/sel0_b0/or_or_or_B0_or_B1_B2  (\U_AHB/n114 [0], \U_AHB/sel0_b0/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b0/or_or_B6_or_B7_B8_o__o );
  and \U_AHB/sel0_b1/and_b0_0  (\U_AHB/sel0_b1/B0 , \U_AHB/h2h_hrdata [1], \U_AHB/n113 );
  and \U_AHB/sel0_b1/and_b0_1  (\U_AHB/sel0_b1/B1 , pnumcntA[1], \U_AHB/n111 );
  and \U_AHB/sel0_b1/and_b0_10  (\U_AHB/sel0_b1/B10 , pnumcnt1[1], \U_AHB/n84 );
  and \U_AHB/sel0_b1/and_b0_11  (\U_AHB/sel0_b1/B11 , pnumcnt0[1], \U_AHB/h2h_haddr [2]);
  and \U_AHB/sel0_b1/and_b0_2  (\U_AHB/sel0_b1/B2 , pnumcnt9[1], \U_AHB/n108 );
  and \U_AHB/sel0_b1/and_b0_3  (\U_AHB/sel0_b1/B3 , pnumcnt8[1], \U_AHB/n105 );
  and \U_AHB/sel0_b1/and_b0_4  (\U_AHB/sel0_b1/B4 , pnumcnt7[1], \U_AHB/n102 );
  and \U_AHB/sel0_b1/and_b0_5  (\U_AHB/sel0_b1/B5 , pnumcnt6[1], \U_AHB/n99 );
  and \U_AHB/sel0_b1/and_b0_6  (\U_AHB/sel0_b1/B6 , pnumcnt5[1], \U_AHB/n96 );
  and \U_AHB/sel0_b1/and_b0_7  (\U_AHB/sel0_b1/B7 , pnumcnt4[1], \U_AHB/n93 );
  and \U_AHB/sel0_b1/and_b0_8  (\U_AHB/sel0_b1/B8 , pnumcnt3[1], \U_AHB/n90 );
  and \U_AHB/sel0_b1/and_b0_9  (\U_AHB/sel0_b1/B9 , pnumcnt2[1], \U_AHB/n87 );
  or \U_AHB/sel0_b1/or_B0_or_B1_B2_o  (\U_AHB/sel0_b1/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b1/B0 , \U_AHB/sel0_b1/or_B1_B2_o );
  or \U_AHB/sel0_b1/or_B10_B11  (\U_AHB/sel0_b1/or_B10_B11_o , \U_AHB/sel0_b1/B10 , \U_AHB/sel0_b1/B11 );
  or \U_AHB/sel0_b1/or_B1_B2  (\U_AHB/sel0_b1/or_B1_B2_o , \U_AHB/sel0_b1/B1 , \U_AHB/sel0_b1/B2 );
  or \U_AHB/sel0_b1/or_B3_or_B4_B5_o  (\U_AHB/sel0_b1/or_B3_or_B4_B5_o_o , \U_AHB/sel0_b1/B3 , \U_AHB/sel0_b1/or_B4_B5_o );
  or \U_AHB/sel0_b1/or_B4_B5  (\U_AHB/sel0_b1/or_B4_B5_o , \U_AHB/sel0_b1/B4 , \U_AHB/sel0_b1/B5 );
  or \U_AHB/sel0_b1/or_B6_or_B7_B8_o  (\U_AHB/sel0_b1/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b1/B6 , \U_AHB/sel0_b1/or_B7_B8_o );
  or \U_AHB/sel0_b1/or_B7_B8  (\U_AHB/sel0_b1/or_B7_B8_o , \U_AHB/sel0_b1/B7 , \U_AHB/sel0_b1/B8 );
  or \U_AHB/sel0_b1/or_B9_or_B10_B11_o  (\U_AHB/sel0_b1/or_B9_or_B10_B11_o_o , \U_AHB/sel0_b1/B9 , \U_AHB/sel0_b1/or_B10_B11_o );
  or \U_AHB/sel0_b1/or_or_B0_or_B1_B2_o_  (\U_AHB/sel0_b1/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b1/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b1/or_B3_or_B4_B5_o_o );
  or \U_AHB/sel0_b1/or_or_B6_or_B7_B8_o_  (\U_AHB/sel0_b1/or_or_B6_or_B7_B8_o__o , \U_AHB/sel0_b1/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b1/or_B9_or_B10_B11_o_o );
  or \U_AHB/sel0_b1/or_or_or_B0_or_B1_B2  (\U_AHB/n114 [1], \U_AHB/sel0_b1/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b1/or_or_B6_or_B7_B8_o__o );
  and \U_AHB/sel0_b10/and_b0_0  (\U_AHB/sel0_b10/B0 , \U_AHB/h2h_hrdata [10], \U_AHB/n113 );
  and \U_AHB/sel0_b10/and_b0_1  (\U_AHB/sel0_b10/B1 , pnumcntA[10], \U_AHB/n111 );
  and \U_AHB/sel0_b10/and_b0_10  (\U_AHB/sel0_b10/B10 , pnumcnt1[10], \U_AHB/n84 );
  and \U_AHB/sel0_b10/and_b0_11  (\U_AHB/sel0_b10/B11 , pnumcnt0[10], \U_AHB/h2h_haddr [2]);
  and \U_AHB/sel0_b10/and_b0_2  (\U_AHB/sel0_b10/B2 , pnumcnt9[10], \U_AHB/n108 );
  and \U_AHB/sel0_b10/and_b0_3  (\U_AHB/sel0_b10/B3 , pnumcnt8[10], \U_AHB/n105 );
  and \U_AHB/sel0_b10/and_b0_4  (\U_AHB/sel0_b10/B4 , pnumcnt7[10], \U_AHB/n102 );
  and \U_AHB/sel0_b10/and_b0_5  (\U_AHB/sel0_b10/B5 , pnumcnt6[10], \U_AHB/n99 );
  and \U_AHB/sel0_b10/and_b0_6  (\U_AHB/sel0_b10/B6 , pnumcnt5[10], \U_AHB/n96 );
  and \U_AHB/sel0_b10/and_b0_7  (\U_AHB/sel0_b10/B7 , pnumcnt4[10], \U_AHB/n93 );
  and \U_AHB/sel0_b10/and_b0_8  (\U_AHB/sel0_b10/B8 , pnumcnt3[10], \U_AHB/n90 );
  and \U_AHB/sel0_b10/and_b0_9  (\U_AHB/sel0_b10/B9 , pnumcnt2[10], \U_AHB/n87 );
  or \U_AHB/sel0_b10/or_B0_or_B1_B2_o  (\U_AHB/sel0_b10/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b10/B0 , \U_AHB/sel0_b10/or_B1_B2_o );
  or \U_AHB/sel0_b10/or_B10_B11  (\U_AHB/sel0_b10/or_B10_B11_o , \U_AHB/sel0_b10/B10 , \U_AHB/sel0_b10/B11 );
  or \U_AHB/sel0_b10/or_B1_B2  (\U_AHB/sel0_b10/or_B1_B2_o , \U_AHB/sel0_b10/B1 , \U_AHB/sel0_b10/B2 );
  or \U_AHB/sel0_b10/or_B3_or_B4_B5_o  (\U_AHB/sel0_b10/or_B3_or_B4_B5_o_o , \U_AHB/sel0_b10/B3 , \U_AHB/sel0_b10/or_B4_B5_o );
  or \U_AHB/sel0_b10/or_B4_B5  (\U_AHB/sel0_b10/or_B4_B5_o , \U_AHB/sel0_b10/B4 , \U_AHB/sel0_b10/B5 );
  or \U_AHB/sel0_b10/or_B6_or_B7_B8_o  (\U_AHB/sel0_b10/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b10/B6 , \U_AHB/sel0_b10/or_B7_B8_o );
  or \U_AHB/sel0_b10/or_B7_B8  (\U_AHB/sel0_b10/or_B7_B8_o , \U_AHB/sel0_b10/B7 , \U_AHB/sel0_b10/B8 );
  or \U_AHB/sel0_b10/or_B9_or_B10_B11_o  (\U_AHB/sel0_b10/or_B9_or_B10_B11_o_o , \U_AHB/sel0_b10/B9 , \U_AHB/sel0_b10/or_B10_B11_o );
  or \U_AHB/sel0_b10/or_or_B0_or_B1_B2_o_  (\U_AHB/sel0_b10/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b10/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b10/or_B3_or_B4_B5_o_o );
  or \U_AHB/sel0_b10/or_or_B6_or_B7_B8_o_  (\U_AHB/sel0_b10/or_or_B6_or_B7_B8_o__o , \U_AHB/sel0_b10/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b10/or_B9_or_B10_B11_o_o );
  or \U_AHB/sel0_b10/or_or_or_B0_or_B1_B2  (\U_AHB/n114 [10], \U_AHB/sel0_b10/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b10/or_or_B6_or_B7_B8_o__o );
  and \U_AHB/sel0_b11/and_b0_0  (\U_AHB/sel0_b11/B0 , \U_AHB/h2h_hrdata [11], \U_AHB/n113 );
  and \U_AHB/sel0_b11/and_b0_1  (\U_AHB/sel0_b11/B1 , pnumcntA[11], \U_AHB/n111 );
  and \U_AHB/sel0_b11/and_b0_10  (\U_AHB/sel0_b11/B10 , pnumcnt1[11], \U_AHB/n84 );
  and \U_AHB/sel0_b11/and_b0_11  (\U_AHB/sel0_b11/B11 , pnumcnt0[11], \U_AHB/h2h_haddr [2]);
  and \U_AHB/sel0_b11/and_b0_2  (\U_AHB/sel0_b11/B2 , pnumcnt9[11], \U_AHB/n108 );
  and \U_AHB/sel0_b11/and_b0_3  (\U_AHB/sel0_b11/B3 , pnumcnt8[11], \U_AHB/n105 );
  and \U_AHB/sel0_b11/and_b0_4  (\U_AHB/sel0_b11/B4 , pnumcnt7[11], \U_AHB/n102 );
  and \U_AHB/sel0_b11/and_b0_5  (\U_AHB/sel0_b11/B5 , pnumcnt6[11], \U_AHB/n99 );
  and \U_AHB/sel0_b11/and_b0_6  (\U_AHB/sel0_b11/B6 , pnumcnt5[11], \U_AHB/n96 );
  and \U_AHB/sel0_b11/and_b0_7  (\U_AHB/sel0_b11/B7 , pnumcnt4[11], \U_AHB/n93 );
  and \U_AHB/sel0_b11/and_b0_8  (\U_AHB/sel0_b11/B8 , pnumcnt3[11], \U_AHB/n90 );
  and \U_AHB/sel0_b11/and_b0_9  (\U_AHB/sel0_b11/B9 , pnumcnt2[11], \U_AHB/n87 );
  or \U_AHB/sel0_b11/or_B0_or_B1_B2_o  (\U_AHB/sel0_b11/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b11/B0 , \U_AHB/sel0_b11/or_B1_B2_o );
  or \U_AHB/sel0_b11/or_B10_B11  (\U_AHB/sel0_b11/or_B10_B11_o , \U_AHB/sel0_b11/B10 , \U_AHB/sel0_b11/B11 );
  or \U_AHB/sel0_b11/or_B1_B2  (\U_AHB/sel0_b11/or_B1_B2_o , \U_AHB/sel0_b11/B1 , \U_AHB/sel0_b11/B2 );
  or \U_AHB/sel0_b11/or_B3_or_B4_B5_o  (\U_AHB/sel0_b11/or_B3_or_B4_B5_o_o , \U_AHB/sel0_b11/B3 , \U_AHB/sel0_b11/or_B4_B5_o );
  or \U_AHB/sel0_b11/or_B4_B5  (\U_AHB/sel0_b11/or_B4_B5_o , \U_AHB/sel0_b11/B4 , \U_AHB/sel0_b11/B5 );
  or \U_AHB/sel0_b11/or_B6_or_B7_B8_o  (\U_AHB/sel0_b11/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b11/B6 , \U_AHB/sel0_b11/or_B7_B8_o );
  or \U_AHB/sel0_b11/or_B7_B8  (\U_AHB/sel0_b11/or_B7_B8_o , \U_AHB/sel0_b11/B7 , \U_AHB/sel0_b11/B8 );
  or \U_AHB/sel0_b11/or_B9_or_B10_B11_o  (\U_AHB/sel0_b11/or_B9_or_B10_B11_o_o , \U_AHB/sel0_b11/B9 , \U_AHB/sel0_b11/or_B10_B11_o );
  or \U_AHB/sel0_b11/or_or_B0_or_B1_B2_o_  (\U_AHB/sel0_b11/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b11/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b11/or_B3_or_B4_B5_o_o );
  or \U_AHB/sel0_b11/or_or_B6_or_B7_B8_o_  (\U_AHB/sel0_b11/or_or_B6_or_B7_B8_o__o , \U_AHB/sel0_b11/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b11/or_B9_or_B10_B11_o_o );
  or \U_AHB/sel0_b11/or_or_or_B0_or_B1_B2  (\U_AHB/n114 [11], \U_AHB/sel0_b11/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b11/or_or_B6_or_B7_B8_o__o );
  and \U_AHB/sel0_b12/and_b0_0  (\U_AHB/sel0_b12/B0 , \U_AHB/h2h_hrdata [12], \U_AHB/n113 );
  and \U_AHB/sel0_b12/and_b0_1  (\U_AHB/sel0_b12/B1 , pnumcntA[12], \U_AHB/n111 );
  and \U_AHB/sel0_b12/and_b0_10  (\U_AHB/sel0_b12/B10 , pnumcnt1[12], \U_AHB/n84 );
  and \U_AHB/sel0_b12/and_b0_11  (\U_AHB/sel0_b12/B11 , pnumcnt0[12], \U_AHB/h2h_haddr [2]);
  and \U_AHB/sel0_b12/and_b0_2  (\U_AHB/sel0_b12/B2 , pnumcnt9[12], \U_AHB/n108 );
  and \U_AHB/sel0_b12/and_b0_3  (\U_AHB/sel0_b12/B3 , pnumcnt8[12], \U_AHB/n105 );
  and \U_AHB/sel0_b12/and_b0_4  (\U_AHB/sel0_b12/B4 , pnumcnt7[12], \U_AHB/n102 );
  and \U_AHB/sel0_b12/and_b0_5  (\U_AHB/sel0_b12/B5 , pnumcnt6[12], \U_AHB/n99 );
  and \U_AHB/sel0_b12/and_b0_6  (\U_AHB/sel0_b12/B6 , pnumcnt5[12], \U_AHB/n96 );
  and \U_AHB/sel0_b12/and_b0_7  (\U_AHB/sel0_b12/B7 , pnumcnt4[12], \U_AHB/n93 );
  and \U_AHB/sel0_b12/and_b0_8  (\U_AHB/sel0_b12/B8 , pnumcnt3[12], \U_AHB/n90 );
  and \U_AHB/sel0_b12/and_b0_9  (\U_AHB/sel0_b12/B9 , pnumcnt2[12], \U_AHB/n87 );
  or \U_AHB/sel0_b12/or_B0_or_B1_B2_o  (\U_AHB/sel0_b12/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b12/B0 , \U_AHB/sel0_b12/or_B1_B2_o );
  or \U_AHB/sel0_b12/or_B10_B11  (\U_AHB/sel0_b12/or_B10_B11_o , \U_AHB/sel0_b12/B10 , \U_AHB/sel0_b12/B11 );
  or \U_AHB/sel0_b12/or_B1_B2  (\U_AHB/sel0_b12/or_B1_B2_o , \U_AHB/sel0_b12/B1 , \U_AHB/sel0_b12/B2 );
  or \U_AHB/sel0_b12/or_B3_or_B4_B5_o  (\U_AHB/sel0_b12/or_B3_or_B4_B5_o_o , \U_AHB/sel0_b12/B3 , \U_AHB/sel0_b12/or_B4_B5_o );
  or \U_AHB/sel0_b12/or_B4_B5  (\U_AHB/sel0_b12/or_B4_B5_o , \U_AHB/sel0_b12/B4 , \U_AHB/sel0_b12/B5 );
  or \U_AHB/sel0_b12/or_B6_or_B7_B8_o  (\U_AHB/sel0_b12/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b12/B6 , \U_AHB/sel0_b12/or_B7_B8_o );
  or \U_AHB/sel0_b12/or_B7_B8  (\U_AHB/sel0_b12/or_B7_B8_o , \U_AHB/sel0_b12/B7 , \U_AHB/sel0_b12/B8 );
  or \U_AHB/sel0_b12/or_B9_or_B10_B11_o  (\U_AHB/sel0_b12/or_B9_or_B10_B11_o_o , \U_AHB/sel0_b12/B9 , \U_AHB/sel0_b12/or_B10_B11_o );
  or \U_AHB/sel0_b12/or_or_B0_or_B1_B2_o_  (\U_AHB/sel0_b12/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b12/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b12/or_B3_or_B4_B5_o_o );
  or \U_AHB/sel0_b12/or_or_B6_or_B7_B8_o_  (\U_AHB/sel0_b12/or_or_B6_or_B7_B8_o__o , \U_AHB/sel0_b12/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b12/or_B9_or_B10_B11_o_o );
  or \U_AHB/sel0_b12/or_or_or_B0_or_B1_B2  (\U_AHB/n114 [12], \U_AHB/sel0_b12/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b12/or_or_B6_or_B7_B8_o__o );
  and \U_AHB/sel0_b13/and_b0_0  (\U_AHB/sel0_b13/B0 , \U_AHB/h2h_hrdata [13], \U_AHB/n113 );
  and \U_AHB/sel0_b13/and_b0_1  (\U_AHB/sel0_b13/B1 , pnumcntA[13], \U_AHB/n111 );
  and \U_AHB/sel0_b13/and_b0_10  (\U_AHB/sel0_b13/B10 , pnumcnt1[13], \U_AHB/n84 );
  and \U_AHB/sel0_b13/and_b0_11  (\U_AHB/sel0_b13/B11 , pnumcnt0[13], \U_AHB/h2h_haddr [2]);
  and \U_AHB/sel0_b13/and_b0_2  (\U_AHB/sel0_b13/B2 , pnumcnt9[13], \U_AHB/n108 );
  and \U_AHB/sel0_b13/and_b0_3  (\U_AHB/sel0_b13/B3 , pnumcnt8[13], \U_AHB/n105 );
  and \U_AHB/sel0_b13/and_b0_4  (\U_AHB/sel0_b13/B4 , pnumcnt7[13], \U_AHB/n102 );
  and \U_AHB/sel0_b13/and_b0_5  (\U_AHB/sel0_b13/B5 , pnumcnt6[13], \U_AHB/n99 );
  and \U_AHB/sel0_b13/and_b0_6  (\U_AHB/sel0_b13/B6 , pnumcnt5[13], \U_AHB/n96 );
  and \U_AHB/sel0_b13/and_b0_7  (\U_AHB/sel0_b13/B7 , pnumcnt4[13], \U_AHB/n93 );
  and \U_AHB/sel0_b13/and_b0_8  (\U_AHB/sel0_b13/B8 , pnumcnt3[13], \U_AHB/n90 );
  and \U_AHB/sel0_b13/and_b0_9  (\U_AHB/sel0_b13/B9 , pnumcnt2[13], \U_AHB/n87 );
  or \U_AHB/sel0_b13/or_B0_or_B1_B2_o  (\U_AHB/sel0_b13/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b13/B0 , \U_AHB/sel0_b13/or_B1_B2_o );
  or \U_AHB/sel0_b13/or_B10_B11  (\U_AHB/sel0_b13/or_B10_B11_o , \U_AHB/sel0_b13/B10 , \U_AHB/sel0_b13/B11 );
  or \U_AHB/sel0_b13/or_B1_B2  (\U_AHB/sel0_b13/or_B1_B2_o , \U_AHB/sel0_b13/B1 , \U_AHB/sel0_b13/B2 );
  or \U_AHB/sel0_b13/or_B3_or_B4_B5_o  (\U_AHB/sel0_b13/or_B3_or_B4_B5_o_o , \U_AHB/sel0_b13/B3 , \U_AHB/sel0_b13/or_B4_B5_o );
  or \U_AHB/sel0_b13/or_B4_B5  (\U_AHB/sel0_b13/or_B4_B5_o , \U_AHB/sel0_b13/B4 , \U_AHB/sel0_b13/B5 );
  or \U_AHB/sel0_b13/or_B6_or_B7_B8_o  (\U_AHB/sel0_b13/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b13/B6 , \U_AHB/sel0_b13/or_B7_B8_o );
  or \U_AHB/sel0_b13/or_B7_B8  (\U_AHB/sel0_b13/or_B7_B8_o , \U_AHB/sel0_b13/B7 , \U_AHB/sel0_b13/B8 );
  or \U_AHB/sel0_b13/or_B9_or_B10_B11_o  (\U_AHB/sel0_b13/or_B9_or_B10_B11_o_o , \U_AHB/sel0_b13/B9 , \U_AHB/sel0_b13/or_B10_B11_o );
  or \U_AHB/sel0_b13/or_or_B0_or_B1_B2_o_  (\U_AHB/sel0_b13/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b13/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b13/or_B3_or_B4_B5_o_o );
  or \U_AHB/sel0_b13/or_or_B6_or_B7_B8_o_  (\U_AHB/sel0_b13/or_or_B6_or_B7_B8_o__o , \U_AHB/sel0_b13/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b13/or_B9_or_B10_B11_o_o );
  or \U_AHB/sel0_b13/or_or_or_B0_or_B1_B2  (\U_AHB/n114 [13], \U_AHB/sel0_b13/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b13/or_or_B6_or_B7_B8_o__o );
  and \U_AHB/sel0_b14/and_b0_0  (\U_AHB/sel0_b14/B0 , \U_AHB/h2h_hrdata [14], \U_AHB/n113 );
  and \U_AHB/sel0_b14/and_b0_1  (\U_AHB/sel0_b14/B1 , pnumcntA[14], \U_AHB/n111 );
  and \U_AHB/sel0_b14/and_b0_10  (\U_AHB/sel0_b14/B10 , pnumcnt1[14], \U_AHB/n84 );
  and \U_AHB/sel0_b14/and_b0_11  (\U_AHB/sel0_b14/B11 , pnumcnt0[14], \U_AHB/h2h_haddr [2]);
  and \U_AHB/sel0_b14/and_b0_2  (\U_AHB/sel0_b14/B2 , pnumcnt9[14], \U_AHB/n108 );
  and \U_AHB/sel0_b14/and_b0_3  (\U_AHB/sel0_b14/B3 , pnumcnt8[14], \U_AHB/n105 );
  and \U_AHB/sel0_b14/and_b0_4  (\U_AHB/sel0_b14/B4 , pnumcnt7[14], \U_AHB/n102 );
  and \U_AHB/sel0_b14/and_b0_5  (\U_AHB/sel0_b14/B5 , pnumcnt6[14], \U_AHB/n99 );
  and \U_AHB/sel0_b14/and_b0_6  (\U_AHB/sel0_b14/B6 , pnumcnt5[14], \U_AHB/n96 );
  and \U_AHB/sel0_b14/and_b0_7  (\U_AHB/sel0_b14/B7 , pnumcnt4[14], \U_AHB/n93 );
  and \U_AHB/sel0_b14/and_b0_8  (\U_AHB/sel0_b14/B8 , pnumcnt3[14], \U_AHB/n90 );
  and \U_AHB/sel0_b14/and_b0_9  (\U_AHB/sel0_b14/B9 , pnumcnt2[14], \U_AHB/n87 );
  or \U_AHB/sel0_b14/or_B0_or_B1_B2_o  (\U_AHB/sel0_b14/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b14/B0 , \U_AHB/sel0_b14/or_B1_B2_o );
  or \U_AHB/sel0_b14/or_B10_B11  (\U_AHB/sel0_b14/or_B10_B11_o , \U_AHB/sel0_b14/B10 , \U_AHB/sel0_b14/B11 );
  or \U_AHB/sel0_b14/or_B1_B2  (\U_AHB/sel0_b14/or_B1_B2_o , \U_AHB/sel0_b14/B1 , \U_AHB/sel0_b14/B2 );
  or \U_AHB/sel0_b14/or_B3_or_B4_B5_o  (\U_AHB/sel0_b14/or_B3_or_B4_B5_o_o , \U_AHB/sel0_b14/B3 , \U_AHB/sel0_b14/or_B4_B5_o );
  or \U_AHB/sel0_b14/or_B4_B5  (\U_AHB/sel0_b14/or_B4_B5_o , \U_AHB/sel0_b14/B4 , \U_AHB/sel0_b14/B5 );
  or \U_AHB/sel0_b14/or_B6_or_B7_B8_o  (\U_AHB/sel0_b14/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b14/B6 , \U_AHB/sel0_b14/or_B7_B8_o );
  or \U_AHB/sel0_b14/or_B7_B8  (\U_AHB/sel0_b14/or_B7_B8_o , \U_AHB/sel0_b14/B7 , \U_AHB/sel0_b14/B8 );
  or \U_AHB/sel0_b14/or_B9_or_B10_B11_o  (\U_AHB/sel0_b14/or_B9_or_B10_B11_o_o , \U_AHB/sel0_b14/B9 , \U_AHB/sel0_b14/or_B10_B11_o );
  or \U_AHB/sel0_b14/or_or_B0_or_B1_B2_o_  (\U_AHB/sel0_b14/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b14/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b14/or_B3_or_B4_B5_o_o );
  or \U_AHB/sel0_b14/or_or_B6_or_B7_B8_o_  (\U_AHB/sel0_b14/or_or_B6_or_B7_B8_o__o , \U_AHB/sel0_b14/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b14/or_B9_or_B10_B11_o_o );
  or \U_AHB/sel0_b14/or_or_or_B0_or_B1_B2  (\U_AHB/n114 [14], \U_AHB/sel0_b14/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b14/or_or_B6_or_B7_B8_o__o );
  and \U_AHB/sel0_b15/and_b0_0  (\U_AHB/sel0_b15/B0 , \U_AHB/h2h_hrdata [15], \U_AHB/n113 );
  and \U_AHB/sel0_b15/and_b0_1  (\U_AHB/sel0_b15/B1 , pnumcntA[15], \U_AHB/n111 );
  and \U_AHB/sel0_b15/and_b0_10  (\U_AHB/sel0_b15/B10 , pnumcnt1[15], \U_AHB/n84 );
  and \U_AHB/sel0_b15/and_b0_11  (\U_AHB/sel0_b15/B11 , pnumcnt0[15], \U_AHB/h2h_haddr [2]);
  and \U_AHB/sel0_b15/and_b0_2  (\U_AHB/sel0_b15/B2 , pnumcnt9[15], \U_AHB/n108 );
  and \U_AHB/sel0_b15/and_b0_3  (\U_AHB/sel0_b15/B3 , pnumcnt8[15], \U_AHB/n105 );
  and \U_AHB/sel0_b15/and_b0_4  (\U_AHB/sel0_b15/B4 , pnumcnt7[15], \U_AHB/n102 );
  and \U_AHB/sel0_b15/and_b0_5  (\U_AHB/sel0_b15/B5 , pnumcnt6[15], \U_AHB/n99 );
  and \U_AHB/sel0_b15/and_b0_6  (\U_AHB/sel0_b15/B6 , pnumcnt5[15], \U_AHB/n96 );
  and \U_AHB/sel0_b15/and_b0_7  (\U_AHB/sel0_b15/B7 , pnumcnt4[15], \U_AHB/n93 );
  and \U_AHB/sel0_b15/and_b0_8  (\U_AHB/sel0_b15/B8 , pnumcnt3[15], \U_AHB/n90 );
  and \U_AHB/sel0_b15/and_b0_9  (\U_AHB/sel0_b15/B9 , pnumcnt2[15], \U_AHB/n87 );
  or \U_AHB/sel0_b15/or_B0_or_B1_B2_o  (\U_AHB/sel0_b15/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b15/B0 , \U_AHB/sel0_b15/or_B1_B2_o );
  or \U_AHB/sel0_b15/or_B10_B11  (\U_AHB/sel0_b15/or_B10_B11_o , \U_AHB/sel0_b15/B10 , \U_AHB/sel0_b15/B11 );
  or \U_AHB/sel0_b15/or_B1_B2  (\U_AHB/sel0_b15/or_B1_B2_o , \U_AHB/sel0_b15/B1 , \U_AHB/sel0_b15/B2 );
  or \U_AHB/sel0_b15/or_B3_or_B4_B5_o  (\U_AHB/sel0_b15/or_B3_or_B4_B5_o_o , \U_AHB/sel0_b15/B3 , \U_AHB/sel0_b15/or_B4_B5_o );
  or \U_AHB/sel0_b15/or_B4_B5  (\U_AHB/sel0_b15/or_B4_B5_o , \U_AHB/sel0_b15/B4 , \U_AHB/sel0_b15/B5 );
  or \U_AHB/sel0_b15/or_B6_or_B7_B8_o  (\U_AHB/sel0_b15/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b15/B6 , \U_AHB/sel0_b15/or_B7_B8_o );
  or \U_AHB/sel0_b15/or_B7_B8  (\U_AHB/sel0_b15/or_B7_B8_o , \U_AHB/sel0_b15/B7 , \U_AHB/sel0_b15/B8 );
  or \U_AHB/sel0_b15/or_B9_or_B10_B11_o  (\U_AHB/sel0_b15/or_B9_or_B10_B11_o_o , \U_AHB/sel0_b15/B9 , \U_AHB/sel0_b15/or_B10_B11_o );
  or \U_AHB/sel0_b15/or_or_B0_or_B1_B2_o_  (\U_AHB/sel0_b15/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b15/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b15/or_B3_or_B4_B5_o_o );
  or \U_AHB/sel0_b15/or_or_B6_or_B7_B8_o_  (\U_AHB/sel0_b15/or_or_B6_or_B7_B8_o__o , \U_AHB/sel0_b15/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b15/or_B9_or_B10_B11_o_o );
  or \U_AHB/sel0_b15/or_or_or_B0_or_B1_B2  (\U_AHB/n114 [15], \U_AHB/sel0_b15/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b15/or_or_B6_or_B7_B8_o__o );
  and \U_AHB/sel0_b16/and_b0_0  (\U_AHB/sel0_b16/B0 , \U_AHB/h2h_hrdata [16], \U_AHB/n113 );
  and \U_AHB/sel0_b16/and_b0_1  (\U_AHB/sel0_b16/B1 , pnumcntA[16], \U_AHB/n111 );
  and \U_AHB/sel0_b16/and_b0_10  (\U_AHB/sel0_b16/B10 , pnumcnt1[16], \U_AHB/n84 );
  and \U_AHB/sel0_b16/and_b0_11  (\U_AHB/sel0_b16/B11 , pnumcnt0[16], \U_AHB/h2h_haddr [2]);
  and \U_AHB/sel0_b16/and_b0_2  (\U_AHB/sel0_b16/B2 , pnumcnt9[16], \U_AHB/n108 );
  and \U_AHB/sel0_b16/and_b0_3  (\U_AHB/sel0_b16/B3 , pnumcnt8[16], \U_AHB/n105 );
  and \U_AHB/sel0_b16/and_b0_4  (\U_AHB/sel0_b16/B4 , pnumcnt7[16], \U_AHB/n102 );
  and \U_AHB/sel0_b16/and_b0_5  (\U_AHB/sel0_b16/B5 , pnumcnt6[16], \U_AHB/n99 );
  and \U_AHB/sel0_b16/and_b0_6  (\U_AHB/sel0_b16/B6 , pnumcnt5[16], \U_AHB/n96 );
  and \U_AHB/sel0_b16/and_b0_7  (\U_AHB/sel0_b16/B7 , pnumcnt4[16], \U_AHB/n93 );
  and \U_AHB/sel0_b16/and_b0_8  (\U_AHB/sel0_b16/B8 , pnumcnt3[16], \U_AHB/n90 );
  and \U_AHB/sel0_b16/and_b0_9  (\U_AHB/sel0_b16/B9 , pnumcnt2[16], \U_AHB/n87 );
  or \U_AHB/sel0_b16/or_B0_or_B1_B2_o  (\U_AHB/sel0_b16/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b16/B0 , \U_AHB/sel0_b16/or_B1_B2_o );
  or \U_AHB/sel0_b16/or_B10_B11  (\U_AHB/sel0_b16/or_B10_B11_o , \U_AHB/sel0_b16/B10 , \U_AHB/sel0_b16/B11 );
  or \U_AHB/sel0_b16/or_B1_B2  (\U_AHB/sel0_b16/or_B1_B2_o , \U_AHB/sel0_b16/B1 , \U_AHB/sel0_b16/B2 );
  or \U_AHB/sel0_b16/or_B3_or_B4_B5_o  (\U_AHB/sel0_b16/or_B3_or_B4_B5_o_o , \U_AHB/sel0_b16/B3 , \U_AHB/sel0_b16/or_B4_B5_o );
  or \U_AHB/sel0_b16/or_B4_B5  (\U_AHB/sel0_b16/or_B4_B5_o , \U_AHB/sel0_b16/B4 , \U_AHB/sel0_b16/B5 );
  or \U_AHB/sel0_b16/or_B6_or_B7_B8_o  (\U_AHB/sel0_b16/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b16/B6 , \U_AHB/sel0_b16/or_B7_B8_o );
  or \U_AHB/sel0_b16/or_B7_B8  (\U_AHB/sel0_b16/or_B7_B8_o , \U_AHB/sel0_b16/B7 , \U_AHB/sel0_b16/B8 );
  or \U_AHB/sel0_b16/or_B9_or_B10_B11_o  (\U_AHB/sel0_b16/or_B9_or_B10_B11_o_o , \U_AHB/sel0_b16/B9 , \U_AHB/sel0_b16/or_B10_B11_o );
  or \U_AHB/sel0_b16/or_or_B0_or_B1_B2_o_  (\U_AHB/sel0_b16/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b16/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b16/or_B3_or_B4_B5_o_o );
  or \U_AHB/sel0_b16/or_or_B6_or_B7_B8_o_  (\U_AHB/sel0_b16/or_or_B6_or_B7_B8_o__o , \U_AHB/sel0_b16/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b16/or_B9_or_B10_B11_o_o );
  or \U_AHB/sel0_b16/or_or_or_B0_or_B1_B2  (\U_AHB/n114 [16], \U_AHB/sel0_b16/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b16/or_or_B6_or_B7_B8_o__o );
  and \U_AHB/sel0_b17/and_b0_0  (\U_AHB/sel0_b17/B0 , \U_AHB/h2h_hrdata [17], \U_AHB/n113 );
  and \U_AHB/sel0_b17/and_b0_1  (\U_AHB/sel0_b17/B1 , pnumcntA[17], \U_AHB/n111 );
  and \U_AHB/sel0_b17/and_b0_10  (\U_AHB/sel0_b17/B10 , pnumcnt1[17], \U_AHB/n84 );
  and \U_AHB/sel0_b17/and_b0_11  (\U_AHB/sel0_b17/B11 , pnumcnt0[17], \U_AHB/h2h_haddr [2]);
  and \U_AHB/sel0_b17/and_b0_2  (\U_AHB/sel0_b17/B2 , pnumcnt9[17], \U_AHB/n108 );
  and \U_AHB/sel0_b17/and_b0_3  (\U_AHB/sel0_b17/B3 , pnumcnt8[17], \U_AHB/n105 );
  and \U_AHB/sel0_b17/and_b0_4  (\U_AHB/sel0_b17/B4 , pnumcnt7[17], \U_AHB/n102 );
  and \U_AHB/sel0_b17/and_b0_5  (\U_AHB/sel0_b17/B5 , pnumcnt6[17], \U_AHB/n99 );
  and \U_AHB/sel0_b17/and_b0_6  (\U_AHB/sel0_b17/B6 , pnumcnt5[17], \U_AHB/n96 );
  and \U_AHB/sel0_b17/and_b0_7  (\U_AHB/sel0_b17/B7 , pnumcnt4[17], \U_AHB/n93 );
  and \U_AHB/sel0_b17/and_b0_8  (\U_AHB/sel0_b17/B8 , pnumcnt3[17], \U_AHB/n90 );
  and \U_AHB/sel0_b17/and_b0_9  (\U_AHB/sel0_b17/B9 , pnumcnt2[17], \U_AHB/n87 );
  or \U_AHB/sel0_b17/or_B0_or_B1_B2_o  (\U_AHB/sel0_b17/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b17/B0 , \U_AHB/sel0_b17/or_B1_B2_o );
  or \U_AHB/sel0_b17/or_B10_B11  (\U_AHB/sel0_b17/or_B10_B11_o , \U_AHB/sel0_b17/B10 , \U_AHB/sel0_b17/B11 );
  or \U_AHB/sel0_b17/or_B1_B2  (\U_AHB/sel0_b17/or_B1_B2_o , \U_AHB/sel0_b17/B1 , \U_AHB/sel0_b17/B2 );
  or \U_AHB/sel0_b17/or_B3_or_B4_B5_o  (\U_AHB/sel0_b17/or_B3_or_B4_B5_o_o , \U_AHB/sel0_b17/B3 , \U_AHB/sel0_b17/or_B4_B5_o );
  or \U_AHB/sel0_b17/or_B4_B5  (\U_AHB/sel0_b17/or_B4_B5_o , \U_AHB/sel0_b17/B4 , \U_AHB/sel0_b17/B5 );
  or \U_AHB/sel0_b17/or_B6_or_B7_B8_o  (\U_AHB/sel0_b17/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b17/B6 , \U_AHB/sel0_b17/or_B7_B8_o );
  or \U_AHB/sel0_b17/or_B7_B8  (\U_AHB/sel0_b17/or_B7_B8_o , \U_AHB/sel0_b17/B7 , \U_AHB/sel0_b17/B8 );
  or \U_AHB/sel0_b17/or_B9_or_B10_B11_o  (\U_AHB/sel0_b17/or_B9_or_B10_B11_o_o , \U_AHB/sel0_b17/B9 , \U_AHB/sel0_b17/or_B10_B11_o );
  or \U_AHB/sel0_b17/or_or_B0_or_B1_B2_o_  (\U_AHB/sel0_b17/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b17/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b17/or_B3_or_B4_B5_o_o );
  or \U_AHB/sel0_b17/or_or_B6_or_B7_B8_o_  (\U_AHB/sel0_b17/or_or_B6_or_B7_B8_o__o , \U_AHB/sel0_b17/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b17/or_B9_or_B10_B11_o_o );
  or \U_AHB/sel0_b17/or_or_or_B0_or_B1_B2  (\U_AHB/n114 [17], \U_AHB/sel0_b17/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b17/or_or_B6_or_B7_B8_o__o );
  and \U_AHB/sel0_b18/and_b0_0  (\U_AHB/sel0_b18/B0 , \U_AHB/h2h_hrdata [18], \U_AHB/n113 );
  and \U_AHB/sel0_b18/and_b0_1  (\U_AHB/sel0_b18/B1 , pnumcntA[18], \U_AHB/n111 );
  and \U_AHB/sel0_b18/and_b0_10  (\U_AHB/sel0_b18/B10 , pnumcnt1[18], \U_AHB/n84 );
  and \U_AHB/sel0_b18/and_b0_11  (\U_AHB/sel0_b18/B11 , pnumcnt0[18], \U_AHB/h2h_haddr [2]);
  and \U_AHB/sel0_b18/and_b0_2  (\U_AHB/sel0_b18/B2 , pnumcnt9[18], \U_AHB/n108 );
  and \U_AHB/sel0_b18/and_b0_3  (\U_AHB/sel0_b18/B3 , pnumcnt8[18], \U_AHB/n105 );
  and \U_AHB/sel0_b18/and_b0_4  (\U_AHB/sel0_b18/B4 , pnumcnt7[18], \U_AHB/n102 );
  and \U_AHB/sel0_b18/and_b0_5  (\U_AHB/sel0_b18/B5 , pnumcnt6[18], \U_AHB/n99 );
  and \U_AHB/sel0_b18/and_b0_6  (\U_AHB/sel0_b18/B6 , pnumcnt5[18], \U_AHB/n96 );
  and \U_AHB/sel0_b18/and_b0_7  (\U_AHB/sel0_b18/B7 , pnumcnt4[18], \U_AHB/n93 );
  and \U_AHB/sel0_b18/and_b0_8  (\U_AHB/sel0_b18/B8 , pnumcnt3[18], \U_AHB/n90 );
  and \U_AHB/sel0_b18/and_b0_9  (\U_AHB/sel0_b18/B9 , pnumcnt2[18], \U_AHB/n87 );
  or \U_AHB/sel0_b18/or_B0_or_B1_B2_o  (\U_AHB/sel0_b18/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b18/B0 , \U_AHB/sel0_b18/or_B1_B2_o );
  or \U_AHB/sel0_b18/or_B10_B11  (\U_AHB/sel0_b18/or_B10_B11_o , \U_AHB/sel0_b18/B10 , \U_AHB/sel0_b18/B11 );
  or \U_AHB/sel0_b18/or_B1_B2  (\U_AHB/sel0_b18/or_B1_B2_o , \U_AHB/sel0_b18/B1 , \U_AHB/sel0_b18/B2 );
  or \U_AHB/sel0_b18/or_B3_or_B4_B5_o  (\U_AHB/sel0_b18/or_B3_or_B4_B5_o_o , \U_AHB/sel0_b18/B3 , \U_AHB/sel0_b18/or_B4_B5_o );
  or \U_AHB/sel0_b18/or_B4_B5  (\U_AHB/sel0_b18/or_B4_B5_o , \U_AHB/sel0_b18/B4 , \U_AHB/sel0_b18/B5 );
  or \U_AHB/sel0_b18/or_B6_or_B7_B8_o  (\U_AHB/sel0_b18/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b18/B6 , \U_AHB/sel0_b18/or_B7_B8_o );
  or \U_AHB/sel0_b18/or_B7_B8  (\U_AHB/sel0_b18/or_B7_B8_o , \U_AHB/sel0_b18/B7 , \U_AHB/sel0_b18/B8 );
  or \U_AHB/sel0_b18/or_B9_or_B10_B11_o  (\U_AHB/sel0_b18/or_B9_or_B10_B11_o_o , \U_AHB/sel0_b18/B9 , \U_AHB/sel0_b18/or_B10_B11_o );
  or \U_AHB/sel0_b18/or_or_B0_or_B1_B2_o_  (\U_AHB/sel0_b18/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b18/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b18/or_B3_or_B4_B5_o_o );
  or \U_AHB/sel0_b18/or_or_B6_or_B7_B8_o_  (\U_AHB/sel0_b18/or_or_B6_or_B7_B8_o__o , \U_AHB/sel0_b18/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b18/or_B9_or_B10_B11_o_o );
  or \U_AHB/sel0_b18/or_or_or_B0_or_B1_B2  (\U_AHB/n114 [18], \U_AHB/sel0_b18/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b18/or_or_B6_or_B7_B8_o__o );
  and \U_AHB/sel0_b19/and_b0_0  (\U_AHB/sel0_b19/B0 , \U_AHB/h2h_hrdata [19], \U_AHB/n113 );
  and \U_AHB/sel0_b19/and_b0_1  (\U_AHB/sel0_b19/B1 , pnumcntA[19], \U_AHB/n111 );
  and \U_AHB/sel0_b19/and_b0_10  (\U_AHB/sel0_b19/B10 , pnumcnt1[19], \U_AHB/n84 );
  and \U_AHB/sel0_b19/and_b0_11  (\U_AHB/sel0_b19/B11 , pnumcnt0[19], \U_AHB/h2h_haddr [2]);
  and \U_AHB/sel0_b19/and_b0_2  (\U_AHB/sel0_b19/B2 , pnumcnt9[19], \U_AHB/n108 );
  and \U_AHB/sel0_b19/and_b0_3  (\U_AHB/sel0_b19/B3 , pnumcnt8[19], \U_AHB/n105 );
  and \U_AHB/sel0_b19/and_b0_4  (\U_AHB/sel0_b19/B4 , pnumcnt7[19], \U_AHB/n102 );
  and \U_AHB/sel0_b19/and_b0_5  (\U_AHB/sel0_b19/B5 , pnumcnt6[19], \U_AHB/n99 );
  and \U_AHB/sel0_b19/and_b0_6  (\U_AHB/sel0_b19/B6 , pnumcnt5[19], \U_AHB/n96 );
  and \U_AHB/sel0_b19/and_b0_7  (\U_AHB/sel0_b19/B7 , pnumcnt4[19], \U_AHB/n93 );
  and \U_AHB/sel0_b19/and_b0_8  (\U_AHB/sel0_b19/B8 , pnumcnt3[19], \U_AHB/n90 );
  and \U_AHB/sel0_b19/and_b0_9  (\U_AHB/sel0_b19/B9 , pnumcnt2[19], \U_AHB/n87 );
  or \U_AHB/sel0_b19/or_B0_or_B1_B2_o  (\U_AHB/sel0_b19/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b19/B0 , \U_AHB/sel0_b19/or_B1_B2_o );
  or \U_AHB/sel0_b19/or_B10_B11  (\U_AHB/sel0_b19/or_B10_B11_o , \U_AHB/sel0_b19/B10 , \U_AHB/sel0_b19/B11 );
  or \U_AHB/sel0_b19/or_B1_B2  (\U_AHB/sel0_b19/or_B1_B2_o , \U_AHB/sel0_b19/B1 , \U_AHB/sel0_b19/B2 );
  or \U_AHB/sel0_b19/or_B3_or_B4_B5_o  (\U_AHB/sel0_b19/or_B3_or_B4_B5_o_o , \U_AHB/sel0_b19/B3 , \U_AHB/sel0_b19/or_B4_B5_o );
  or \U_AHB/sel0_b19/or_B4_B5  (\U_AHB/sel0_b19/or_B4_B5_o , \U_AHB/sel0_b19/B4 , \U_AHB/sel0_b19/B5 );
  or \U_AHB/sel0_b19/or_B6_or_B7_B8_o  (\U_AHB/sel0_b19/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b19/B6 , \U_AHB/sel0_b19/or_B7_B8_o );
  or \U_AHB/sel0_b19/or_B7_B8  (\U_AHB/sel0_b19/or_B7_B8_o , \U_AHB/sel0_b19/B7 , \U_AHB/sel0_b19/B8 );
  or \U_AHB/sel0_b19/or_B9_or_B10_B11_o  (\U_AHB/sel0_b19/or_B9_or_B10_B11_o_o , \U_AHB/sel0_b19/B9 , \U_AHB/sel0_b19/or_B10_B11_o );
  or \U_AHB/sel0_b19/or_or_B0_or_B1_B2_o_  (\U_AHB/sel0_b19/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b19/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b19/or_B3_or_B4_B5_o_o );
  or \U_AHB/sel0_b19/or_or_B6_or_B7_B8_o_  (\U_AHB/sel0_b19/or_or_B6_or_B7_B8_o__o , \U_AHB/sel0_b19/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b19/or_B9_or_B10_B11_o_o );
  or \U_AHB/sel0_b19/or_or_or_B0_or_B1_B2  (\U_AHB/n114 [19], \U_AHB/sel0_b19/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b19/or_or_B6_or_B7_B8_o__o );
  and \U_AHB/sel0_b2/and_b0_0  (\U_AHB/sel0_b2/B0 , \U_AHB/h2h_hrdata [2], \U_AHB/n113 );
  and \U_AHB/sel0_b2/and_b0_1  (\U_AHB/sel0_b2/B1 , pnumcntA[2], \U_AHB/n111 );
  and \U_AHB/sel0_b2/and_b0_10  (\U_AHB/sel0_b2/B10 , pnumcnt1[2], \U_AHB/n84 );
  and \U_AHB/sel0_b2/and_b0_11  (\U_AHB/sel0_b2/B11 , pnumcnt0[2], \U_AHB/h2h_haddr [2]);
  and \U_AHB/sel0_b2/and_b0_2  (\U_AHB/sel0_b2/B2 , pnumcnt9[2], \U_AHB/n108 );
  and \U_AHB/sel0_b2/and_b0_3  (\U_AHB/sel0_b2/B3 , pnumcnt8[2], \U_AHB/n105 );
  and \U_AHB/sel0_b2/and_b0_4  (\U_AHB/sel0_b2/B4 , pnumcnt7[2], \U_AHB/n102 );
  and \U_AHB/sel0_b2/and_b0_5  (\U_AHB/sel0_b2/B5 , pnumcnt6[2], \U_AHB/n99 );
  and \U_AHB/sel0_b2/and_b0_6  (\U_AHB/sel0_b2/B6 , pnumcnt5[2], \U_AHB/n96 );
  and \U_AHB/sel0_b2/and_b0_7  (\U_AHB/sel0_b2/B7 , pnumcnt4[2], \U_AHB/n93 );
  and \U_AHB/sel0_b2/and_b0_8  (\U_AHB/sel0_b2/B8 , pnumcnt3[2], \U_AHB/n90 );
  and \U_AHB/sel0_b2/and_b0_9  (\U_AHB/sel0_b2/B9 , pnumcnt2[2], \U_AHB/n87 );
  or \U_AHB/sel0_b2/or_B0_or_B1_B2_o  (\U_AHB/sel0_b2/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b2/B0 , \U_AHB/sel0_b2/or_B1_B2_o );
  or \U_AHB/sel0_b2/or_B10_B11  (\U_AHB/sel0_b2/or_B10_B11_o , \U_AHB/sel0_b2/B10 , \U_AHB/sel0_b2/B11 );
  or \U_AHB/sel0_b2/or_B1_B2  (\U_AHB/sel0_b2/or_B1_B2_o , \U_AHB/sel0_b2/B1 , \U_AHB/sel0_b2/B2 );
  or \U_AHB/sel0_b2/or_B3_or_B4_B5_o  (\U_AHB/sel0_b2/or_B3_or_B4_B5_o_o , \U_AHB/sel0_b2/B3 , \U_AHB/sel0_b2/or_B4_B5_o );
  or \U_AHB/sel0_b2/or_B4_B5  (\U_AHB/sel0_b2/or_B4_B5_o , \U_AHB/sel0_b2/B4 , \U_AHB/sel0_b2/B5 );
  or \U_AHB/sel0_b2/or_B6_or_B7_B8_o  (\U_AHB/sel0_b2/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b2/B6 , \U_AHB/sel0_b2/or_B7_B8_o );
  or \U_AHB/sel0_b2/or_B7_B8  (\U_AHB/sel0_b2/or_B7_B8_o , \U_AHB/sel0_b2/B7 , \U_AHB/sel0_b2/B8 );
  or \U_AHB/sel0_b2/or_B9_or_B10_B11_o  (\U_AHB/sel0_b2/or_B9_or_B10_B11_o_o , \U_AHB/sel0_b2/B9 , \U_AHB/sel0_b2/or_B10_B11_o );
  or \U_AHB/sel0_b2/or_or_B0_or_B1_B2_o_  (\U_AHB/sel0_b2/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b2/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b2/or_B3_or_B4_B5_o_o );
  or \U_AHB/sel0_b2/or_or_B6_or_B7_B8_o_  (\U_AHB/sel0_b2/or_or_B6_or_B7_B8_o__o , \U_AHB/sel0_b2/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b2/or_B9_or_B10_B11_o_o );
  or \U_AHB/sel0_b2/or_or_or_B0_or_B1_B2  (\U_AHB/n114 [2], \U_AHB/sel0_b2/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b2/or_or_B6_or_B7_B8_o__o );
  and \U_AHB/sel0_b20/and_b0_0  (\U_AHB/sel0_b20/B0 , \U_AHB/h2h_hrdata [20], \U_AHB/n113 );
  and \U_AHB/sel0_b20/and_b0_1  (\U_AHB/sel0_b20/B1 , pnumcntA[20], \U_AHB/n111 );
  and \U_AHB/sel0_b20/and_b0_10  (\U_AHB/sel0_b20/B10 , pnumcnt1[20], \U_AHB/n84 );
  and \U_AHB/sel0_b20/and_b0_11  (\U_AHB/sel0_b20/B11 , pnumcnt0[20], \U_AHB/h2h_haddr [2]);
  and \U_AHB/sel0_b20/and_b0_2  (\U_AHB/sel0_b20/B2 , pnumcnt9[20], \U_AHB/n108 );
  and \U_AHB/sel0_b20/and_b0_3  (\U_AHB/sel0_b20/B3 , pnumcnt8[20], \U_AHB/n105 );
  and \U_AHB/sel0_b20/and_b0_4  (\U_AHB/sel0_b20/B4 , pnumcnt7[20], \U_AHB/n102 );
  and \U_AHB/sel0_b20/and_b0_5  (\U_AHB/sel0_b20/B5 , pnumcnt6[20], \U_AHB/n99 );
  and \U_AHB/sel0_b20/and_b0_6  (\U_AHB/sel0_b20/B6 , pnumcnt5[20], \U_AHB/n96 );
  and \U_AHB/sel0_b20/and_b0_7  (\U_AHB/sel0_b20/B7 , pnumcnt4[20], \U_AHB/n93 );
  and \U_AHB/sel0_b20/and_b0_8  (\U_AHB/sel0_b20/B8 , pnumcnt3[20], \U_AHB/n90 );
  and \U_AHB/sel0_b20/and_b0_9  (\U_AHB/sel0_b20/B9 , pnumcnt2[20], \U_AHB/n87 );
  or \U_AHB/sel0_b20/or_B0_or_B1_B2_o  (\U_AHB/sel0_b20/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b20/B0 , \U_AHB/sel0_b20/or_B1_B2_o );
  or \U_AHB/sel0_b20/or_B10_B11  (\U_AHB/sel0_b20/or_B10_B11_o , \U_AHB/sel0_b20/B10 , \U_AHB/sel0_b20/B11 );
  or \U_AHB/sel0_b20/or_B1_B2  (\U_AHB/sel0_b20/or_B1_B2_o , \U_AHB/sel0_b20/B1 , \U_AHB/sel0_b20/B2 );
  or \U_AHB/sel0_b20/or_B3_or_B4_B5_o  (\U_AHB/sel0_b20/or_B3_or_B4_B5_o_o , \U_AHB/sel0_b20/B3 , \U_AHB/sel0_b20/or_B4_B5_o );
  or \U_AHB/sel0_b20/or_B4_B5  (\U_AHB/sel0_b20/or_B4_B5_o , \U_AHB/sel0_b20/B4 , \U_AHB/sel0_b20/B5 );
  or \U_AHB/sel0_b20/or_B6_or_B7_B8_o  (\U_AHB/sel0_b20/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b20/B6 , \U_AHB/sel0_b20/or_B7_B8_o );
  or \U_AHB/sel0_b20/or_B7_B8  (\U_AHB/sel0_b20/or_B7_B8_o , \U_AHB/sel0_b20/B7 , \U_AHB/sel0_b20/B8 );
  or \U_AHB/sel0_b20/or_B9_or_B10_B11_o  (\U_AHB/sel0_b20/or_B9_or_B10_B11_o_o , \U_AHB/sel0_b20/B9 , \U_AHB/sel0_b20/or_B10_B11_o );
  or \U_AHB/sel0_b20/or_or_B0_or_B1_B2_o_  (\U_AHB/sel0_b20/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b20/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b20/or_B3_or_B4_B5_o_o );
  or \U_AHB/sel0_b20/or_or_B6_or_B7_B8_o_  (\U_AHB/sel0_b20/or_or_B6_or_B7_B8_o__o , \U_AHB/sel0_b20/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b20/or_B9_or_B10_B11_o_o );
  or \U_AHB/sel0_b20/or_or_or_B0_or_B1_B2  (\U_AHB/n114 [20], \U_AHB/sel0_b20/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b20/or_or_B6_or_B7_B8_o__o );
  and \U_AHB/sel0_b21/and_b0_0  (\U_AHB/sel0_b21/B0 , \U_AHB/h2h_hrdata [21], \U_AHB/n113 );
  and \U_AHB/sel0_b21/and_b0_1  (\U_AHB/sel0_b21/B1 , pnumcntA[21], \U_AHB/n111 );
  and \U_AHB/sel0_b21/and_b0_10  (\U_AHB/sel0_b21/B10 , pnumcnt1[21], \U_AHB/n84 );
  and \U_AHB/sel0_b21/and_b0_11  (\U_AHB/sel0_b21/B11 , pnumcnt0[21], \U_AHB/h2h_haddr [2]);
  and \U_AHB/sel0_b21/and_b0_2  (\U_AHB/sel0_b21/B2 , pnumcnt9[21], \U_AHB/n108 );
  and \U_AHB/sel0_b21/and_b0_3  (\U_AHB/sel0_b21/B3 , pnumcnt8[21], \U_AHB/n105 );
  and \U_AHB/sel0_b21/and_b0_4  (\U_AHB/sel0_b21/B4 , pnumcnt7[21], \U_AHB/n102 );
  and \U_AHB/sel0_b21/and_b0_5  (\U_AHB/sel0_b21/B5 , pnumcnt6[21], \U_AHB/n99 );
  and \U_AHB/sel0_b21/and_b0_6  (\U_AHB/sel0_b21/B6 , pnumcnt5[21], \U_AHB/n96 );
  and \U_AHB/sel0_b21/and_b0_7  (\U_AHB/sel0_b21/B7 , pnumcnt4[21], \U_AHB/n93 );
  and \U_AHB/sel0_b21/and_b0_8  (\U_AHB/sel0_b21/B8 , pnumcnt3[21], \U_AHB/n90 );
  and \U_AHB/sel0_b21/and_b0_9  (\U_AHB/sel0_b21/B9 , pnumcnt2[21], \U_AHB/n87 );
  or \U_AHB/sel0_b21/or_B0_or_B1_B2_o  (\U_AHB/sel0_b21/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b21/B0 , \U_AHB/sel0_b21/or_B1_B2_o );
  or \U_AHB/sel0_b21/or_B10_B11  (\U_AHB/sel0_b21/or_B10_B11_o , \U_AHB/sel0_b21/B10 , \U_AHB/sel0_b21/B11 );
  or \U_AHB/sel0_b21/or_B1_B2  (\U_AHB/sel0_b21/or_B1_B2_o , \U_AHB/sel0_b21/B1 , \U_AHB/sel0_b21/B2 );
  or \U_AHB/sel0_b21/or_B3_or_B4_B5_o  (\U_AHB/sel0_b21/or_B3_or_B4_B5_o_o , \U_AHB/sel0_b21/B3 , \U_AHB/sel0_b21/or_B4_B5_o );
  or \U_AHB/sel0_b21/or_B4_B5  (\U_AHB/sel0_b21/or_B4_B5_o , \U_AHB/sel0_b21/B4 , \U_AHB/sel0_b21/B5 );
  or \U_AHB/sel0_b21/or_B6_or_B7_B8_o  (\U_AHB/sel0_b21/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b21/B6 , \U_AHB/sel0_b21/or_B7_B8_o );
  or \U_AHB/sel0_b21/or_B7_B8  (\U_AHB/sel0_b21/or_B7_B8_o , \U_AHB/sel0_b21/B7 , \U_AHB/sel0_b21/B8 );
  or \U_AHB/sel0_b21/or_B9_or_B10_B11_o  (\U_AHB/sel0_b21/or_B9_or_B10_B11_o_o , \U_AHB/sel0_b21/B9 , \U_AHB/sel0_b21/or_B10_B11_o );
  or \U_AHB/sel0_b21/or_or_B0_or_B1_B2_o_  (\U_AHB/sel0_b21/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b21/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b21/or_B3_or_B4_B5_o_o );
  or \U_AHB/sel0_b21/or_or_B6_or_B7_B8_o_  (\U_AHB/sel0_b21/or_or_B6_or_B7_B8_o__o , \U_AHB/sel0_b21/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b21/or_B9_or_B10_B11_o_o );
  or \U_AHB/sel0_b21/or_or_or_B0_or_B1_B2  (\U_AHB/n114 [21], \U_AHB/sel0_b21/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b21/or_or_B6_or_B7_B8_o__o );
  and \U_AHB/sel0_b22/and_b0_0  (\U_AHB/sel0_b22/B0 , \U_AHB/h2h_hrdata [22], \U_AHB/n113 );
  and \U_AHB/sel0_b22/and_b0_1  (\U_AHB/sel0_b22/B1 , pnumcntA[22], \U_AHB/n111 );
  and \U_AHB/sel0_b22/and_b0_10  (\U_AHB/sel0_b22/B10 , pnumcnt1[22], \U_AHB/n84 );
  and \U_AHB/sel0_b22/and_b0_11  (\U_AHB/sel0_b22/B11 , pnumcnt0[22], \U_AHB/h2h_haddr [2]);
  and \U_AHB/sel0_b22/and_b0_2  (\U_AHB/sel0_b22/B2 , pnumcnt9[22], \U_AHB/n108 );
  and \U_AHB/sel0_b22/and_b0_3  (\U_AHB/sel0_b22/B3 , pnumcnt8[22], \U_AHB/n105 );
  and \U_AHB/sel0_b22/and_b0_4  (\U_AHB/sel0_b22/B4 , pnumcnt7[22], \U_AHB/n102 );
  and \U_AHB/sel0_b22/and_b0_5  (\U_AHB/sel0_b22/B5 , pnumcnt6[22], \U_AHB/n99 );
  and \U_AHB/sel0_b22/and_b0_6  (\U_AHB/sel0_b22/B6 , pnumcnt5[22], \U_AHB/n96 );
  and \U_AHB/sel0_b22/and_b0_7  (\U_AHB/sel0_b22/B7 , pnumcnt4[22], \U_AHB/n93 );
  and \U_AHB/sel0_b22/and_b0_8  (\U_AHB/sel0_b22/B8 , pnumcnt3[22], \U_AHB/n90 );
  and \U_AHB/sel0_b22/and_b0_9  (\U_AHB/sel0_b22/B9 , pnumcnt2[22], \U_AHB/n87 );
  or \U_AHB/sel0_b22/or_B0_or_B1_B2_o  (\U_AHB/sel0_b22/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b22/B0 , \U_AHB/sel0_b22/or_B1_B2_o );
  or \U_AHB/sel0_b22/or_B10_B11  (\U_AHB/sel0_b22/or_B10_B11_o , \U_AHB/sel0_b22/B10 , \U_AHB/sel0_b22/B11 );
  or \U_AHB/sel0_b22/or_B1_B2  (\U_AHB/sel0_b22/or_B1_B2_o , \U_AHB/sel0_b22/B1 , \U_AHB/sel0_b22/B2 );
  or \U_AHB/sel0_b22/or_B3_or_B4_B5_o  (\U_AHB/sel0_b22/or_B3_or_B4_B5_o_o , \U_AHB/sel0_b22/B3 , \U_AHB/sel0_b22/or_B4_B5_o );
  or \U_AHB/sel0_b22/or_B4_B5  (\U_AHB/sel0_b22/or_B4_B5_o , \U_AHB/sel0_b22/B4 , \U_AHB/sel0_b22/B5 );
  or \U_AHB/sel0_b22/or_B6_or_B7_B8_o  (\U_AHB/sel0_b22/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b22/B6 , \U_AHB/sel0_b22/or_B7_B8_o );
  or \U_AHB/sel0_b22/or_B7_B8  (\U_AHB/sel0_b22/or_B7_B8_o , \U_AHB/sel0_b22/B7 , \U_AHB/sel0_b22/B8 );
  or \U_AHB/sel0_b22/or_B9_or_B10_B11_o  (\U_AHB/sel0_b22/or_B9_or_B10_B11_o_o , \U_AHB/sel0_b22/B9 , \U_AHB/sel0_b22/or_B10_B11_o );
  or \U_AHB/sel0_b22/or_or_B0_or_B1_B2_o_  (\U_AHB/sel0_b22/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b22/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b22/or_B3_or_B4_B5_o_o );
  or \U_AHB/sel0_b22/or_or_B6_or_B7_B8_o_  (\U_AHB/sel0_b22/or_or_B6_or_B7_B8_o__o , \U_AHB/sel0_b22/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b22/or_B9_or_B10_B11_o_o );
  or \U_AHB/sel0_b22/or_or_or_B0_or_B1_B2  (\U_AHB/n114 [22], \U_AHB/sel0_b22/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b22/or_or_B6_or_B7_B8_o__o );
  and \U_AHB/sel0_b23/and_b0_0  (\U_AHB/sel0_b23/B0 , \U_AHB/h2h_hrdata [23], \U_AHB/n113 );
  and \U_AHB/sel0_b23/and_b0_1  (\U_AHB/sel0_b23/B1 , pnumcntA[23], \U_AHB/n111 );
  and \U_AHB/sel0_b23/and_b0_10  (\U_AHB/sel0_b23/B10 , pnumcnt1[23], \U_AHB/n84 );
  and \U_AHB/sel0_b23/and_b0_11  (\U_AHB/sel0_b23/B11 , pnumcnt0[23], \U_AHB/h2h_haddr [2]);
  and \U_AHB/sel0_b23/and_b0_2  (\U_AHB/sel0_b23/B2 , pnumcnt9[23], \U_AHB/n108 );
  and \U_AHB/sel0_b23/and_b0_3  (\U_AHB/sel0_b23/B3 , pnumcnt8[23], \U_AHB/n105 );
  and \U_AHB/sel0_b23/and_b0_4  (\U_AHB/sel0_b23/B4 , pnumcnt7[23], \U_AHB/n102 );
  and \U_AHB/sel0_b23/and_b0_5  (\U_AHB/sel0_b23/B5 , pnumcnt6[23], \U_AHB/n99 );
  and \U_AHB/sel0_b23/and_b0_6  (\U_AHB/sel0_b23/B6 , pnumcnt5[23], \U_AHB/n96 );
  and \U_AHB/sel0_b23/and_b0_7  (\U_AHB/sel0_b23/B7 , pnumcnt4[23], \U_AHB/n93 );
  and \U_AHB/sel0_b23/and_b0_8  (\U_AHB/sel0_b23/B8 , pnumcnt3[23], \U_AHB/n90 );
  and \U_AHB/sel0_b23/and_b0_9  (\U_AHB/sel0_b23/B9 , pnumcnt2[23], \U_AHB/n87 );
  or \U_AHB/sel0_b23/or_B0_or_B1_B2_o  (\U_AHB/sel0_b23/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b23/B0 , \U_AHB/sel0_b23/or_B1_B2_o );
  or \U_AHB/sel0_b23/or_B10_B11  (\U_AHB/sel0_b23/or_B10_B11_o , \U_AHB/sel0_b23/B10 , \U_AHB/sel0_b23/B11 );
  or \U_AHB/sel0_b23/or_B1_B2  (\U_AHB/sel0_b23/or_B1_B2_o , \U_AHB/sel0_b23/B1 , \U_AHB/sel0_b23/B2 );
  or \U_AHB/sel0_b23/or_B3_or_B4_B5_o  (\U_AHB/sel0_b23/or_B3_or_B4_B5_o_o , \U_AHB/sel0_b23/B3 , \U_AHB/sel0_b23/or_B4_B5_o );
  or \U_AHB/sel0_b23/or_B4_B5  (\U_AHB/sel0_b23/or_B4_B5_o , \U_AHB/sel0_b23/B4 , \U_AHB/sel0_b23/B5 );
  or \U_AHB/sel0_b23/or_B6_or_B7_B8_o  (\U_AHB/sel0_b23/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b23/B6 , \U_AHB/sel0_b23/or_B7_B8_o );
  or \U_AHB/sel0_b23/or_B7_B8  (\U_AHB/sel0_b23/or_B7_B8_o , \U_AHB/sel0_b23/B7 , \U_AHB/sel0_b23/B8 );
  or \U_AHB/sel0_b23/or_B9_or_B10_B11_o  (\U_AHB/sel0_b23/or_B9_or_B10_B11_o_o , \U_AHB/sel0_b23/B9 , \U_AHB/sel0_b23/or_B10_B11_o );
  or \U_AHB/sel0_b23/or_or_B0_or_B1_B2_o_  (\U_AHB/sel0_b23/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b23/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b23/or_B3_or_B4_B5_o_o );
  or \U_AHB/sel0_b23/or_or_B6_or_B7_B8_o_  (\U_AHB/sel0_b23/or_or_B6_or_B7_B8_o__o , \U_AHB/sel0_b23/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b23/or_B9_or_B10_B11_o_o );
  or \U_AHB/sel0_b23/or_or_or_B0_or_B1_B2  (\U_AHB/n114 [23], \U_AHB/sel0_b23/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b23/or_or_B6_or_B7_B8_o__o );
  AL_MUX \U_AHB/sel0_b24  (
    .i0(1'b0),
    .i1(\U_AHB/h2h_hrdata [24]),
    .sel(\U_AHB/n113 ),
    .o(\U_AHB/n114 [24]));  // src/AHB.v(101)
  AL_MUX \U_AHB/sel0_b25  (
    .i0(1'b0),
    .i1(\U_AHB/h2h_hrdata [25]),
    .sel(\U_AHB/n113 ),
    .o(\U_AHB/n114 [25]));  // src/AHB.v(101)
  AL_MUX \U_AHB/sel0_b26  (
    .i0(1'b0),
    .i1(\U_AHB/h2h_hrdata [26]),
    .sel(\U_AHB/n113 ),
    .o(\U_AHB/n114 [26]));  // src/AHB.v(101)
  AL_MUX \U_AHB/sel0_b27  (
    .i0(1'b0),
    .i1(\U_AHB/h2h_hrdata [27]),
    .sel(\U_AHB/n113 ),
    .o(\U_AHB/n114 [27]));  // src/AHB.v(101)
  AL_MUX \U_AHB/sel0_b28  (
    .i0(1'b0),
    .i1(\U_AHB/h2h_hrdata [28]),
    .sel(\U_AHB/n113 ),
    .o(\U_AHB/n114 [28]));  // src/AHB.v(101)
  AL_MUX \U_AHB/sel0_b29  (
    .i0(1'b0),
    .i1(\U_AHB/h2h_hrdata [29]),
    .sel(\U_AHB/n113 ),
    .o(\U_AHB/n114 [29]));  // src/AHB.v(101)
  and \U_AHB/sel0_b3/and_b0_0  (\U_AHB/sel0_b3/B0 , \U_AHB/h2h_hrdata [3], \U_AHB/n113 );
  and \U_AHB/sel0_b3/and_b0_1  (\U_AHB/sel0_b3/B1 , pnumcntA[3], \U_AHB/n111 );
  and \U_AHB/sel0_b3/and_b0_10  (\U_AHB/sel0_b3/B10 , pnumcnt1[3], \U_AHB/n84 );
  and \U_AHB/sel0_b3/and_b0_11  (\U_AHB/sel0_b3/B11 , pnumcnt0[3], \U_AHB/h2h_haddr [2]);
  and \U_AHB/sel0_b3/and_b0_2  (\U_AHB/sel0_b3/B2 , pnumcnt9[3], \U_AHB/n108 );
  and \U_AHB/sel0_b3/and_b0_3  (\U_AHB/sel0_b3/B3 , pnumcnt8[3], \U_AHB/n105 );
  and \U_AHB/sel0_b3/and_b0_4  (\U_AHB/sel0_b3/B4 , pnumcnt7[3], \U_AHB/n102 );
  and \U_AHB/sel0_b3/and_b0_5  (\U_AHB/sel0_b3/B5 , pnumcnt6[3], \U_AHB/n99 );
  and \U_AHB/sel0_b3/and_b0_6  (\U_AHB/sel0_b3/B6 , pnumcnt5[3], \U_AHB/n96 );
  and \U_AHB/sel0_b3/and_b0_7  (\U_AHB/sel0_b3/B7 , pnumcnt4[3], \U_AHB/n93 );
  and \U_AHB/sel0_b3/and_b0_8  (\U_AHB/sel0_b3/B8 , pnumcnt3[3], \U_AHB/n90 );
  and \U_AHB/sel0_b3/and_b0_9  (\U_AHB/sel0_b3/B9 , pnumcnt2[3], \U_AHB/n87 );
  or \U_AHB/sel0_b3/or_B0_or_B1_B2_o  (\U_AHB/sel0_b3/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b3/B0 , \U_AHB/sel0_b3/or_B1_B2_o );
  or \U_AHB/sel0_b3/or_B10_B11  (\U_AHB/sel0_b3/or_B10_B11_o , \U_AHB/sel0_b3/B10 , \U_AHB/sel0_b3/B11 );
  or \U_AHB/sel0_b3/or_B1_B2  (\U_AHB/sel0_b3/or_B1_B2_o , \U_AHB/sel0_b3/B1 , \U_AHB/sel0_b3/B2 );
  or \U_AHB/sel0_b3/or_B3_or_B4_B5_o  (\U_AHB/sel0_b3/or_B3_or_B4_B5_o_o , \U_AHB/sel0_b3/B3 , \U_AHB/sel0_b3/or_B4_B5_o );
  or \U_AHB/sel0_b3/or_B4_B5  (\U_AHB/sel0_b3/or_B4_B5_o , \U_AHB/sel0_b3/B4 , \U_AHB/sel0_b3/B5 );
  or \U_AHB/sel0_b3/or_B6_or_B7_B8_o  (\U_AHB/sel0_b3/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b3/B6 , \U_AHB/sel0_b3/or_B7_B8_o );
  or \U_AHB/sel0_b3/or_B7_B8  (\U_AHB/sel0_b3/or_B7_B8_o , \U_AHB/sel0_b3/B7 , \U_AHB/sel0_b3/B8 );
  or \U_AHB/sel0_b3/or_B9_or_B10_B11_o  (\U_AHB/sel0_b3/or_B9_or_B10_B11_o_o , \U_AHB/sel0_b3/B9 , \U_AHB/sel0_b3/or_B10_B11_o );
  or \U_AHB/sel0_b3/or_or_B0_or_B1_B2_o_  (\U_AHB/sel0_b3/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b3/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b3/or_B3_or_B4_B5_o_o );
  or \U_AHB/sel0_b3/or_or_B6_or_B7_B8_o_  (\U_AHB/sel0_b3/or_or_B6_or_B7_B8_o__o , \U_AHB/sel0_b3/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b3/or_B9_or_B10_B11_o_o );
  or \U_AHB/sel0_b3/or_or_or_B0_or_B1_B2  (\U_AHB/n114 [3], \U_AHB/sel0_b3/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b3/or_or_B6_or_B7_B8_o__o );
  AL_MUX \U_AHB/sel0_b30  (
    .i0(1'b0),
    .i1(\U_AHB/h2h_hrdata [30]),
    .sel(\U_AHB/n113 ),
    .o(\U_AHB/n114 [30]));  // src/AHB.v(101)
  AL_MUX \U_AHB/sel0_b31  (
    .i0(1'b0),
    .i1(\U_AHB/h2h_hrdata [31]),
    .sel(\U_AHB/n113 ),
    .o(\U_AHB/n114 [31]));  // src/AHB.v(101)
  and \U_AHB/sel0_b4/and_b0_0  (\U_AHB/sel0_b4/B0 , \U_AHB/h2h_hrdata [4], \U_AHB/n113 );
  and \U_AHB/sel0_b4/and_b0_1  (\U_AHB/sel0_b4/B1 , pnumcntA[4], \U_AHB/n111 );
  and \U_AHB/sel0_b4/and_b0_10  (\U_AHB/sel0_b4/B10 , pnumcnt1[4], \U_AHB/n84 );
  and \U_AHB/sel0_b4/and_b0_11  (\U_AHB/sel0_b4/B11 , pnumcnt0[4], \U_AHB/h2h_haddr [2]);
  and \U_AHB/sel0_b4/and_b0_2  (\U_AHB/sel0_b4/B2 , pnumcnt9[4], \U_AHB/n108 );
  and \U_AHB/sel0_b4/and_b0_3  (\U_AHB/sel0_b4/B3 , pnumcnt8[4], \U_AHB/n105 );
  and \U_AHB/sel0_b4/and_b0_4  (\U_AHB/sel0_b4/B4 , pnumcnt7[4], \U_AHB/n102 );
  and \U_AHB/sel0_b4/and_b0_5  (\U_AHB/sel0_b4/B5 , pnumcnt6[4], \U_AHB/n99 );
  and \U_AHB/sel0_b4/and_b0_6  (\U_AHB/sel0_b4/B6 , pnumcnt5[4], \U_AHB/n96 );
  and \U_AHB/sel0_b4/and_b0_7  (\U_AHB/sel0_b4/B7 , pnumcnt4[4], \U_AHB/n93 );
  and \U_AHB/sel0_b4/and_b0_8  (\U_AHB/sel0_b4/B8 , pnumcnt3[4], \U_AHB/n90 );
  and \U_AHB/sel0_b4/and_b0_9  (\U_AHB/sel0_b4/B9 , pnumcnt2[4], \U_AHB/n87 );
  or \U_AHB/sel0_b4/or_B0_or_B1_B2_o  (\U_AHB/sel0_b4/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b4/B0 , \U_AHB/sel0_b4/or_B1_B2_o );
  or \U_AHB/sel0_b4/or_B10_B11  (\U_AHB/sel0_b4/or_B10_B11_o , \U_AHB/sel0_b4/B10 , \U_AHB/sel0_b4/B11 );
  or \U_AHB/sel0_b4/or_B1_B2  (\U_AHB/sel0_b4/or_B1_B2_o , \U_AHB/sel0_b4/B1 , \U_AHB/sel0_b4/B2 );
  or \U_AHB/sel0_b4/or_B3_or_B4_B5_o  (\U_AHB/sel0_b4/or_B3_or_B4_B5_o_o , \U_AHB/sel0_b4/B3 , \U_AHB/sel0_b4/or_B4_B5_o );
  or \U_AHB/sel0_b4/or_B4_B5  (\U_AHB/sel0_b4/or_B4_B5_o , \U_AHB/sel0_b4/B4 , \U_AHB/sel0_b4/B5 );
  or \U_AHB/sel0_b4/or_B6_or_B7_B8_o  (\U_AHB/sel0_b4/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b4/B6 , \U_AHB/sel0_b4/or_B7_B8_o );
  or \U_AHB/sel0_b4/or_B7_B8  (\U_AHB/sel0_b4/or_B7_B8_o , \U_AHB/sel0_b4/B7 , \U_AHB/sel0_b4/B8 );
  or \U_AHB/sel0_b4/or_B9_or_B10_B11_o  (\U_AHB/sel0_b4/or_B9_or_B10_B11_o_o , \U_AHB/sel0_b4/B9 , \U_AHB/sel0_b4/or_B10_B11_o );
  or \U_AHB/sel0_b4/or_or_B0_or_B1_B2_o_  (\U_AHB/sel0_b4/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b4/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b4/or_B3_or_B4_B5_o_o );
  or \U_AHB/sel0_b4/or_or_B6_or_B7_B8_o_  (\U_AHB/sel0_b4/or_or_B6_or_B7_B8_o__o , \U_AHB/sel0_b4/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b4/or_B9_or_B10_B11_o_o );
  or \U_AHB/sel0_b4/or_or_or_B0_or_B1_B2  (\U_AHB/n114 [4], \U_AHB/sel0_b4/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b4/or_or_B6_or_B7_B8_o__o );
  and \U_AHB/sel0_b5/and_b0_0  (\U_AHB/sel0_b5/B0 , \U_AHB/h2h_hrdata [5], \U_AHB/n113 );
  and \U_AHB/sel0_b5/and_b0_1  (\U_AHB/sel0_b5/B1 , pnumcntA[5], \U_AHB/n111 );
  and \U_AHB/sel0_b5/and_b0_10  (\U_AHB/sel0_b5/B10 , pnumcnt1[5], \U_AHB/n84 );
  and \U_AHB/sel0_b5/and_b0_11  (\U_AHB/sel0_b5/B11 , pnumcnt0[5], \U_AHB/h2h_haddr [2]);
  and \U_AHB/sel0_b5/and_b0_2  (\U_AHB/sel0_b5/B2 , pnumcnt9[5], \U_AHB/n108 );
  and \U_AHB/sel0_b5/and_b0_3  (\U_AHB/sel0_b5/B3 , pnumcnt8[5], \U_AHB/n105 );
  and \U_AHB/sel0_b5/and_b0_4  (\U_AHB/sel0_b5/B4 , pnumcnt7[5], \U_AHB/n102 );
  and \U_AHB/sel0_b5/and_b0_5  (\U_AHB/sel0_b5/B5 , pnumcnt6[5], \U_AHB/n99 );
  and \U_AHB/sel0_b5/and_b0_6  (\U_AHB/sel0_b5/B6 , pnumcnt5[5], \U_AHB/n96 );
  and \U_AHB/sel0_b5/and_b0_7  (\U_AHB/sel0_b5/B7 , pnumcnt4[5], \U_AHB/n93 );
  and \U_AHB/sel0_b5/and_b0_8  (\U_AHB/sel0_b5/B8 , pnumcnt3[5], \U_AHB/n90 );
  and \U_AHB/sel0_b5/and_b0_9  (\U_AHB/sel0_b5/B9 , pnumcnt2[5], \U_AHB/n87 );
  or \U_AHB/sel0_b5/or_B0_or_B1_B2_o  (\U_AHB/sel0_b5/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b5/B0 , \U_AHB/sel0_b5/or_B1_B2_o );
  or \U_AHB/sel0_b5/or_B10_B11  (\U_AHB/sel0_b5/or_B10_B11_o , \U_AHB/sel0_b5/B10 , \U_AHB/sel0_b5/B11 );
  or \U_AHB/sel0_b5/or_B1_B2  (\U_AHB/sel0_b5/or_B1_B2_o , \U_AHB/sel0_b5/B1 , \U_AHB/sel0_b5/B2 );
  or \U_AHB/sel0_b5/or_B3_or_B4_B5_o  (\U_AHB/sel0_b5/or_B3_or_B4_B5_o_o , \U_AHB/sel0_b5/B3 , \U_AHB/sel0_b5/or_B4_B5_o );
  or \U_AHB/sel0_b5/or_B4_B5  (\U_AHB/sel0_b5/or_B4_B5_o , \U_AHB/sel0_b5/B4 , \U_AHB/sel0_b5/B5 );
  or \U_AHB/sel0_b5/or_B6_or_B7_B8_o  (\U_AHB/sel0_b5/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b5/B6 , \U_AHB/sel0_b5/or_B7_B8_o );
  or \U_AHB/sel0_b5/or_B7_B8  (\U_AHB/sel0_b5/or_B7_B8_o , \U_AHB/sel0_b5/B7 , \U_AHB/sel0_b5/B8 );
  or \U_AHB/sel0_b5/or_B9_or_B10_B11_o  (\U_AHB/sel0_b5/or_B9_or_B10_B11_o_o , \U_AHB/sel0_b5/B9 , \U_AHB/sel0_b5/or_B10_B11_o );
  or \U_AHB/sel0_b5/or_or_B0_or_B1_B2_o_  (\U_AHB/sel0_b5/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b5/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b5/or_B3_or_B4_B5_o_o );
  or \U_AHB/sel0_b5/or_or_B6_or_B7_B8_o_  (\U_AHB/sel0_b5/or_or_B6_or_B7_B8_o__o , \U_AHB/sel0_b5/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b5/or_B9_or_B10_B11_o_o );
  or \U_AHB/sel0_b5/or_or_or_B0_or_B1_B2  (\U_AHB/n114 [5], \U_AHB/sel0_b5/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b5/or_or_B6_or_B7_B8_o__o );
  and \U_AHB/sel0_b6/and_b0_0  (\U_AHB/sel0_b6/B0 , \U_AHB/h2h_hrdata [6], \U_AHB/n113 );
  and \U_AHB/sel0_b6/and_b0_1  (\U_AHB/sel0_b6/B1 , pnumcntA[6], \U_AHB/n111 );
  and \U_AHB/sel0_b6/and_b0_10  (\U_AHB/sel0_b6/B10 , pnumcnt1[6], \U_AHB/n84 );
  and \U_AHB/sel0_b6/and_b0_11  (\U_AHB/sel0_b6/B11 , pnumcnt0[6], \U_AHB/h2h_haddr [2]);
  and \U_AHB/sel0_b6/and_b0_2  (\U_AHB/sel0_b6/B2 , pnumcnt9[6], \U_AHB/n108 );
  and \U_AHB/sel0_b6/and_b0_3  (\U_AHB/sel0_b6/B3 , pnumcnt8[6], \U_AHB/n105 );
  and \U_AHB/sel0_b6/and_b0_4  (\U_AHB/sel0_b6/B4 , pnumcnt7[6], \U_AHB/n102 );
  and \U_AHB/sel0_b6/and_b0_5  (\U_AHB/sel0_b6/B5 , pnumcnt6[6], \U_AHB/n99 );
  and \U_AHB/sel0_b6/and_b0_6  (\U_AHB/sel0_b6/B6 , pnumcnt5[6], \U_AHB/n96 );
  and \U_AHB/sel0_b6/and_b0_7  (\U_AHB/sel0_b6/B7 , pnumcnt4[6], \U_AHB/n93 );
  and \U_AHB/sel0_b6/and_b0_8  (\U_AHB/sel0_b6/B8 , pnumcnt3[6], \U_AHB/n90 );
  and \U_AHB/sel0_b6/and_b0_9  (\U_AHB/sel0_b6/B9 , pnumcnt2[6], \U_AHB/n87 );
  or \U_AHB/sel0_b6/or_B0_or_B1_B2_o  (\U_AHB/sel0_b6/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b6/B0 , \U_AHB/sel0_b6/or_B1_B2_o );
  or \U_AHB/sel0_b6/or_B10_B11  (\U_AHB/sel0_b6/or_B10_B11_o , \U_AHB/sel0_b6/B10 , \U_AHB/sel0_b6/B11 );
  or \U_AHB/sel0_b6/or_B1_B2  (\U_AHB/sel0_b6/or_B1_B2_o , \U_AHB/sel0_b6/B1 , \U_AHB/sel0_b6/B2 );
  or \U_AHB/sel0_b6/or_B3_or_B4_B5_o  (\U_AHB/sel0_b6/or_B3_or_B4_B5_o_o , \U_AHB/sel0_b6/B3 , \U_AHB/sel0_b6/or_B4_B5_o );
  or \U_AHB/sel0_b6/or_B4_B5  (\U_AHB/sel0_b6/or_B4_B5_o , \U_AHB/sel0_b6/B4 , \U_AHB/sel0_b6/B5 );
  or \U_AHB/sel0_b6/or_B6_or_B7_B8_o  (\U_AHB/sel0_b6/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b6/B6 , \U_AHB/sel0_b6/or_B7_B8_o );
  or \U_AHB/sel0_b6/or_B7_B8  (\U_AHB/sel0_b6/or_B7_B8_o , \U_AHB/sel0_b6/B7 , \U_AHB/sel0_b6/B8 );
  or \U_AHB/sel0_b6/or_B9_or_B10_B11_o  (\U_AHB/sel0_b6/or_B9_or_B10_B11_o_o , \U_AHB/sel0_b6/B9 , \U_AHB/sel0_b6/or_B10_B11_o );
  or \U_AHB/sel0_b6/or_or_B0_or_B1_B2_o_  (\U_AHB/sel0_b6/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b6/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b6/or_B3_or_B4_B5_o_o );
  or \U_AHB/sel0_b6/or_or_B6_or_B7_B8_o_  (\U_AHB/sel0_b6/or_or_B6_or_B7_B8_o__o , \U_AHB/sel0_b6/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b6/or_B9_or_B10_B11_o_o );
  or \U_AHB/sel0_b6/or_or_or_B0_or_B1_B2  (\U_AHB/n114 [6], \U_AHB/sel0_b6/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b6/or_or_B6_or_B7_B8_o__o );
  and \U_AHB/sel0_b7/and_b0_0  (\U_AHB/sel0_b7/B0 , \U_AHB/h2h_hrdata [7], \U_AHB/n113 );
  and \U_AHB/sel0_b7/and_b0_1  (\U_AHB/sel0_b7/B1 , pnumcntA[7], \U_AHB/n111 );
  and \U_AHB/sel0_b7/and_b0_10  (\U_AHB/sel0_b7/B10 , pnumcnt1[7], \U_AHB/n84 );
  and \U_AHB/sel0_b7/and_b0_11  (\U_AHB/sel0_b7/B11 , pnumcnt0[7], \U_AHB/h2h_haddr [2]);
  and \U_AHB/sel0_b7/and_b0_2  (\U_AHB/sel0_b7/B2 , pnumcnt9[7], \U_AHB/n108 );
  and \U_AHB/sel0_b7/and_b0_3  (\U_AHB/sel0_b7/B3 , pnumcnt8[7], \U_AHB/n105 );
  and \U_AHB/sel0_b7/and_b0_4  (\U_AHB/sel0_b7/B4 , pnumcnt7[7], \U_AHB/n102 );
  and \U_AHB/sel0_b7/and_b0_5  (\U_AHB/sel0_b7/B5 , pnumcnt6[7], \U_AHB/n99 );
  and \U_AHB/sel0_b7/and_b0_6  (\U_AHB/sel0_b7/B6 , pnumcnt5[7], \U_AHB/n96 );
  and \U_AHB/sel0_b7/and_b0_7  (\U_AHB/sel0_b7/B7 , pnumcnt4[7], \U_AHB/n93 );
  and \U_AHB/sel0_b7/and_b0_8  (\U_AHB/sel0_b7/B8 , pnumcnt3[7], \U_AHB/n90 );
  and \U_AHB/sel0_b7/and_b0_9  (\U_AHB/sel0_b7/B9 , pnumcnt2[7], \U_AHB/n87 );
  or \U_AHB/sel0_b7/or_B0_or_B1_B2_o  (\U_AHB/sel0_b7/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b7/B0 , \U_AHB/sel0_b7/or_B1_B2_o );
  or \U_AHB/sel0_b7/or_B10_B11  (\U_AHB/sel0_b7/or_B10_B11_o , \U_AHB/sel0_b7/B10 , \U_AHB/sel0_b7/B11 );
  or \U_AHB/sel0_b7/or_B1_B2  (\U_AHB/sel0_b7/or_B1_B2_o , \U_AHB/sel0_b7/B1 , \U_AHB/sel0_b7/B2 );
  or \U_AHB/sel0_b7/or_B3_or_B4_B5_o  (\U_AHB/sel0_b7/or_B3_or_B4_B5_o_o , \U_AHB/sel0_b7/B3 , \U_AHB/sel0_b7/or_B4_B5_o );
  or \U_AHB/sel0_b7/or_B4_B5  (\U_AHB/sel0_b7/or_B4_B5_o , \U_AHB/sel0_b7/B4 , \U_AHB/sel0_b7/B5 );
  or \U_AHB/sel0_b7/or_B6_or_B7_B8_o  (\U_AHB/sel0_b7/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b7/B6 , \U_AHB/sel0_b7/or_B7_B8_o );
  or \U_AHB/sel0_b7/or_B7_B8  (\U_AHB/sel0_b7/or_B7_B8_o , \U_AHB/sel0_b7/B7 , \U_AHB/sel0_b7/B8 );
  or \U_AHB/sel0_b7/or_B9_or_B10_B11_o  (\U_AHB/sel0_b7/or_B9_or_B10_B11_o_o , \U_AHB/sel0_b7/B9 , \U_AHB/sel0_b7/or_B10_B11_o );
  or \U_AHB/sel0_b7/or_or_B0_or_B1_B2_o_  (\U_AHB/sel0_b7/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b7/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b7/or_B3_or_B4_B5_o_o );
  or \U_AHB/sel0_b7/or_or_B6_or_B7_B8_o_  (\U_AHB/sel0_b7/or_or_B6_or_B7_B8_o__o , \U_AHB/sel0_b7/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b7/or_B9_or_B10_B11_o_o );
  or \U_AHB/sel0_b7/or_or_or_B0_or_B1_B2  (\U_AHB/n114 [7], \U_AHB/sel0_b7/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b7/or_or_B6_or_B7_B8_o__o );
  and \U_AHB/sel0_b8/and_b0_0  (\U_AHB/sel0_b8/B0 , \U_AHB/h2h_hrdata [8], \U_AHB/n113 );
  and \U_AHB/sel0_b8/and_b0_1  (\U_AHB/sel0_b8/B1 , pnumcntA[8], \U_AHB/n111 );
  and \U_AHB/sel0_b8/and_b0_10  (\U_AHB/sel0_b8/B10 , pnumcnt1[8], \U_AHB/n84 );
  and \U_AHB/sel0_b8/and_b0_11  (\U_AHB/sel0_b8/B11 , pnumcnt0[8], \U_AHB/h2h_haddr [2]);
  and \U_AHB/sel0_b8/and_b0_2  (\U_AHB/sel0_b8/B2 , pnumcnt9[8], \U_AHB/n108 );
  and \U_AHB/sel0_b8/and_b0_3  (\U_AHB/sel0_b8/B3 , pnumcnt8[8], \U_AHB/n105 );
  and \U_AHB/sel0_b8/and_b0_4  (\U_AHB/sel0_b8/B4 , pnumcnt7[8], \U_AHB/n102 );
  and \U_AHB/sel0_b8/and_b0_5  (\U_AHB/sel0_b8/B5 , pnumcnt6[8], \U_AHB/n99 );
  and \U_AHB/sel0_b8/and_b0_6  (\U_AHB/sel0_b8/B6 , pnumcnt5[8], \U_AHB/n96 );
  and \U_AHB/sel0_b8/and_b0_7  (\U_AHB/sel0_b8/B7 , pnumcnt4[8], \U_AHB/n93 );
  and \U_AHB/sel0_b8/and_b0_8  (\U_AHB/sel0_b8/B8 , pnumcnt3[8], \U_AHB/n90 );
  and \U_AHB/sel0_b8/and_b0_9  (\U_AHB/sel0_b8/B9 , pnumcnt2[8], \U_AHB/n87 );
  or \U_AHB/sel0_b8/or_B0_or_B1_B2_o  (\U_AHB/sel0_b8/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b8/B0 , \U_AHB/sel0_b8/or_B1_B2_o );
  or \U_AHB/sel0_b8/or_B10_B11  (\U_AHB/sel0_b8/or_B10_B11_o , \U_AHB/sel0_b8/B10 , \U_AHB/sel0_b8/B11 );
  or \U_AHB/sel0_b8/or_B1_B2  (\U_AHB/sel0_b8/or_B1_B2_o , \U_AHB/sel0_b8/B1 , \U_AHB/sel0_b8/B2 );
  or \U_AHB/sel0_b8/or_B3_or_B4_B5_o  (\U_AHB/sel0_b8/or_B3_or_B4_B5_o_o , \U_AHB/sel0_b8/B3 , \U_AHB/sel0_b8/or_B4_B5_o );
  or \U_AHB/sel0_b8/or_B4_B5  (\U_AHB/sel0_b8/or_B4_B5_o , \U_AHB/sel0_b8/B4 , \U_AHB/sel0_b8/B5 );
  or \U_AHB/sel0_b8/or_B6_or_B7_B8_o  (\U_AHB/sel0_b8/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b8/B6 , \U_AHB/sel0_b8/or_B7_B8_o );
  or \U_AHB/sel0_b8/or_B7_B8  (\U_AHB/sel0_b8/or_B7_B8_o , \U_AHB/sel0_b8/B7 , \U_AHB/sel0_b8/B8 );
  or \U_AHB/sel0_b8/or_B9_or_B10_B11_o  (\U_AHB/sel0_b8/or_B9_or_B10_B11_o_o , \U_AHB/sel0_b8/B9 , \U_AHB/sel0_b8/or_B10_B11_o );
  or \U_AHB/sel0_b8/or_or_B0_or_B1_B2_o_  (\U_AHB/sel0_b8/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b8/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b8/or_B3_or_B4_B5_o_o );
  or \U_AHB/sel0_b8/or_or_B6_or_B7_B8_o_  (\U_AHB/sel0_b8/or_or_B6_or_B7_B8_o__o , \U_AHB/sel0_b8/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b8/or_B9_or_B10_B11_o_o );
  or \U_AHB/sel0_b8/or_or_or_B0_or_B1_B2  (\U_AHB/n114 [8], \U_AHB/sel0_b8/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b8/or_or_B6_or_B7_B8_o__o );
  and \U_AHB/sel0_b9/and_b0_0  (\U_AHB/sel0_b9/B0 , \U_AHB/h2h_hrdata [9], \U_AHB/n113 );
  and \U_AHB/sel0_b9/and_b0_1  (\U_AHB/sel0_b9/B1 , pnumcntA[9], \U_AHB/n111 );
  and \U_AHB/sel0_b9/and_b0_10  (\U_AHB/sel0_b9/B10 , pnumcnt1[9], \U_AHB/n84 );
  and \U_AHB/sel0_b9/and_b0_11  (\U_AHB/sel0_b9/B11 , pnumcnt0[9], \U_AHB/h2h_haddr [2]);
  and \U_AHB/sel0_b9/and_b0_2  (\U_AHB/sel0_b9/B2 , pnumcnt9[9], \U_AHB/n108 );
  and \U_AHB/sel0_b9/and_b0_3  (\U_AHB/sel0_b9/B3 , pnumcnt8[9], \U_AHB/n105 );
  and \U_AHB/sel0_b9/and_b0_4  (\U_AHB/sel0_b9/B4 , pnumcnt7[9], \U_AHB/n102 );
  and \U_AHB/sel0_b9/and_b0_5  (\U_AHB/sel0_b9/B5 , pnumcnt6[9], \U_AHB/n99 );
  and \U_AHB/sel0_b9/and_b0_6  (\U_AHB/sel0_b9/B6 , pnumcnt5[9], \U_AHB/n96 );
  and \U_AHB/sel0_b9/and_b0_7  (\U_AHB/sel0_b9/B7 , pnumcnt4[9], \U_AHB/n93 );
  and \U_AHB/sel0_b9/and_b0_8  (\U_AHB/sel0_b9/B8 , pnumcnt3[9], \U_AHB/n90 );
  and \U_AHB/sel0_b9/and_b0_9  (\U_AHB/sel0_b9/B9 , pnumcnt2[9], \U_AHB/n87 );
  or \U_AHB/sel0_b9/or_B0_or_B1_B2_o  (\U_AHB/sel0_b9/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b9/B0 , \U_AHB/sel0_b9/or_B1_B2_o );
  or \U_AHB/sel0_b9/or_B10_B11  (\U_AHB/sel0_b9/or_B10_B11_o , \U_AHB/sel0_b9/B10 , \U_AHB/sel0_b9/B11 );
  or \U_AHB/sel0_b9/or_B1_B2  (\U_AHB/sel0_b9/or_B1_B2_o , \U_AHB/sel0_b9/B1 , \U_AHB/sel0_b9/B2 );
  or \U_AHB/sel0_b9/or_B3_or_B4_B5_o  (\U_AHB/sel0_b9/or_B3_or_B4_B5_o_o , \U_AHB/sel0_b9/B3 , \U_AHB/sel0_b9/or_B4_B5_o );
  or \U_AHB/sel0_b9/or_B4_B5  (\U_AHB/sel0_b9/or_B4_B5_o , \U_AHB/sel0_b9/B4 , \U_AHB/sel0_b9/B5 );
  or \U_AHB/sel0_b9/or_B6_or_B7_B8_o  (\U_AHB/sel0_b9/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b9/B6 , \U_AHB/sel0_b9/or_B7_B8_o );
  or \U_AHB/sel0_b9/or_B7_B8  (\U_AHB/sel0_b9/or_B7_B8_o , \U_AHB/sel0_b9/B7 , \U_AHB/sel0_b9/B8 );
  or \U_AHB/sel0_b9/or_B9_or_B10_B11_o  (\U_AHB/sel0_b9/or_B9_or_B10_B11_o_o , \U_AHB/sel0_b9/B9 , \U_AHB/sel0_b9/or_B10_B11_o );
  or \U_AHB/sel0_b9/or_or_B0_or_B1_B2_o_  (\U_AHB/sel0_b9/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b9/or_B0_or_B1_B2_o_o , \U_AHB/sel0_b9/or_B3_or_B4_B5_o_o );
  or \U_AHB/sel0_b9/or_or_B6_or_B7_B8_o_  (\U_AHB/sel0_b9/or_or_B6_or_B7_B8_o__o , \U_AHB/sel0_b9/or_B6_or_B7_B8_o_o , \U_AHB/sel0_b9/or_B9_or_B10_B11_o_o );
  or \U_AHB/sel0_b9/or_or_or_B0_or_B1_B2  (\U_AHB/n114 [9], \U_AHB/sel0_b9/or_or_B0_or_B1_B2_o__o , \U_AHB/sel0_b9/or_or_B6_or_B7_B8_o__o );
  and \U_AHB/sel1_b0/and_b0_0  (\U_AHB/sel1_b0/B0 , \U_AHB/h2h_hrdata [0], \U_AHB/n104 );
  and \U_AHB/sel1_b0/and_b0_1  (\U_AHB/sel1_b0/B1 , limit_r[0], \U_AHB/n102 );
  and \U_AHB/sel1_b0/and_b0_3  (\U_AHB/sel1_b0/B3 , pwm_state_read[0], \U_AHB/n96 );
  and \U_AHB/sel1_b0/and_b0_4  (\U_AHB/sel1_b0/B4 , pnumcntF[0], \U_AHB/n93 );
  and \U_AHB/sel1_b0/and_b0_5  (\U_AHB/sel1_b0/B5 , pnumcntE[0], \U_AHB/n90 );
  and \U_AHB/sel1_b0/and_b0_6  (\U_AHB/sel1_b0/B6 , pnumcntD[0], \U_AHB/n87 );
  and \U_AHB/sel1_b0/and_b0_7  (\U_AHB/sel1_b0/B7 , pnumcntC[0], \U_AHB/n84 );
  and \U_AHB/sel1_b0/and_b0_8  (\U_AHB/sel1_b0/B8 , pnumcntB[0], \U_AHB/h2h_haddr [2]);
  or \U_AHB/sel1_b0/or_B0_B1  (\U_AHB/sel1_b0/or_B0_B1_o , \U_AHB/sel1_b0/B0 , \U_AHB/sel1_b0/B1 );
  or \U_AHB/sel1_b0/or_B4_B5  (\U_AHB/sel1_b0/or_B4_B5_o , \U_AHB/sel1_b0/B4 , \U_AHB/sel1_b0/B5 );
  or \U_AHB/sel1_b0/or_B6_or_B7_B8_o  (\U_AHB/sel1_b0/or_B6_or_B7_B8_o_o , \U_AHB/sel1_b0/B6 , \U_AHB/sel1_b0/or_B7_B8_o );
  or \U_AHB/sel1_b0/or_B7_B8  (\U_AHB/sel1_b0/or_B7_B8_o , \U_AHB/sel1_b0/B7 , \U_AHB/sel1_b0/B8 );
  or \U_AHB/sel1_b0/or_or_B0_B1_o_or_B2_  (\U_AHB/sel1_b0/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b0/or_B0_B1_o , \U_AHB/sel1_b0/B3 );
  or \U_AHB/sel1_b0/or_or_B4_B5_o_or_B6_  (\U_AHB/sel1_b0/or_or_B4_B5_o_or_B6__o , \U_AHB/sel1_b0/or_B4_B5_o , \U_AHB/sel1_b0/or_B6_or_B7_B8_o_o );
  or \U_AHB/sel1_b0/or_or_or_B0_B1_o_or_  (\U_AHB/n116 [0], \U_AHB/sel1_b0/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b0/or_or_B4_B5_o_or_B6__o );
  and \U_AHB/sel1_b1/and_b0_0  (\U_AHB/sel1_b1/B0 , \U_AHB/h2h_hrdata [1], \U_AHB/n104 );
  and \U_AHB/sel1_b1/and_b0_1  (\U_AHB/sel1_b1/B1 , limit_r[1], \U_AHB/n102 );
  and \U_AHB/sel1_b1/and_b0_3  (\U_AHB/sel1_b1/B3 , pwm_state_read[1], \U_AHB/n96 );
  and \U_AHB/sel1_b1/and_b0_4  (\U_AHB/sel1_b1/B4 , pnumcntF[1], \U_AHB/n93 );
  and \U_AHB/sel1_b1/and_b0_5  (\U_AHB/sel1_b1/B5 , pnumcntE[1], \U_AHB/n90 );
  and \U_AHB/sel1_b1/and_b0_6  (\U_AHB/sel1_b1/B6 , pnumcntD[1], \U_AHB/n87 );
  and \U_AHB/sel1_b1/and_b0_7  (\U_AHB/sel1_b1/B7 , pnumcntC[1], \U_AHB/n84 );
  and \U_AHB/sel1_b1/and_b0_8  (\U_AHB/sel1_b1/B8 , pnumcntB[1], \U_AHB/h2h_haddr [2]);
  or \U_AHB/sel1_b1/or_B0_B1  (\U_AHB/sel1_b1/or_B0_B1_o , \U_AHB/sel1_b1/B0 , \U_AHB/sel1_b1/B1 );
  or \U_AHB/sel1_b1/or_B4_B5  (\U_AHB/sel1_b1/or_B4_B5_o , \U_AHB/sel1_b1/B4 , \U_AHB/sel1_b1/B5 );
  or \U_AHB/sel1_b1/or_B6_or_B7_B8_o  (\U_AHB/sel1_b1/or_B6_or_B7_B8_o_o , \U_AHB/sel1_b1/B6 , \U_AHB/sel1_b1/or_B7_B8_o );
  or \U_AHB/sel1_b1/or_B7_B8  (\U_AHB/sel1_b1/or_B7_B8_o , \U_AHB/sel1_b1/B7 , \U_AHB/sel1_b1/B8 );
  or \U_AHB/sel1_b1/or_or_B0_B1_o_or_B2_  (\U_AHB/sel1_b1/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b1/or_B0_B1_o , \U_AHB/sel1_b1/B3 );
  or \U_AHB/sel1_b1/or_or_B4_B5_o_or_B6_  (\U_AHB/sel1_b1/or_or_B4_B5_o_or_B6__o , \U_AHB/sel1_b1/or_B4_B5_o , \U_AHB/sel1_b1/or_B6_or_B7_B8_o_o );
  or \U_AHB/sel1_b1/or_or_or_B0_B1_o_or_  (\U_AHB/n116 [1], \U_AHB/sel1_b1/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b1/or_or_B4_B5_o_or_B6__o );
  and \U_AHB/sel1_b10/and_b0_0  (\U_AHB/sel1_b10/B0 , \U_AHB/h2h_hrdata [10], \U_AHB/n104 );
  and \U_AHB/sel1_b10/and_b0_1  (\U_AHB/sel1_b10/B1 , limit_r[10], \U_AHB/n102 );
  and \U_AHB/sel1_b10/and_b0_3  (\U_AHB/sel1_b10/B3 , pwm_state_read[10], \U_AHB/n96 );
  and \U_AHB/sel1_b10/and_b0_4  (\U_AHB/sel1_b10/B4 , pnumcntF[10], \U_AHB/n93 );
  and \U_AHB/sel1_b10/and_b0_5  (\U_AHB/sel1_b10/B5 , pnumcntE[10], \U_AHB/n90 );
  and \U_AHB/sel1_b10/and_b0_6  (\U_AHB/sel1_b10/B6 , pnumcntD[10], \U_AHB/n87 );
  and \U_AHB/sel1_b10/and_b0_7  (\U_AHB/sel1_b10/B7 , pnumcntC[10], \U_AHB/n84 );
  and \U_AHB/sel1_b10/and_b0_8  (\U_AHB/sel1_b10/B8 , pnumcntB[10], \U_AHB/h2h_haddr [2]);
  or \U_AHB/sel1_b10/or_B0_B1  (\U_AHB/sel1_b10/or_B0_B1_o , \U_AHB/sel1_b10/B0 , \U_AHB/sel1_b10/B1 );
  or \U_AHB/sel1_b10/or_B4_B5  (\U_AHB/sel1_b10/or_B4_B5_o , \U_AHB/sel1_b10/B4 , \U_AHB/sel1_b10/B5 );
  or \U_AHB/sel1_b10/or_B6_or_B7_B8_o  (\U_AHB/sel1_b10/or_B6_or_B7_B8_o_o , \U_AHB/sel1_b10/B6 , \U_AHB/sel1_b10/or_B7_B8_o );
  or \U_AHB/sel1_b10/or_B7_B8  (\U_AHB/sel1_b10/or_B7_B8_o , \U_AHB/sel1_b10/B7 , \U_AHB/sel1_b10/B8 );
  or \U_AHB/sel1_b10/or_or_B0_B1_o_or_B2_  (\U_AHB/sel1_b10/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b10/or_B0_B1_o , \U_AHB/sel1_b10/B3 );
  or \U_AHB/sel1_b10/or_or_B4_B5_o_or_B6_  (\U_AHB/sel1_b10/or_or_B4_B5_o_or_B6__o , \U_AHB/sel1_b10/or_B4_B5_o , \U_AHB/sel1_b10/or_B6_or_B7_B8_o_o );
  or \U_AHB/sel1_b10/or_or_or_B0_B1_o_or_  (\U_AHB/n116 [10], \U_AHB/sel1_b10/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b10/or_or_B4_B5_o_or_B6__o );
  and \U_AHB/sel1_b11/and_b0_0  (\U_AHB/sel1_b11/B0 , \U_AHB/h2h_hrdata [11], \U_AHB/n104 );
  and \U_AHB/sel1_b11/and_b0_1  (\U_AHB/sel1_b11/B1 , limit_r[11], \U_AHB/n102 );
  and \U_AHB/sel1_b11/and_b0_3  (\U_AHB/sel1_b11/B3 , pwm_state_read[11], \U_AHB/n96 );
  and \U_AHB/sel1_b11/and_b0_4  (\U_AHB/sel1_b11/B4 , pnumcntF[11], \U_AHB/n93 );
  and \U_AHB/sel1_b11/and_b0_5  (\U_AHB/sel1_b11/B5 , pnumcntE[11], \U_AHB/n90 );
  and \U_AHB/sel1_b11/and_b0_6  (\U_AHB/sel1_b11/B6 , pnumcntD[11], \U_AHB/n87 );
  and \U_AHB/sel1_b11/and_b0_7  (\U_AHB/sel1_b11/B7 , pnumcntC[11], \U_AHB/n84 );
  and \U_AHB/sel1_b11/and_b0_8  (\U_AHB/sel1_b11/B8 , pnumcntB[11], \U_AHB/h2h_haddr [2]);
  or \U_AHB/sel1_b11/or_B0_B1  (\U_AHB/sel1_b11/or_B0_B1_o , \U_AHB/sel1_b11/B0 , \U_AHB/sel1_b11/B1 );
  or \U_AHB/sel1_b11/or_B4_B5  (\U_AHB/sel1_b11/or_B4_B5_o , \U_AHB/sel1_b11/B4 , \U_AHB/sel1_b11/B5 );
  or \U_AHB/sel1_b11/or_B6_or_B7_B8_o  (\U_AHB/sel1_b11/or_B6_or_B7_B8_o_o , \U_AHB/sel1_b11/B6 , \U_AHB/sel1_b11/or_B7_B8_o );
  or \U_AHB/sel1_b11/or_B7_B8  (\U_AHB/sel1_b11/or_B7_B8_o , \U_AHB/sel1_b11/B7 , \U_AHB/sel1_b11/B8 );
  or \U_AHB/sel1_b11/or_or_B0_B1_o_or_B2_  (\U_AHB/sel1_b11/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b11/or_B0_B1_o , \U_AHB/sel1_b11/B3 );
  or \U_AHB/sel1_b11/or_or_B4_B5_o_or_B6_  (\U_AHB/sel1_b11/or_or_B4_B5_o_or_B6__o , \U_AHB/sel1_b11/or_B4_B5_o , \U_AHB/sel1_b11/or_B6_or_B7_B8_o_o );
  or \U_AHB/sel1_b11/or_or_or_B0_B1_o_or_  (\U_AHB/n116 [11], \U_AHB/sel1_b11/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b11/or_or_B4_B5_o_or_B6__o );
  and \U_AHB/sel1_b12/and_b0_0  (\U_AHB/sel1_b12/B0 , \U_AHB/h2h_hrdata [12], \U_AHB/n104 );
  and \U_AHB/sel1_b12/and_b0_1  (\U_AHB/sel1_b12/B1 , limit_r[12], \U_AHB/n102 );
  and \U_AHB/sel1_b12/and_b0_3  (\U_AHB/sel1_b12/B3 , pwm_state_read[12], \U_AHB/n96 );
  and \U_AHB/sel1_b12/and_b0_4  (\U_AHB/sel1_b12/B4 , pnumcntF[12], \U_AHB/n93 );
  and \U_AHB/sel1_b12/and_b0_5  (\U_AHB/sel1_b12/B5 , pnumcntE[12], \U_AHB/n90 );
  and \U_AHB/sel1_b12/and_b0_6  (\U_AHB/sel1_b12/B6 , pnumcntD[12], \U_AHB/n87 );
  and \U_AHB/sel1_b12/and_b0_7  (\U_AHB/sel1_b12/B7 , pnumcntC[12], \U_AHB/n84 );
  and \U_AHB/sel1_b12/and_b0_8  (\U_AHB/sel1_b12/B8 , pnumcntB[12], \U_AHB/h2h_haddr [2]);
  or \U_AHB/sel1_b12/or_B0_B1  (\U_AHB/sel1_b12/or_B0_B1_o , \U_AHB/sel1_b12/B0 , \U_AHB/sel1_b12/B1 );
  or \U_AHB/sel1_b12/or_B4_B5  (\U_AHB/sel1_b12/or_B4_B5_o , \U_AHB/sel1_b12/B4 , \U_AHB/sel1_b12/B5 );
  or \U_AHB/sel1_b12/or_B6_or_B7_B8_o  (\U_AHB/sel1_b12/or_B6_or_B7_B8_o_o , \U_AHB/sel1_b12/B6 , \U_AHB/sel1_b12/or_B7_B8_o );
  or \U_AHB/sel1_b12/or_B7_B8  (\U_AHB/sel1_b12/or_B7_B8_o , \U_AHB/sel1_b12/B7 , \U_AHB/sel1_b12/B8 );
  or \U_AHB/sel1_b12/or_or_B0_B1_o_or_B2_  (\U_AHB/sel1_b12/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b12/or_B0_B1_o , \U_AHB/sel1_b12/B3 );
  or \U_AHB/sel1_b12/or_or_B4_B5_o_or_B6_  (\U_AHB/sel1_b12/or_or_B4_B5_o_or_B6__o , \U_AHB/sel1_b12/or_B4_B5_o , \U_AHB/sel1_b12/or_B6_or_B7_B8_o_o );
  or \U_AHB/sel1_b12/or_or_or_B0_B1_o_or_  (\U_AHB/n116 [12], \U_AHB/sel1_b12/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b12/or_or_B4_B5_o_or_B6__o );
  and \U_AHB/sel1_b13/and_b0_0  (\U_AHB/sel1_b13/B0 , \U_AHB/h2h_hrdata [13], \U_AHB/n104 );
  and \U_AHB/sel1_b13/and_b0_1  (\U_AHB/sel1_b13/B1 , limit_r[13], \U_AHB/n102 );
  and \U_AHB/sel1_b13/and_b0_3  (\U_AHB/sel1_b13/B3 , pwm_state_read[13], \U_AHB/n96 );
  and \U_AHB/sel1_b13/and_b0_4  (\U_AHB/sel1_b13/B4 , pnumcntF[13], \U_AHB/n93 );
  and \U_AHB/sel1_b13/and_b0_5  (\U_AHB/sel1_b13/B5 , pnumcntE[13], \U_AHB/n90 );
  and \U_AHB/sel1_b13/and_b0_6  (\U_AHB/sel1_b13/B6 , pnumcntD[13], \U_AHB/n87 );
  and \U_AHB/sel1_b13/and_b0_7  (\U_AHB/sel1_b13/B7 , pnumcntC[13], \U_AHB/n84 );
  and \U_AHB/sel1_b13/and_b0_8  (\U_AHB/sel1_b13/B8 , pnumcntB[13], \U_AHB/h2h_haddr [2]);
  or \U_AHB/sel1_b13/or_B0_B1  (\U_AHB/sel1_b13/or_B0_B1_o , \U_AHB/sel1_b13/B0 , \U_AHB/sel1_b13/B1 );
  or \U_AHB/sel1_b13/or_B4_B5  (\U_AHB/sel1_b13/or_B4_B5_o , \U_AHB/sel1_b13/B4 , \U_AHB/sel1_b13/B5 );
  or \U_AHB/sel1_b13/or_B6_or_B7_B8_o  (\U_AHB/sel1_b13/or_B6_or_B7_B8_o_o , \U_AHB/sel1_b13/B6 , \U_AHB/sel1_b13/or_B7_B8_o );
  or \U_AHB/sel1_b13/or_B7_B8  (\U_AHB/sel1_b13/or_B7_B8_o , \U_AHB/sel1_b13/B7 , \U_AHB/sel1_b13/B8 );
  or \U_AHB/sel1_b13/or_or_B0_B1_o_or_B2_  (\U_AHB/sel1_b13/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b13/or_B0_B1_o , \U_AHB/sel1_b13/B3 );
  or \U_AHB/sel1_b13/or_or_B4_B5_o_or_B6_  (\U_AHB/sel1_b13/or_or_B4_B5_o_or_B6__o , \U_AHB/sel1_b13/or_B4_B5_o , \U_AHB/sel1_b13/or_B6_or_B7_B8_o_o );
  or \U_AHB/sel1_b13/or_or_or_B0_B1_o_or_  (\U_AHB/n116 [13], \U_AHB/sel1_b13/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b13/or_or_B4_B5_o_or_B6__o );
  and \U_AHB/sel1_b14/and_b0_0  (\U_AHB/sel1_b14/B0 , \U_AHB/h2h_hrdata [14], \U_AHB/n104 );
  and \U_AHB/sel1_b14/and_b0_1  (\U_AHB/sel1_b14/B1 , limit_r[14], \U_AHB/n102 );
  and \U_AHB/sel1_b14/and_b0_3  (\U_AHB/sel1_b14/B3 , pwm_state_read[14], \U_AHB/n96 );
  and \U_AHB/sel1_b14/and_b0_4  (\U_AHB/sel1_b14/B4 , pnumcntF[14], \U_AHB/n93 );
  and \U_AHB/sel1_b14/and_b0_5  (\U_AHB/sel1_b14/B5 , pnumcntE[14], \U_AHB/n90 );
  and \U_AHB/sel1_b14/and_b0_6  (\U_AHB/sel1_b14/B6 , pnumcntD[14], \U_AHB/n87 );
  and \U_AHB/sel1_b14/and_b0_7  (\U_AHB/sel1_b14/B7 , pnumcntC[14], \U_AHB/n84 );
  and \U_AHB/sel1_b14/and_b0_8  (\U_AHB/sel1_b14/B8 , pnumcntB[14], \U_AHB/h2h_haddr [2]);
  or \U_AHB/sel1_b14/or_B0_B1  (\U_AHB/sel1_b14/or_B0_B1_o , \U_AHB/sel1_b14/B0 , \U_AHB/sel1_b14/B1 );
  or \U_AHB/sel1_b14/or_B4_B5  (\U_AHB/sel1_b14/or_B4_B5_o , \U_AHB/sel1_b14/B4 , \U_AHB/sel1_b14/B5 );
  or \U_AHB/sel1_b14/or_B6_or_B7_B8_o  (\U_AHB/sel1_b14/or_B6_or_B7_B8_o_o , \U_AHB/sel1_b14/B6 , \U_AHB/sel1_b14/or_B7_B8_o );
  or \U_AHB/sel1_b14/or_B7_B8  (\U_AHB/sel1_b14/or_B7_B8_o , \U_AHB/sel1_b14/B7 , \U_AHB/sel1_b14/B8 );
  or \U_AHB/sel1_b14/or_or_B0_B1_o_or_B2_  (\U_AHB/sel1_b14/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b14/or_B0_B1_o , \U_AHB/sel1_b14/B3 );
  or \U_AHB/sel1_b14/or_or_B4_B5_o_or_B6_  (\U_AHB/sel1_b14/or_or_B4_B5_o_or_B6__o , \U_AHB/sel1_b14/or_B4_B5_o , \U_AHB/sel1_b14/or_B6_or_B7_B8_o_o );
  or \U_AHB/sel1_b14/or_or_or_B0_B1_o_or_  (\U_AHB/n116 [14], \U_AHB/sel1_b14/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b14/or_or_B4_B5_o_or_B6__o );
  and \U_AHB/sel1_b15/and_b0_0  (\U_AHB/sel1_b15/B0 , \U_AHB/h2h_hrdata [15], \U_AHB/n104 );
  and \U_AHB/sel1_b15/and_b0_1  (\U_AHB/sel1_b15/B1 , limit_r[15], \U_AHB/n102 );
  and \U_AHB/sel1_b15/and_b0_3  (\U_AHB/sel1_b15/B3 , pwm_state_read[15], \U_AHB/n96 );
  and \U_AHB/sel1_b15/and_b0_4  (\U_AHB/sel1_b15/B4 , pnumcntF[15], \U_AHB/n93 );
  and \U_AHB/sel1_b15/and_b0_5  (\U_AHB/sel1_b15/B5 , pnumcntE[15], \U_AHB/n90 );
  and \U_AHB/sel1_b15/and_b0_6  (\U_AHB/sel1_b15/B6 , pnumcntD[15], \U_AHB/n87 );
  and \U_AHB/sel1_b15/and_b0_7  (\U_AHB/sel1_b15/B7 , pnumcntC[15], \U_AHB/n84 );
  and \U_AHB/sel1_b15/and_b0_8  (\U_AHB/sel1_b15/B8 , pnumcntB[15], \U_AHB/h2h_haddr [2]);
  or \U_AHB/sel1_b15/or_B0_B1  (\U_AHB/sel1_b15/or_B0_B1_o , \U_AHB/sel1_b15/B0 , \U_AHB/sel1_b15/B1 );
  or \U_AHB/sel1_b15/or_B4_B5  (\U_AHB/sel1_b15/or_B4_B5_o , \U_AHB/sel1_b15/B4 , \U_AHB/sel1_b15/B5 );
  or \U_AHB/sel1_b15/or_B6_or_B7_B8_o  (\U_AHB/sel1_b15/or_B6_or_B7_B8_o_o , \U_AHB/sel1_b15/B6 , \U_AHB/sel1_b15/or_B7_B8_o );
  or \U_AHB/sel1_b15/or_B7_B8  (\U_AHB/sel1_b15/or_B7_B8_o , \U_AHB/sel1_b15/B7 , \U_AHB/sel1_b15/B8 );
  or \U_AHB/sel1_b15/or_or_B0_B1_o_or_B2_  (\U_AHB/sel1_b15/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b15/or_B0_B1_o , \U_AHB/sel1_b15/B3 );
  or \U_AHB/sel1_b15/or_or_B4_B5_o_or_B6_  (\U_AHB/sel1_b15/or_or_B4_B5_o_or_B6__o , \U_AHB/sel1_b15/or_B4_B5_o , \U_AHB/sel1_b15/or_B6_or_B7_B8_o_o );
  or \U_AHB/sel1_b15/or_or_or_B0_B1_o_or_  (\U_AHB/n116 [15], \U_AHB/sel1_b15/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b15/or_or_B4_B5_o_or_B6__o );
  and \U_AHB/sel1_b16/and_b0_0  (\U_AHB/sel1_b16/B0 , \U_AHB/h2h_hrdata [16], \U_AHB/n104 );
  and \U_AHB/sel1_b16/and_b0_1  (\U_AHB/sel1_b16/B1 , limit_l[0], \U_AHB/n102 );
  and \U_AHB/sel1_b16/and_b0_4  (\U_AHB/sel1_b16/B4 , pnumcntF[16], \U_AHB/n93 );
  and \U_AHB/sel1_b16/and_b0_5  (\U_AHB/sel1_b16/B5 , pnumcntE[16], \U_AHB/n90 );
  and \U_AHB/sel1_b16/and_b0_6  (\U_AHB/sel1_b16/B6 , pnumcntD[16], \U_AHB/n87 );
  and \U_AHB/sel1_b16/and_b0_7  (\U_AHB/sel1_b16/B7 , pnumcntC[16], \U_AHB/n84 );
  and \U_AHB/sel1_b16/and_b0_8  (\U_AHB/sel1_b16/B8 , pnumcntB[16], \U_AHB/h2h_haddr [2]);
  or \U_AHB/sel1_b16/or_B0_B1  (\U_AHB/sel1_b16/or_B0_B1_o , \U_AHB/sel1_b16/B0 , \U_AHB/sel1_b16/B1 );
  or \U_AHB/sel1_b16/or_B4_B5  (\U_AHB/sel1_b16/or_B4_B5_o , \U_AHB/sel1_b16/B4 , \U_AHB/sel1_b16/B5 );
  or \U_AHB/sel1_b16/or_B6_or_B7_B8_o  (\U_AHB/sel1_b16/or_B6_or_B7_B8_o_o , \U_AHB/sel1_b16/B6 , \U_AHB/sel1_b16/or_B7_B8_o );
  or \U_AHB/sel1_b16/or_B7_B8  (\U_AHB/sel1_b16/or_B7_B8_o , \U_AHB/sel1_b16/B7 , \U_AHB/sel1_b16/B8 );
  or \U_AHB/sel1_b16/or_or_B0_B1_o_or_B2_  (\U_AHB/sel1_b16/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b16/or_B0_B1_o , \U_AHB/sel1_b0/B3 );
  or \U_AHB/sel1_b16/or_or_B4_B5_o_or_B6_  (\U_AHB/sel1_b16/or_or_B4_B5_o_or_B6__o , \U_AHB/sel1_b16/or_B4_B5_o , \U_AHB/sel1_b16/or_B6_or_B7_B8_o_o );
  or \U_AHB/sel1_b16/or_or_or_B0_B1_o_or_  (\U_AHB/n116 [16], \U_AHB/sel1_b16/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b16/or_or_B4_B5_o_or_B6__o );
  and \U_AHB/sel1_b17/and_b0_0  (\U_AHB/sel1_b17/B0 , \U_AHB/h2h_hrdata [17], \U_AHB/n104 );
  and \U_AHB/sel1_b17/and_b0_1  (\U_AHB/sel1_b17/B1 , limit_l[1], \U_AHB/n102 );
  and \U_AHB/sel1_b17/and_b0_4  (\U_AHB/sel1_b17/B4 , pnumcntF[17], \U_AHB/n93 );
  and \U_AHB/sel1_b17/and_b0_5  (\U_AHB/sel1_b17/B5 , pnumcntE[17], \U_AHB/n90 );
  and \U_AHB/sel1_b17/and_b0_6  (\U_AHB/sel1_b17/B6 , pnumcntD[17], \U_AHB/n87 );
  and \U_AHB/sel1_b17/and_b0_7  (\U_AHB/sel1_b17/B7 , pnumcntC[17], \U_AHB/n84 );
  and \U_AHB/sel1_b17/and_b0_8  (\U_AHB/sel1_b17/B8 , pnumcntB[17], \U_AHB/h2h_haddr [2]);
  or \U_AHB/sel1_b17/or_B0_B1  (\U_AHB/sel1_b17/or_B0_B1_o , \U_AHB/sel1_b17/B0 , \U_AHB/sel1_b17/B1 );
  or \U_AHB/sel1_b17/or_B4_B5  (\U_AHB/sel1_b17/or_B4_B5_o , \U_AHB/sel1_b17/B4 , \U_AHB/sel1_b17/B5 );
  or \U_AHB/sel1_b17/or_B6_or_B7_B8_o  (\U_AHB/sel1_b17/or_B6_or_B7_B8_o_o , \U_AHB/sel1_b17/B6 , \U_AHB/sel1_b17/or_B7_B8_o );
  or \U_AHB/sel1_b17/or_B7_B8  (\U_AHB/sel1_b17/or_B7_B8_o , \U_AHB/sel1_b17/B7 , \U_AHB/sel1_b17/B8 );
  or \U_AHB/sel1_b17/or_or_B0_B1_o_or_B2_  (\U_AHB/sel1_b17/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b17/or_B0_B1_o , \U_AHB/sel1_b1/B3 );
  or \U_AHB/sel1_b17/or_or_B4_B5_o_or_B6_  (\U_AHB/sel1_b17/or_or_B4_B5_o_or_B6__o , \U_AHB/sel1_b17/or_B4_B5_o , \U_AHB/sel1_b17/or_B6_or_B7_B8_o_o );
  or \U_AHB/sel1_b17/or_or_or_B0_B1_o_or_  (\U_AHB/n116 [17], \U_AHB/sel1_b17/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b17/or_or_B4_B5_o_or_B6__o );
  and \U_AHB/sel1_b18/and_b0_0  (\U_AHB/sel1_b18/B0 , \U_AHB/h2h_hrdata [18], \U_AHB/n104 );
  and \U_AHB/sel1_b18/and_b0_1  (\U_AHB/sel1_b18/B1 , limit_l[2], \U_AHB/n102 );
  and \U_AHB/sel1_b18/and_b0_3  (\U_AHB/sel1_b18/B3 , pwm_state_read[2], \U_AHB/n96 );
  and \U_AHB/sel1_b18/and_b0_4  (\U_AHB/sel1_b18/B4 , pnumcntF[18], \U_AHB/n93 );
  and \U_AHB/sel1_b18/and_b0_5  (\U_AHB/sel1_b18/B5 , pnumcntE[18], \U_AHB/n90 );
  and \U_AHB/sel1_b18/and_b0_6  (\U_AHB/sel1_b18/B6 , pnumcntD[18], \U_AHB/n87 );
  and \U_AHB/sel1_b18/and_b0_7  (\U_AHB/sel1_b18/B7 , pnumcntC[18], \U_AHB/n84 );
  and \U_AHB/sel1_b18/and_b0_8  (\U_AHB/sel1_b18/B8 , pnumcntB[18], \U_AHB/h2h_haddr [2]);
  or \U_AHB/sel1_b18/or_B0_B1  (\U_AHB/sel1_b18/or_B0_B1_o , \U_AHB/sel1_b18/B0 , \U_AHB/sel1_b18/B1 );
  or \U_AHB/sel1_b18/or_B4_B5  (\U_AHB/sel1_b18/or_B4_B5_o , \U_AHB/sel1_b18/B4 , \U_AHB/sel1_b18/B5 );
  or \U_AHB/sel1_b18/or_B6_or_B7_B8_o  (\U_AHB/sel1_b18/or_B6_or_B7_B8_o_o , \U_AHB/sel1_b18/B6 , \U_AHB/sel1_b18/or_B7_B8_o );
  or \U_AHB/sel1_b18/or_B7_B8  (\U_AHB/sel1_b18/or_B7_B8_o , \U_AHB/sel1_b18/B7 , \U_AHB/sel1_b18/B8 );
  or \U_AHB/sel1_b18/or_or_B0_B1_o_or_B2_  (\U_AHB/sel1_b18/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b18/or_B0_B1_o , \U_AHB/sel1_b18/B3 );
  or \U_AHB/sel1_b18/or_or_B4_B5_o_or_B6_  (\U_AHB/sel1_b18/or_or_B4_B5_o_or_B6__o , \U_AHB/sel1_b18/or_B4_B5_o , \U_AHB/sel1_b18/or_B6_or_B7_B8_o_o );
  or \U_AHB/sel1_b18/or_or_or_B0_B1_o_or_  (\U_AHB/n116 [18], \U_AHB/sel1_b18/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b18/or_or_B4_B5_o_or_B6__o );
  and \U_AHB/sel1_b19/and_b0_0  (\U_AHB/sel1_b19/B0 , \U_AHB/h2h_hrdata [19], \U_AHB/n104 );
  and \U_AHB/sel1_b19/and_b0_1  (\U_AHB/sel1_b19/B1 , limit_l[3], \U_AHB/n102 );
  and \U_AHB/sel1_b19/and_b0_3  (\U_AHB/sel1_b19/B3 , pwm_state_read[3], \U_AHB/n96 );
  and \U_AHB/sel1_b19/and_b0_4  (\U_AHB/sel1_b19/B4 , pnumcntF[19], \U_AHB/n93 );
  and \U_AHB/sel1_b19/and_b0_5  (\U_AHB/sel1_b19/B5 , pnumcntE[19], \U_AHB/n90 );
  and \U_AHB/sel1_b19/and_b0_6  (\U_AHB/sel1_b19/B6 , pnumcntD[19], \U_AHB/n87 );
  and \U_AHB/sel1_b19/and_b0_7  (\U_AHB/sel1_b19/B7 , pnumcntC[19], \U_AHB/n84 );
  and \U_AHB/sel1_b19/and_b0_8  (\U_AHB/sel1_b19/B8 , pnumcntB[19], \U_AHB/h2h_haddr [2]);
  or \U_AHB/sel1_b19/or_B0_B1  (\U_AHB/sel1_b19/or_B0_B1_o , \U_AHB/sel1_b19/B0 , \U_AHB/sel1_b19/B1 );
  or \U_AHB/sel1_b19/or_B4_B5  (\U_AHB/sel1_b19/or_B4_B5_o , \U_AHB/sel1_b19/B4 , \U_AHB/sel1_b19/B5 );
  or \U_AHB/sel1_b19/or_B6_or_B7_B8_o  (\U_AHB/sel1_b19/or_B6_or_B7_B8_o_o , \U_AHB/sel1_b19/B6 , \U_AHB/sel1_b19/or_B7_B8_o );
  or \U_AHB/sel1_b19/or_B7_B8  (\U_AHB/sel1_b19/or_B7_B8_o , \U_AHB/sel1_b19/B7 , \U_AHB/sel1_b19/B8 );
  or \U_AHB/sel1_b19/or_or_B0_B1_o_or_B2_  (\U_AHB/sel1_b19/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b19/or_B0_B1_o , \U_AHB/sel1_b19/B3 );
  or \U_AHB/sel1_b19/or_or_B4_B5_o_or_B6_  (\U_AHB/sel1_b19/or_or_B4_B5_o_or_B6__o , \U_AHB/sel1_b19/or_B4_B5_o , \U_AHB/sel1_b19/or_B6_or_B7_B8_o_o );
  or \U_AHB/sel1_b19/or_or_or_B0_B1_o_or_  (\U_AHB/n116 [19], \U_AHB/sel1_b19/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b19/or_or_B4_B5_o_or_B6__o );
  and \U_AHB/sel1_b2/and_b0_0  (\U_AHB/sel1_b2/B0 , \U_AHB/h2h_hrdata [2], \U_AHB/n104 );
  and \U_AHB/sel1_b2/and_b0_1  (\U_AHB/sel1_b2/B1 , limit_r[2], \U_AHB/n102 );
  and \U_AHB/sel1_b2/and_b0_4  (\U_AHB/sel1_b2/B4 , pnumcntF[2], \U_AHB/n93 );
  and \U_AHB/sel1_b2/and_b0_5  (\U_AHB/sel1_b2/B5 , pnumcntE[2], \U_AHB/n90 );
  and \U_AHB/sel1_b2/and_b0_6  (\U_AHB/sel1_b2/B6 , pnumcntD[2], \U_AHB/n87 );
  and \U_AHB/sel1_b2/and_b0_7  (\U_AHB/sel1_b2/B7 , pnumcntC[2], \U_AHB/n84 );
  and \U_AHB/sel1_b2/and_b0_8  (\U_AHB/sel1_b2/B8 , pnumcntB[2], \U_AHB/h2h_haddr [2]);
  or \U_AHB/sel1_b2/or_B0_B1  (\U_AHB/sel1_b2/or_B0_B1_o , \U_AHB/sel1_b2/B0 , \U_AHB/sel1_b2/B1 );
  or \U_AHB/sel1_b2/or_B4_B5  (\U_AHB/sel1_b2/or_B4_B5_o , \U_AHB/sel1_b2/B4 , \U_AHB/sel1_b2/B5 );
  or \U_AHB/sel1_b2/or_B6_or_B7_B8_o  (\U_AHB/sel1_b2/or_B6_or_B7_B8_o_o , \U_AHB/sel1_b2/B6 , \U_AHB/sel1_b2/or_B7_B8_o );
  or \U_AHB/sel1_b2/or_B7_B8  (\U_AHB/sel1_b2/or_B7_B8_o , \U_AHB/sel1_b2/B7 , \U_AHB/sel1_b2/B8 );
  or \U_AHB/sel1_b2/or_or_B0_B1_o_or_B2_  (\U_AHB/sel1_b2/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b2/or_B0_B1_o , \U_AHB/sel1_b18/B3 );
  or \U_AHB/sel1_b2/or_or_B4_B5_o_or_B6_  (\U_AHB/sel1_b2/or_or_B4_B5_o_or_B6__o , \U_AHB/sel1_b2/or_B4_B5_o , \U_AHB/sel1_b2/or_B6_or_B7_B8_o_o );
  or \U_AHB/sel1_b2/or_or_or_B0_B1_o_or_  (\U_AHB/n116 [2], \U_AHB/sel1_b2/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b2/or_or_B4_B5_o_or_B6__o );
  and \U_AHB/sel1_b20/and_b0_0  (\U_AHB/sel1_b20/B0 , \U_AHB/h2h_hrdata [20], \U_AHB/n104 );
  and \U_AHB/sel1_b20/and_b0_1  (\U_AHB/sel1_b20/B1 , limit_l[4], \U_AHB/n102 );
  and \U_AHB/sel1_b20/and_b0_3  (\U_AHB/sel1_b20/B3 , pwm_state_read[4], \U_AHB/n96 );
  and \U_AHB/sel1_b20/and_b0_4  (\U_AHB/sel1_b20/B4 , pnumcntF[20], \U_AHB/n93 );
  and \U_AHB/sel1_b20/and_b0_5  (\U_AHB/sel1_b20/B5 , pnumcntE[20], \U_AHB/n90 );
  and \U_AHB/sel1_b20/and_b0_6  (\U_AHB/sel1_b20/B6 , pnumcntD[20], \U_AHB/n87 );
  and \U_AHB/sel1_b20/and_b0_7  (\U_AHB/sel1_b20/B7 , pnumcntC[20], \U_AHB/n84 );
  and \U_AHB/sel1_b20/and_b0_8  (\U_AHB/sel1_b20/B8 , pnumcntB[20], \U_AHB/h2h_haddr [2]);
  or \U_AHB/sel1_b20/or_B0_B1  (\U_AHB/sel1_b20/or_B0_B1_o , \U_AHB/sel1_b20/B0 , \U_AHB/sel1_b20/B1 );
  or \U_AHB/sel1_b20/or_B4_B5  (\U_AHB/sel1_b20/or_B4_B5_o , \U_AHB/sel1_b20/B4 , \U_AHB/sel1_b20/B5 );
  or \U_AHB/sel1_b20/or_B6_or_B7_B8_o  (\U_AHB/sel1_b20/or_B6_or_B7_B8_o_o , \U_AHB/sel1_b20/B6 , \U_AHB/sel1_b20/or_B7_B8_o );
  or \U_AHB/sel1_b20/or_B7_B8  (\U_AHB/sel1_b20/or_B7_B8_o , \U_AHB/sel1_b20/B7 , \U_AHB/sel1_b20/B8 );
  or \U_AHB/sel1_b20/or_or_B0_B1_o_or_B2_  (\U_AHB/sel1_b20/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b20/or_B0_B1_o , \U_AHB/sel1_b20/B3 );
  or \U_AHB/sel1_b20/or_or_B4_B5_o_or_B6_  (\U_AHB/sel1_b20/or_or_B4_B5_o_or_B6__o , \U_AHB/sel1_b20/or_B4_B5_o , \U_AHB/sel1_b20/or_B6_or_B7_B8_o_o );
  or \U_AHB/sel1_b20/or_or_or_B0_B1_o_or_  (\U_AHB/n116 [20], \U_AHB/sel1_b20/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b20/or_or_B4_B5_o_or_B6__o );
  and \U_AHB/sel1_b21/and_b0_0  (\U_AHB/sel1_b21/B0 , \U_AHB/h2h_hrdata [21], \U_AHB/n104 );
  and \U_AHB/sel1_b21/and_b0_1  (\U_AHB/sel1_b21/B1 , limit_l[5], \U_AHB/n102 );
  and \U_AHB/sel1_b21/and_b0_3  (\U_AHB/sel1_b21/B3 , pwm_state_read[5], \U_AHB/n96 );
  and \U_AHB/sel1_b21/and_b0_4  (\U_AHB/sel1_b21/B4 , pnumcntF[21], \U_AHB/n93 );
  and \U_AHB/sel1_b21/and_b0_5  (\U_AHB/sel1_b21/B5 , pnumcntE[21], \U_AHB/n90 );
  and \U_AHB/sel1_b21/and_b0_6  (\U_AHB/sel1_b21/B6 , pnumcntD[21], \U_AHB/n87 );
  and \U_AHB/sel1_b21/and_b0_7  (\U_AHB/sel1_b21/B7 , pnumcntC[21], \U_AHB/n84 );
  and \U_AHB/sel1_b21/and_b0_8  (\U_AHB/sel1_b21/B8 , pnumcntB[21], \U_AHB/h2h_haddr [2]);
  or \U_AHB/sel1_b21/or_B0_B1  (\U_AHB/sel1_b21/or_B0_B1_o , \U_AHB/sel1_b21/B0 , \U_AHB/sel1_b21/B1 );
  or \U_AHB/sel1_b21/or_B4_B5  (\U_AHB/sel1_b21/or_B4_B5_o , \U_AHB/sel1_b21/B4 , \U_AHB/sel1_b21/B5 );
  or \U_AHB/sel1_b21/or_B6_or_B7_B8_o  (\U_AHB/sel1_b21/or_B6_or_B7_B8_o_o , \U_AHB/sel1_b21/B6 , \U_AHB/sel1_b21/or_B7_B8_o );
  or \U_AHB/sel1_b21/or_B7_B8  (\U_AHB/sel1_b21/or_B7_B8_o , \U_AHB/sel1_b21/B7 , \U_AHB/sel1_b21/B8 );
  or \U_AHB/sel1_b21/or_or_B0_B1_o_or_B2_  (\U_AHB/sel1_b21/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b21/or_B0_B1_o , \U_AHB/sel1_b21/B3 );
  or \U_AHB/sel1_b21/or_or_B4_B5_o_or_B6_  (\U_AHB/sel1_b21/or_or_B4_B5_o_or_B6__o , \U_AHB/sel1_b21/or_B4_B5_o , \U_AHB/sel1_b21/or_B6_or_B7_B8_o_o );
  or \U_AHB/sel1_b21/or_or_or_B0_B1_o_or_  (\U_AHB/n116 [21], \U_AHB/sel1_b21/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b21/or_or_B4_B5_o_or_B6__o );
  and \U_AHB/sel1_b22/and_b0_0  (\U_AHB/sel1_b22/B0 , \U_AHB/h2h_hrdata [22], \U_AHB/n104 );
  and \U_AHB/sel1_b22/and_b0_1  (\U_AHB/sel1_b22/B1 , limit_l[6], \U_AHB/n102 );
  and \U_AHB/sel1_b22/and_b0_3  (\U_AHB/sel1_b22/B3 , pwm_state_read[6], \U_AHB/n96 );
  and \U_AHB/sel1_b22/and_b0_4  (\U_AHB/sel1_b22/B4 , pnumcntF[22], \U_AHB/n93 );
  and \U_AHB/sel1_b22/and_b0_5  (\U_AHB/sel1_b22/B5 , pnumcntE[22], \U_AHB/n90 );
  and \U_AHB/sel1_b22/and_b0_6  (\U_AHB/sel1_b22/B6 , pnumcntD[22], \U_AHB/n87 );
  and \U_AHB/sel1_b22/and_b0_7  (\U_AHB/sel1_b22/B7 , pnumcntC[22], \U_AHB/n84 );
  and \U_AHB/sel1_b22/and_b0_8  (\U_AHB/sel1_b22/B8 , pnumcntB[22], \U_AHB/h2h_haddr [2]);
  or \U_AHB/sel1_b22/or_B0_B1  (\U_AHB/sel1_b22/or_B0_B1_o , \U_AHB/sel1_b22/B0 , \U_AHB/sel1_b22/B1 );
  or \U_AHB/sel1_b22/or_B4_B5  (\U_AHB/sel1_b22/or_B4_B5_o , \U_AHB/sel1_b22/B4 , \U_AHB/sel1_b22/B5 );
  or \U_AHB/sel1_b22/or_B6_or_B7_B8_o  (\U_AHB/sel1_b22/or_B6_or_B7_B8_o_o , \U_AHB/sel1_b22/B6 , \U_AHB/sel1_b22/or_B7_B8_o );
  or \U_AHB/sel1_b22/or_B7_B8  (\U_AHB/sel1_b22/or_B7_B8_o , \U_AHB/sel1_b22/B7 , \U_AHB/sel1_b22/B8 );
  or \U_AHB/sel1_b22/or_or_B0_B1_o_or_B2_  (\U_AHB/sel1_b22/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b22/or_B0_B1_o , \U_AHB/sel1_b22/B3 );
  or \U_AHB/sel1_b22/or_or_B4_B5_o_or_B6_  (\U_AHB/sel1_b22/or_or_B4_B5_o_or_B6__o , \U_AHB/sel1_b22/or_B4_B5_o , \U_AHB/sel1_b22/or_B6_or_B7_B8_o_o );
  or \U_AHB/sel1_b22/or_or_or_B0_B1_o_or_  (\U_AHB/n116 [22], \U_AHB/sel1_b22/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b22/or_or_B4_B5_o_or_B6__o );
  and \U_AHB/sel1_b23/and_b0_0  (\U_AHB/sel1_b23/B0 , \U_AHB/h2h_hrdata [23], \U_AHB/n104 );
  and \U_AHB/sel1_b23/and_b0_1  (\U_AHB/sel1_b23/B1 , limit_l[7], \U_AHB/n102 );
  and \U_AHB/sel1_b23/and_b0_3  (\U_AHB/sel1_b23/B3 , pwm_state_read[7], \U_AHB/n96 );
  and \U_AHB/sel1_b23/and_b0_4  (\U_AHB/sel1_b23/B4 , pnumcntF[23], \U_AHB/n93 );
  and \U_AHB/sel1_b23/and_b0_5  (\U_AHB/sel1_b23/B5 , pnumcntE[23], \U_AHB/n90 );
  and \U_AHB/sel1_b23/and_b0_6  (\U_AHB/sel1_b23/B6 , pnumcntD[23], \U_AHB/n87 );
  and \U_AHB/sel1_b23/and_b0_7  (\U_AHB/sel1_b23/B7 , pnumcntC[23], \U_AHB/n84 );
  and \U_AHB/sel1_b23/and_b0_8  (\U_AHB/sel1_b23/B8 , pnumcntB[23], \U_AHB/h2h_haddr [2]);
  or \U_AHB/sel1_b23/or_B0_B1  (\U_AHB/sel1_b23/or_B0_B1_o , \U_AHB/sel1_b23/B0 , \U_AHB/sel1_b23/B1 );
  or \U_AHB/sel1_b23/or_B4_B5  (\U_AHB/sel1_b23/or_B4_B5_o , \U_AHB/sel1_b23/B4 , \U_AHB/sel1_b23/B5 );
  or \U_AHB/sel1_b23/or_B6_or_B7_B8_o  (\U_AHB/sel1_b23/or_B6_or_B7_B8_o_o , \U_AHB/sel1_b23/B6 , \U_AHB/sel1_b23/or_B7_B8_o );
  or \U_AHB/sel1_b23/or_B7_B8  (\U_AHB/sel1_b23/or_B7_B8_o , \U_AHB/sel1_b23/B7 , \U_AHB/sel1_b23/B8 );
  or \U_AHB/sel1_b23/or_or_B0_B1_o_or_B2_  (\U_AHB/sel1_b23/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b23/or_B0_B1_o , \U_AHB/sel1_b23/B3 );
  or \U_AHB/sel1_b23/or_or_B4_B5_o_or_B6_  (\U_AHB/sel1_b23/or_or_B4_B5_o_or_B6__o , \U_AHB/sel1_b23/or_B4_B5_o , \U_AHB/sel1_b23/or_B6_or_B7_B8_o_o );
  or \U_AHB/sel1_b23/or_or_or_B0_B1_o_or_  (\U_AHB/n116 [23], \U_AHB/sel1_b23/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b23/or_or_B4_B5_o_or_B6__o );
  and \U_AHB/sel1_b24/and_b0_0  (\U_AHB/sel1_b24/B0 , \U_AHB/h2h_hrdata [24], \U_AHB/n104 );
  and \U_AHB/sel1_b24/and_b0_1  (\U_AHB/sel1_b24/B1 , limit_l[8], \U_AHB/n102 );
  and \U_AHB/sel1_b24/and_b0_3  (\U_AHB/sel1_b24/B3 , pwm_state_read[8], \U_AHB/n96 );
  or \U_AHB/sel1_b24/or_B0_B1  (\U_AHB/sel1_b24/or_B0_B1_o , \U_AHB/sel1_b24/B0 , \U_AHB/sel1_b24/B1 );
  or \U_AHB/sel1_b24/or_or_B0_B1_o_or_B2_  (\U_AHB/sel1_b24/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b24/or_B0_B1_o , \U_AHB/sel1_b24/B3 );
  and \U_AHB/sel1_b25/and_b0_0  (\U_AHB/sel1_b25/B0 , \U_AHB/h2h_hrdata [25], \U_AHB/n104 );
  and \U_AHB/sel1_b25/and_b0_1  (\U_AHB/sel1_b25/B1 , limit_l[9], \U_AHB/n102 );
  and \U_AHB/sel1_b25/and_b0_3  (\U_AHB/sel1_b25/B3 , pwm_state_read[9], \U_AHB/n96 );
  or \U_AHB/sel1_b25/or_B0_B1  (\U_AHB/sel1_b25/or_B0_B1_o , \U_AHB/sel1_b25/B0 , \U_AHB/sel1_b25/B1 );
  or \U_AHB/sel1_b25/or_or_B0_B1_o_or_B2_  (\U_AHB/sel1_b25/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b25/or_B0_B1_o , \U_AHB/sel1_b25/B3 );
  and \U_AHB/sel1_b26/and_b0_0  (\U_AHB/sel1_b26/B0 , \U_AHB/h2h_hrdata [26], \U_AHB/n104 );
  and \U_AHB/sel1_b26/and_b0_1  (\U_AHB/sel1_b26/B1 , limit_l[10], \U_AHB/n102 );
  or \U_AHB/sel1_b26/or_B0_B1  (\U_AHB/sel1_b26/or_B0_B1_o , \U_AHB/sel1_b26/B0 , \U_AHB/sel1_b26/B1 );
  or \U_AHB/sel1_b26/or_or_B0_B1_o_or_B2_  (\U_AHB/sel1_b26/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b26/or_B0_B1_o , \U_AHB/sel1_b10/B3 );
  and \U_AHB/sel1_b27/and_b0_0  (\U_AHB/sel1_b27/B0 , \U_AHB/h2h_hrdata [27], \U_AHB/n104 );
  and \U_AHB/sel1_b27/and_b0_1  (\U_AHB/sel1_b27/B1 , limit_l[11], \U_AHB/n102 );
  or \U_AHB/sel1_b27/or_B0_B1  (\U_AHB/sel1_b27/or_B0_B1_o , \U_AHB/sel1_b27/B0 , \U_AHB/sel1_b27/B1 );
  or \U_AHB/sel1_b27/or_or_B0_B1_o_or_B2_  (\U_AHB/sel1_b27/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b27/or_B0_B1_o , \U_AHB/sel1_b11/B3 );
  and \U_AHB/sel1_b28/and_b0_0  (\U_AHB/sel1_b28/B0 , \U_AHB/h2h_hrdata [28], \U_AHB/n104 );
  and \U_AHB/sel1_b28/and_b0_1  (\U_AHB/sel1_b28/B1 , limit_l[12], \U_AHB/n102 );
  or \U_AHB/sel1_b28/or_B0_B1  (\U_AHB/sel1_b28/or_B0_B1_o , \U_AHB/sel1_b28/B0 , \U_AHB/sel1_b28/B1 );
  or \U_AHB/sel1_b28/or_or_B0_B1_o_or_B2_  (\U_AHB/sel1_b28/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b28/or_B0_B1_o , \U_AHB/sel1_b12/B3 );
  and \U_AHB/sel1_b29/and_b0_0  (\U_AHB/sel1_b29/B0 , \U_AHB/h2h_hrdata [29], \U_AHB/n104 );
  and \U_AHB/sel1_b29/and_b0_1  (\U_AHB/sel1_b29/B1 , limit_l[13], \U_AHB/n102 );
  or \U_AHB/sel1_b29/or_B0_B1  (\U_AHB/sel1_b29/or_B0_B1_o , \U_AHB/sel1_b29/B0 , \U_AHB/sel1_b29/B1 );
  or \U_AHB/sel1_b29/or_or_B0_B1_o_or_B2_  (\U_AHB/sel1_b29/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b29/or_B0_B1_o , \U_AHB/sel1_b13/B3 );
  and \U_AHB/sel1_b3/and_b0_0  (\U_AHB/sel1_b3/B0 , \U_AHB/h2h_hrdata [3], \U_AHB/n104 );
  and \U_AHB/sel1_b3/and_b0_1  (\U_AHB/sel1_b3/B1 , limit_r[3], \U_AHB/n102 );
  and \U_AHB/sel1_b3/and_b0_4  (\U_AHB/sel1_b3/B4 , pnumcntF[3], \U_AHB/n93 );
  and \U_AHB/sel1_b3/and_b0_5  (\U_AHB/sel1_b3/B5 , pnumcntE[3], \U_AHB/n90 );
  and \U_AHB/sel1_b3/and_b0_6  (\U_AHB/sel1_b3/B6 , pnumcntD[3], \U_AHB/n87 );
  and \U_AHB/sel1_b3/and_b0_7  (\U_AHB/sel1_b3/B7 , pnumcntC[3], \U_AHB/n84 );
  and \U_AHB/sel1_b3/and_b0_8  (\U_AHB/sel1_b3/B8 , pnumcntB[3], \U_AHB/h2h_haddr [2]);
  or \U_AHB/sel1_b3/or_B0_B1  (\U_AHB/sel1_b3/or_B0_B1_o , \U_AHB/sel1_b3/B0 , \U_AHB/sel1_b3/B1 );
  or \U_AHB/sel1_b3/or_B4_B5  (\U_AHB/sel1_b3/or_B4_B5_o , \U_AHB/sel1_b3/B4 , \U_AHB/sel1_b3/B5 );
  or \U_AHB/sel1_b3/or_B6_or_B7_B8_o  (\U_AHB/sel1_b3/or_B6_or_B7_B8_o_o , \U_AHB/sel1_b3/B6 , \U_AHB/sel1_b3/or_B7_B8_o );
  or \U_AHB/sel1_b3/or_B7_B8  (\U_AHB/sel1_b3/or_B7_B8_o , \U_AHB/sel1_b3/B7 , \U_AHB/sel1_b3/B8 );
  or \U_AHB/sel1_b3/or_or_B0_B1_o_or_B2_  (\U_AHB/sel1_b3/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b3/or_B0_B1_o , \U_AHB/sel1_b19/B3 );
  or \U_AHB/sel1_b3/or_or_B4_B5_o_or_B6_  (\U_AHB/sel1_b3/or_or_B4_B5_o_or_B6__o , \U_AHB/sel1_b3/or_B4_B5_o , \U_AHB/sel1_b3/or_B6_or_B7_B8_o_o );
  or \U_AHB/sel1_b3/or_or_or_B0_B1_o_or_  (\U_AHB/n116 [3], \U_AHB/sel1_b3/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b3/or_or_B4_B5_o_or_B6__o );
  and \U_AHB/sel1_b30/and_b0_0  (\U_AHB/sel1_b30/B0 , \U_AHB/h2h_hrdata [30], \U_AHB/n104 );
  and \U_AHB/sel1_b30/and_b0_1  (\U_AHB/sel1_b30/B1 , limit_l[14], \U_AHB/n102 );
  or \U_AHB/sel1_b30/or_B0_B1  (\U_AHB/sel1_b30/or_B0_B1_o , \U_AHB/sel1_b30/B0 , \U_AHB/sel1_b30/B1 );
  or \U_AHB/sel1_b30/or_or_B0_B1_o_or_B2_  (\U_AHB/sel1_b30/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b30/or_B0_B1_o , \U_AHB/sel1_b14/B3 );
  and \U_AHB/sel1_b31/and_b0_0  (\U_AHB/sel1_b31/B0 , \U_AHB/h2h_hrdata [31], \U_AHB/n104 );
  and \U_AHB/sel1_b31/and_b0_1  (\U_AHB/sel1_b31/B1 , limit_l[15], \U_AHB/n102 );
  or \U_AHB/sel1_b31/or_B0_B1  (\U_AHB/sel1_b31/or_B0_B1_o , \U_AHB/sel1_b31/B0 , \U_AHB/sel1_b31/B1 );
  or \U_AHB/sel1_b31/or_or_B0_B1_o_or_B2_  (\U_AHB/sel1_b31/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b31/or_B0_B1_o , \U_AHB/sel1_b15/B3 );
  and \U_AHB/sel1_b4/and_b0_0  (\U_AHB/sel1_b4/B0 , \U_AHB/h2h_hrdata [4], \U_AHB/n104 );
  and \U_AHB/sel1_b4/and_b0_1  (\U_AHB/sel1_b4/B1 , limit_r[4], \U_AHB/n102 );
  and \U_AHB/sel1_b4/and_b0_4  (\U_AHB/sel1_b4/B4 , pnumcntF[4], \U_AHB/n93 );
  and \U_AHB/sel1_b4/and_b0_5  (\U_AHB/sel1_b4/B5 , pnumcntE[4], \U_AHB/n90 );
  and \U_AHB/sel1_b4/and_b0_6  (\U_AHB/sel1_b4/B6 , pnumcntD[4], \U_AHB/n87 );
  and \U_AHB/sel1_b4/and_b0_7  (\U_AHB/sel1_b4/B7 , pnumcntC[4], \U_AHB/n84 );
  and \U_AHB/sel1_b4/and_b0_8  (\U_AHB/sel1_b4/B8 , pnumcntB[4], \U_AHB/h2h_haddr [2]);
  or \U_AHB/sel1_b4/or_B0_B1  (\U_AHB/sel1_b4/or_B0_B1_o , \U_AHB/sel1_b4/B0 , \U_AHB/sel1_b4/B1 );
  or \U_AHB/sel1_b4/or_B4_B5  (\U_AHB/sel1_b4/or_B4_B5_o , \U_AHB/sel1_b4/B4 , \U_AHB/sel1_b4/B5 );
  or \U_AHB/sel1_b4/or_B6_or_B7_B8_o  (\U_AHB/sel1_b4/or_B6_or_B7_B8_o_o , \U_AHB/sel1_b4/B6 , \U_AHB/sel1_b4/or_B7_B8_o );
  or \U_AHB/sel1_b4/or_B7_B8  (\U_AHB/sel1_b4/or_B7_B8_o , \U_AHB/sel1_b4/B7 , \U_AHB/sel1_b4/B8 );
  or \U_AHB/sel1_b4/or_or_B0_B1_o_or_B2_  (\U_AHB/sel1_b4/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b4/or_B0_B1_o , \U_AHB/sel1_b20/B3 );
  or \U_AHB/sel1_b4/or_or_B4_B5_o_or_B6_  (\U_AHB/sel1_b4/or_or_B4_B5_o_or_B6__o , \U_AHB/sel1_b4/or_B4_B5_o , \U_AHB/sel1_b4/or_B6_or_B7_B8_o_o );
  or \U_AHB/sel1_b4/or_or_or_B0_B1_o_or_  (\U_AHB/n116 [4], \U_AHB/sel1_b4/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b4/or_or_B4_B5_o_or_B6__o );
  and \U_AHB/sel1_b5/and_b0_0  (\U_AHB/sel1_b5/B0 , \U_AHB/h2h_hrdata [5], \U_AHB/n104 );
  and \U_AHB/sel1_b5/and_b0_1  (\U_AHB/sel1_b5/B1 , limit_r[5], \U_AHB/n102 );
  and \U_AHB/sel1_b5/and_b0_4  (\U_AHB/sel1_b5/B4 , pnumcntF[5], \U_AHB/n93 );
  and \U_AHB/sel1_b5/and_b0_5  (\U_AHB/sel1_b5/B5 , pnumcntE[5], \U_AHB/n90 );
  and \U_AHB/sel1_b5/and_b0_6  (\U_AHB/sel1_b5/B6 , pnumcntD[5], \U_AHB/n87 );
  and \U_AHB/sel1_b5/and_b0_7  (\U_AHB/sel1_b5/B7 , pnumcntC[5], \U_AHB/n84 );
  and \U_AHB/sel1_b5/and_b0_8  (\U_AHB/sel1_b5/B8 , pnumcntB[5], \U_AHB/h2h_haddr [2]);
  or \U_AHB/sel1_b5/or_B0_B1  (\U_AHB/sel1_b5/or_B0_B1_o , \U_AHB/sel1_b5/B0 , \U_AHB/sel1_b5/B1 );
  or \U_AHB/sel1_b5/or_B4_B5  (\U_AHB/sel1_b5/or_B4_B5_o , \U_AHB/sel1_b5/B4 , \U_AHB/sel1_b5/B5 );
  or \U_AHB/sel1_b5/or_B6_or_B7_B8_o  (\U_AHB/sel1_b5/or_B6_or_B7_B8_o_o , \U_AHB/sel1_b5/B6 , \U_AHB/sel1_b5/or_B7_B8_o );
  or \U_AHB/sel1_b5/or_B7_B8  (\U_AHB/sel1_b5/or_B7_B8_o , \U_AHB/sel1_b5/B7 , \U_AHB/sel1_b5/B8 );
  or \U_AHB/sel1_b5/or_or_B0_B1_o_or_B2_  (\U_AHB/sel1_b5/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b5/or_B0_B1_o , \U_AHB/sel1_b21/B3 );
  or \U_AHB/sel1_b5/or_or_B4_B5_o_or_B6_  (\U_AHB/sel1_b5/or_or_B4_B5_o_or_B6__o , \U_AHB/sel1_b5/or_B4_B5_o , \U_AHB/sel1_b5/or_B6_or_B7_B8_o_o );
  or \U_AHB/sel1_b5/or_or_or_B0_B1_o_or_  (\U_AHB/n116 [5], \U_AHB/sel1_b5/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b5/or_or_B4_B5_o_or_B6__o );
  and \U_AHB/sel1_b6/and_b0_0  (\U_AHB/sel1_b6/B0 , \U_AHB/h2h_hrdata [6], \U_AHB/n104 );
  and \U_AHB/sel1_b6/and_b0_1  (\U_AHB/sel1_b6/B1 , limit_r[6], \U_AHB/n102 );
  and \U_AHB/sel1_b6/and_b0_4  (\U_AHB/sel1_b6/B4 , pnumcntF[6], \U_AHB/n93 );
  and \U_AHB/sel1_b6/and_b0_5  (\U_AHB/sel1_b6/B5 , pnumcntE[6], \U_AHB/n90 );
  and \U_AHB/sel1_b6/and_b0_6  (\U_AHB/sel1_b6/B6 , pnumcntD[6], \U_AHB/n87 );
  and \U_AHB/sel1_b6/and_b0_7  (\U_AHB/sel1_b6/B7 , pnumcntC[6], \U_AHB/n84 );
  and \U_AHB/sel1_b6/and_b0_8  (\U_AHB/sel1_b6/B8 , pnumcntB[6], \U_AHB/h2h_haddr [2]);
  or \U_AHB/sel1_b6/or_B0_B1  (\U_AHB/sel1_b6/or_B0_B1_o , \U_AHB/sel1_b6/B0 , \U_AHB/sel1_b6/B1 );
  or \U_AHB/sel1_b6/or_B4_B5  (\U_AHB/sel1_b6/or_B4_B5_o , \U_AHB/sel1_b6/B4 , \U_AHB/sel1_b6/B5 );
  or \U_AHB/sel1_b6/or_B6_or_B7_B8_o  (\U_AHB/sel1_b6/or_B6_or_B7_B8_o_o , \U_AHB/sel1_b6/B6 , \U_AHB/sel1_b6/or_B7_B8_o );
  or \U_AHB/sel1_b6/or_B7_B8  (\U_AHB/sel1_b6/or_B7_B8_o , \U_AHB/sel1_b6/B7 , \U_AHB/sel1_b6/B8 );
  or \U_AHB/sel1_b6/or_or_B0_B1_o_or_B2_  (\U_AHB/sel1_b6/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b6/or_B0_B1_o , \U_AHB/sel1_b22/B3 );
  or \U_AHB/sel1_b6/or_or_B4_B5_o_or_B6_  (\U_AHB/sel1_b6/or_or_B4_B5_o_or_B6__o , \U_AHB/sel1_b6/or_B4_B5_o , \U_AHB/sel1_b6/or_B6_or_B7_B8_o_o );
  or \U_AHB/sel1_b6/or_or_or_B0_B1_o_or_  (\U_AHB/n116 [6], \U_AHB/sel1_b6/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b6/or_or_B4_B5_o_or_B6__o );
  and \U_AHB/sel1_b7/and_b0_0  (\U_AHB/sel1_b7/B0 , \U_AHB/h2h_hrdata [7], \U_AHB/n104 );
  and \U_AHB/sel1_b7/and_b0_1  (\U_AHB/sel1_b7/B1 , limit_r[7], \U_AHB/n102 );
  and \U_AHB/sel1_b7/and_b0_4  (\U_AHB/sel1_b7/B4 , pnumcntF[7], \U_AHB/n93 );
  and \U_AHB/sel1_b7/and_b0_5  (\U_AHB/sel1_b7/B5 , pnumcntE[7], \U_AHB/n90 );
  and \U_AHB/sel1_b7/and_b0_6  (\U_AHB/sel1_b7/B6 , pnumcntD[7], \U_AHB/n87 );
  and \U_AHB/sel1_b7/and_b0_7  (\U_AHB/sel1_b7/B7 , pnumcntC[7], \U_AHB/n84 );
  and \U_AHB/sel1_b7/and_b0_8  (\U_AHB/sel1_b7/B8 , pnumcntB[7], \U_AHB/h2h_haddr [2]);
  or \U_AHB/sel1_b7/or_B0_B1  (\U_AHB/sel1_b7/or_B0_B1_o , \U_AHB/sel1_b7/B0 , \U_AHB/sel1_b7/B1 );
  or \U_AHB/sel1_b7/or_B4_B5  (\U_AHB/sel1_b7/or_B4_B5_o , \U_AHB/sel1_b7/B4 , \U_AHB/sel1_b7/B5 );
  or \U_AHB/sel1_b7/or_B6_or_B7_B8_o  (\U_AHB/sel1_b7/or_B6_or_B7_B8_o_o , \U_AHB/sel1_b7/B6 , \U_AHB/sel1_b7/or_B7_B8_o );
  or \U_AHB/sel1_b7/or_B7_B8  (\U_AHB/sel1_b7/or_B7_B8_o , \U_AHB/sel1_b7/B7 , \U_AHB/sel1_b7/B8 );
  or \U_AHB/sel1_b7/or_or_B0_B1_o_or_B2_  (\U_AHB/sel1_b7/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b7/or_B0_B1_o , \U_AHB/sel1_b23/B3 );
  or \U_AHB/sel1_b7/or_or_B4_B5_o_or_B6_  (\U_AHB/sel1_b7/or_or_B4_B5_o_or_B6__o , \U_AHB/sel1_b7/or_B4_B5_o , \U_AHB/sel1_b7/or_B6_or_B7_B8_o_o );
  or \U_AHB/sel1_b7/or_or_or_B0_B1_o_or_  (\U_AHB/n116 [7], \U_AHB/sel1_b7/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b7/or_or_B4_B5_o_or_B6__o );
  and \U_AHB/sel1_b8/and_b0_0  (\U_AHB/sel1_b8/B0 , \U_AHB/h2h_hrdata [8], \U_AHB/n104 );
  and \U_AHB/sel1_b8/and_b0_1  (\U_AHB/sel1_b8/B1 , limit_r[8], \U_AHB/n102 );
  and \U_AHB/sel1_b8/and_b0_4  (\U_AHB/sel1_b8/B4 , pnumcntF[8], \U_AHB/n93 );
  and \U_AHB/sel1_b8/and_b0_5  (\U_AHB/sel1_b8/B5 , pnumcntE[8], \U_AHB/n90 );
  and \U_AHB/sel1_b8/and_b0_6  (\U_AHB/sel1_b8/B6 , pnumcntD[8], \U_AHB/n87 );
  and \U_AHB/sel1_b8/and_b0_7  (\U_AHB/sel1_b8/B7 , pnumcntC[8], \U_AHB/n84 );
  and \U_AHB/sel1_b8/and_b0_8  (\U_AHB/sel1_b8/B8 , pnumcntB[8], \U_AHB/h2h_haddr [2]);
  or \U_AHB/sel1_b8/or_B0_B1  (\U_AHB/sel1_b8/or_B0_B1_o , \U_AHB/sel1_b8/B0 , \U_AHB/sel1_b8/B1 );
  or \U_AHB/sel1_b8/or_B4_B5  (\U_AHB/sel1_b8/or_B4_B5_o , \U_AHB/sel1_b8/B4 , \U_AHB/sel1_b8/B5 );
  or \U_AHB/sel1_b8/or_B6_or_B7_B8_o  (\U_AHB/sel1_b8/or_B6_or_B7_B8_o_o , \U_AHB/sel1_b8/B6 , \U_AHB/sel1_b8/or_B7_B8_o );
  or \U_AHB/sel1_b8/or_B7_B8  (\U_AHB/sel1_b8/or_B7_B8_o , \U_AHB/sel1_b8/B7 , \U_AHB/sel1_b8/B8 );
  or \U_AHB/sel1_b8/or_or_B0_B1_o_or_B2_  (\U_AHB/sel1_b8/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b8/or_B0_B1_o , \U_AHB/sel1_b24/B3 );
  or \U_AHB/sel1_b8/or_or_B4_B5_o_or_B6_  (\U_AHB/sel1_b8/or_or_B4_B5_o_or_B6__o , \U_AHB/sel1_b8/or_B4_B5_o , \U_AHB/sel1_b8/or_B6_or_B7_B8_o_o );
  or \U_AHB/sel1_b8/or_or_or_B0_B1_o_or_  (\U_AHB/n116 [8], \U_AHB/sel1_b8/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b8/or_or_B4_B5_o_or_B6__o );
  and \U_AHB/sel1_b9/and_b0_0  (\U_AHB/sel1_b9/B0 , \U_AHB/h2h_hrdata [9], \U_AHB/n104 );
  and \U_AHB/sel1_b9/and_b0_1  (\U_AHB/sel1_b9/B1 , limit_r[9], \U_AHB/n102 );
  and \U_AHB/sel1_b9/and_b0_4  (\U_AHB/sel1_b9/B4 , pnumcntF[9], \U_AHB/n93 );
  and \U_AHB/sel1_b9/and_b0_5  (\U_AHB/sel1_b9/B5 , pnumcntE[9], \U_AHB/n90 );
  and \U_AHB/sel1_b9/and_b0_6  (\U_AHB/sel1_b9/B6 , pnumcntD[9], \U_AHB/n87 );
  and \U_AHB/sel1_b9/and_b0_7  (\U_AHB/sel1_b9/B7 , pnumcntC[9], \U_AHB/n84 );
  and \U_AHB/sel1_b9/and_b0_8  (\U_AHB/sel1_b9/B8 , pnumcntB[9], \U_AHB/h2h_haddr [2]);
  or \U_AHB/sel1_b9/or_B0_B1  (\U_AHB/sel1_b9/or_B0_B1_o , \U_AHB/sel1_b9/B0 , \U_AHB/sel1_b9/B1 );
  or \U_AHB/sel1_b9/or_B4_B5  (\U_AHB/sel1_b9/or_B4_B5_o , \U_AHB/sel1_b9/B4 , \U_AHB/sel1_b9/B5 );
  or \U_AHB/sel1_b9/or_B6_or_B7_B8_o  (\U_AHB/sel1_b9/or_B6_or_B7_B8_o_o , \U_AHB/sel1_b9/B6 , \U_AHB/sel1_b9/or_B7_B8_o );
  or \U_AHB/sel1_b9/or_B7_B8  (\U_AHB/sel1_b9/or_B7_B8_o , \U_AHB/sel1_b9/B7 , \U_AHB/sel1_b9/B8 );
  or \U_AHB/sel1_b9/or_or_B0_B1_o_or_B2_  (\U_AHB/sel1_b9/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b9/or_B0_B1_o , \U_AHB/sel1_b25/B3 );
  or \U_AHB/sel1_b9/or_or_B4_B5_o_or_B6_  (\U_AHB/sel1_b9/or_or_B4_B5_o_or_B6__o , \U_AHB/sel1_b9/or_B4_B5_o , \U_AHB/sel1_b9/or_B6_or_B7_B8_o_o );
  or \U_AHB/sel1_b9/or_or_or_B0_B1_o_or_  (\U_AHB/n116 [9], \U_AHB/sel1_b9/or_or_B0_B1_o_or_B2__o , \U_AHB/sel1_b9/or_or_B4_B5_o_or_B6__o );
  or \U_AHB/u10  (\U_AHB/n37 [21], gpio_out[21], \U_AHB/h2h_hwdata [21]);  // src/AHB.v(63)
  and \U_AHB/u100  (\U_AHB/n40 [27], gpio_out[27], \U_AHB/n39 [27]);  // src/AHB.v(64)
  and \U_AHB/u101  (\U_AHB/n77 , \U_AHB/n44 , \U_AHB/h2h_haddr [4]);  // src/AHB.v(82)
  and \U_AHB/u102  (\U_AHB/n40 [26], gpio_out[26], \U_AHB/n39 [26]);  // src/AHB.v(64)
  and \U_AHB/u103  (\U_AHB/n40 [25], gpio_out[25], \U_AHB/n39 [25]);  // src/AHB.v(64)
  and \U_AHB/u104  (\U_AHB/n79 , \U_AHB/n44 , \U_AHB/h2h_haddr [7]);  // src/AHB.v(83)
  not \U_AHB/u105  (\U_AHB/n81 , \U_AHB/h2h_hwrite );  // src/AHB.v(88)
  and \U_AHB/u106  (\U_AHB/n40 [24], gpio_out[24], \U_AHB/n39 [24]);  // src/AHB.v(64)
  and \U_AHB/u107  (\U_AHB/n82 , \U_AHB/n81 , \U_AHB/n6 );  // src/AHB.v(88)
  not \U_AHB/u108  (\U_AHB/n83 , \U_AHB/h2h_haddr [2]);  // src/AHB.v(101)
  and \U_AHB/u109  (\U_AHB/n84 , \U_AHB/h2h_haddr [3], \U_AHB/n83 );  // src/AHB.v(101)
  and \U_AHB/u11  (\U_AHB/n10 , \U_AHB/n7 , \U_AHB/h2h_haddr [3]);  // src/AHB.v(49)
  or \U_AHB/u110  (\U_AHB/n85 , \U_AHB/h2h_haddr [2], \U_AHB/h2h_haddr [3]);  // src/AHB.v(101)
  not \U_AHB/u111  (\U_AHB/n86 , \U_AHB/n85 );  // src/AHB.v(101)
  and \U_AHB/u112  (\U_AHB/n87 , \U_AHB/h2h_haddr [4], \U_AHB/n86 );  // src/AHB.v(101)
  or \U_AHB/u113  (\U_AHB/n88 , \U_AHB/n85 , \U_AHB/h2h_haddr [4]);  // src/AHB.v(101)
  not \U_AHB/u114  (\U_AHB/n89 , \U_AHB/n88 );  // src/AHB.v(101)
  and \U_AHB/u115  (\U_AHB/n90 , \U_AHB/h2h_haddr [5], \U_AHB/n89 );  // src/AHB.v(101)
  or \U_AHB/u116  (\U_AHB/n91 , \U_AHB/n88 , \U_AHB/h2h_haddr [5]);  // src/AHB.v(101)
  not \U_AHB/u117  (\U_AHB/n92 , \U_AHB/n91 );  // src/AHB.v(101)
  and \U_AHB/u118  (\U_AHB/n93 , \U_AHB/h2h_haddr [6], \U_AHB/n92 );  // src/AHB.v(101)
  or \U_AHB/u119  (\U_AHB/n94 , \U_AHB/n91 , \U_AHB/h2h_haddr [6]);  // src/AHB.v(101)
  or \U_AHB/u12  (\U_AHB/n37 [20], gpio_out[20], \U_AHB/h2h_hwdata [20]);  // src/AHB.v(63)
  not \U_AHB/u120  (\U_AHB/n95 , \U_AHB/n94 );  // src/AHB.v(101)
  and \U_AHB/u121  (\U_AHB/n96 , \U_AHB/h2h_haddr [7], \U_AHB/n95 );  // src/AHB.v(101)
  or \U_AHB/u122  (\U_AHB/n97 , \U_AHB/n94 , \U_AHB/h2h_haddr [7]);  // src/AHB.v(101)
  not \U_AHB/u123  (\U_AHB/n98 , \U_AHB/n97 );  // src/AHB.v(101)
  and \U_AHB/u124  (\U_AHB/n99 , \U_AHB/h2h_haddr [8], \U_AHB/n98 );  // src/AHB.v(101)
  or \U_AHB/u125  (\U_AHB/n100 , \U_AHB/n97 , \U_AHB/h2h_haddr [8]);  // src/AHB.v(101)
  not \U_AHB/u126  (\U_AHB/n101 , \U_AHB/n100 );  // src/AHB.v(101)
  and \U_AHB/u127  (\U_AHB/n102 , \U_AHB/h2h_haddr [9], \U_AHB/n101 );  // src/AHB.v(101)
  or \U_AHB/u128  (\U_AHB/n103 , \U_AHB/n100 , \U_AHB/h2h_haddr [9]);  // src/AHB.v(101)
  not \U_AHB/u129  (\U_AHB/n104 , \U_AHB/n103 );  // src/AHB.v(101)
  or \U_AHB/u13  (\U_AHB/n37 [19], gpio_out[19], \U_AHB/h2h_hwdata [19]);  // src/AHB.v(63)
  and \U_AHB/u130  (\U_AHB/n105 , \U_AHB/h2h_haddr [10], \U_AHB/n104 );  // src/AHB.v(101)
  or \U_AHB/u131  (\U_AHB/n106 , \U_AHB/n103 , \U_AHB/h2h_haddr [10]);  // src/AHB.v(101)
  not \U_AHB/u132  (\U_AHB/n107 , \U_AHB/n106 );  // src/AHB.v(101)
  and \U_AHB/u133  (\U_AHB/n108 , \U_AHB/h2h_haddr [11], \U_AHB/n107 );  // src/AHB.v(101)
  or \U_AHB/u134  (\U_AHB/n109 , \U_AHB/n106 , \U_AHB/h2h_haddr [11]);  // src/AHB.v(101)
  not \U_AHB/u135  (\U_AHB/n110 , \U_AHB/n109 );  // src/AHB.v(101)
  and \U_AHB/u136  (\U_AHB/n111 , \U_AHB/h2h_haddr [12], \U_AHB/n110 );  // src/AHB.v(101)
  or \U_AHB/u137  (\U_AHB/n112 , \U_AHB/n109 , \U_AHB/h2h_haddr [12]);  // src/AHB.v(101)
  not \U_AHB/u138  (\U_AHB/n113 , \U_AHB/n112 );  // src/AHB.v(101)
  and \U_AHB/u139  (\U_AHB/n40 [23], gpio_out[23], \U_AHB/n39 [23]);  // src/AHB.v(64)
  and \U_AHB/u14  (\U_AHB/n12 , \U_AHB/n7 , \U_AHB/h2h_haddr [4]);  // src/AHB.v(50)
  and \U_AHB/u140  (\U_AHB/n40 [22], gpio_out[22], \U_AHB/n39 [22]);  // src/AHB.v(64)
  and \U_AHB/u141  (\U_AHB/n115 , \U_AHB/n81 , \U_AHB/n0 );  // src/AHB.v(103)
  or \U_AHB/u142  (\U_AHB/n37 [31], gpio_out[31], \U_AHB/h2h_hwdata [31]);  // src/AHB.v(63)
  or \U_AHB/u143  (\U_AHB/n37 [30], gpio_out[30], \U_AHB/h2h_hwdata [30]);  // src/AHB.v(63)
  or \U_AHB/u144  (\U_AHB/n37 [29], gpio_out[29], \U_AHB/h2h_hwdata [29]);  // src/AHB.v(63)
  or \U_AHB/u145  (\U_AHB/n37 [28], gpio_out[28], \U_AHB/h2h_hwdata [28]);  // src/AHB.v(63)
  or \U_AHB/u146  (\U_AHB/n37 [27], gpio_out[27], \U_AHB/h2h_hwdata [27]);  // src/AHB.v(63)
  or \U_AHB/u147  (\U_AHB/n37 [26], gpio_out[26], \U_AHB/h2h_hwdata [26]);  // src/AHB.v(63)
  or \U_AHB/u148  (\U_AHB/n37 [25], gpio_out[25], \U_AHB/h2h_hwdata [25]);  // src/AHB.v(63)
  and \U_AHB/u149  (\U_AHB/n40 [21], gpio_out[21], \U_AHB/n39 [21]);  // src/AHB.v(64)
  or \U_AHB/u15  (\U_AHB/n37 [18], gpio_out[18], \U_AHB/h2h_hwdata [18]);  // src/AHB.v(63)
  and \U_AHB/u150  (\U_AHB/n40 [20], gpio_out[20], \U_AHB/n39 [20]);  // src/AHB.v(64)
  and \U_AHB/u151  (\U_AHB/n40 [19], gpio_out[19], \U_AHB/n39 [19]);  // src/AHB.v(64)
  and \U_AHB/u152  (\U_AHB/n40 [18], gpio_out[18], \U_AHB/n39 [18]);  // src/AHB.v(64)
  and \U_AHB/u153  (\U_AHB/n40 [17], gpio_out[17], \U_AHB/n39 [17]);  // src/AHB.v(64)
  and \U_AHB/u154  (\U_AHB/n40 [16], gpio_out[16], \U_AHB/n39 [16]);  // src/AHB.v(64)
  and \U_AHB/u155  (\U_AHB/n40 [15], gpio_out[15], \U_AHB/n39 [15]);  // src/AHB.v(64)
  and \U_AHB/u156  (\U_AHB/n40 [14], gpio_out[14], \U_AHB/n39 [14]);  // src/AHB.v(64)
  and \U_AHB/u157  (\U_AHB/n40 [13], gpio_out[13], \U_AHB/n39 [13]);  // src/AHB.v(64)
  and \U_AHB/u158  (\U_AHB/n40 [12], gpio_out[12], \U_AHB/n39 [12]);  // src/AHB.v(64)
  and \U_AHB/u159  (\U_AHB/n40 [11], gpio_out[11], \U_AHB/n39 [11]);  // src/AHB.v(64)
  or \U_AHB/u16  (\U_AHB/n37 [17], gpio_out[17], \U_AHB/h2h_hwdata [17]);  // src/AHB.v(63)
  and \U_AHB/u160  (\U_AHB/n40 [10], gpio_out[10], \U_AHB/n39 [10]);  // src/AHB.v(64)
  and \U_AHB/u161  (\U_AHB/n40 [9], gpio_out[9], \U_AHB/n39 [9]);  // src/AHB.v(64)
  and \U_AHB/u162  (\U_AHB/n40 [8], gpio_out[8], \U_AHB/n39 [8]);  // src/AHB.v(64)
  and \U_AHB/u163  (\U_AHB/n40 [7], gpio_out[7], \U_AHB/n39 [7]);  // src/AHB.v(64)
  and \U_AHB/u164  (\U_AHB/n40 [6], gpio_out[6], \U_AHB/n39 [6]);  // src/AHB.v(64)
  and \U_AHB/u165  (\U_AHB/n40 [5], gpio_out[5], \U_AHB/n39 [5]);  // src/AHB.v(64)
  and \U_AHB/u166  (\U_AHB/n40 [4], gpio_out[4], \U_AHB/n39 [4]);  // src/AHB.v(64)
  and \U_AHB/u167  (\U_AHB/n40 [3], gpio_out[3], \U_AHB/n39 [3]);  // src/AHB.v(64)
  and \U_AHB/u168  (\U_AHB/n40 [2], gpio_out[2], \U_AHB/n39 [2]);  // src/AHB.v(64)
  and \U_AHB/u169  (\U_AHB/n40 [1], gpio_out[1], \U_AHB/n39 [1]);  // src/AHB.v(64)
  and \U_AHB/u17  (\U_AHB/n14 , \U_AHB/n7 , \U_AHB/h2h_haddr [5]);  // src/AHB.v(51)
  and \U_AHB/u170  (\U_AHB/n40 [0], gpio_out[0], \U_AHB/n39 [0]);  // src/AHB.v(64)
  or \U_AHB/u18  (\U_AHB/n37 [16], gpio_out[16], \U_AHB/h2h_hwdata [16]);  // src/AHB.v(63)
  or \U_AHB/u19  (\U_AHB/n37 [15], gpio_out[15], \U_AHB/h2h_hwdata [15]);  // src/AHB.v(63)
  and \U_AHB/u2  (\U_AHB/n1 , \U_AHB/h2h_hwrite , \U_AHB/n0 );  // src/AHB.v(46)
  and \U_AHB/u20  (\U_AHB/n16 , \U_AHB/n7 , \U_AHB/h2h_haddr [6]);  // src/AHB.v(52)
  or \U_AHB/u21  (\U_AHB/n37 [14], gpio_out[14], \U_AHB/h2h_hwdata [14]);  // src/AHB.v(63)
  or \U_AHB/u22  (\U_AHB/n37 [13], gpio_out[13], \U_AHB/h2h_hwdata [13]);  // src/AHB.v(63)
  and \U_AHB/u23  (\U_AHB/n18 , \U_AHB/n7 , \U_AHB/h2h_haddr [7]);  // src/AHB.v(53)
  or \U_AHB/u24  (\U_AHB/n37 [12], gpio_out[12], \U_AHB/h2h_hwdata [12]);  // src/AHB.v(63)
  or \U_AHB/u25  (\U_AHB/n37 [11], gpio_out[11], \U_AHB/h2h_hwdata [11]);  // src/AHB.v(63)
  and \U_AHB/u26  (\U_AHB/n20 , \U_AHB/n7 , \U_AHB/h2h_haddr [8]);  // src/AHB.v(54)
  or \U_AHB/u27  (\U_AHB/n37 [10], gpio_out[10], \U_AHB/h2h_hwdata [10]);  // src/AHB.v(63)
  or \U_AHB/u28  (\U_AHB/n37 [9], gpio_out[9], \U_AHB/h2h_hwdata [9]);  // src/AHB.v(63)
  and \U_AHB/u29  (\U_AHB/n22 , \U_AHB/n7 , \U_AHB/h2h_haddr [9]);  // src/AHB.v(55)
  and \U_AHB/u3  (\U_AHB/n2 , \U_AHB/n1 , \U_AHB/h2h_haddr [5]);  // src/AHB.v(46)
  or \U_AHB/u30  (\U_AHB/n37 [8], gpio_out[8], \U_AHB/h2h_hwdata [8]);  // src/AHB.v(63)
  or \U_AHB/u31  (\U_AHB/n37 [7], gpio_out[7], \U_AHB/h2h_hwdata [7]);  // src/AHB.v(63)
  and \U_AHB/u32  (\U_AHB/n24 , \U_AHB/n7 , \U_AHB/h2h_haddr [10]);  // src/AHB.v(56)
  or \U_AHB/u33  (\U_AHB/n37 [6], gpio_out[6], \U_AHB/h2h_hwdata [6]);  // src/AHB.v(63)
  or \U_AHB/u34  (\U_AHB/n37 [5], gpio_out[5], \U_AHB/h2h_hwdata [5]);  // src/AHB.v(63)
  and \U_AHB/u35  (\U_AHB/n26 , \U_AHB/n7 , \U_AHB/h2h_haddr [11]);  // src/AHB.v(57)
  or \U_AHB/u36  (\U_AHB/n37 [4], gpio_out[4], \U_AHB/h2h_hwdata [4]);  // src/AHB.v(63)
  or \U_AHB/u37  (\U_AHB/n37 [3], gpio_out[3], \U_AHB/h2h_hwdata [3]);  // src/AHB.v(63)
  and \U_AHB/u38  (\U_AHB/n28 , \U_AHB/n7 , \U_AHB/h2h_haddr [12]);  // src/AHB.v(58)
  or \U_AHB/u39  (\U_AHB/n37 [2], gpio_out[2], \U_AHB/h2h_hwdata [2]);  // src/AHB.v(63)
  or \U_AHB/u4  (\U_AHB/n37 [24], gpio_out[24], \U_AHB/h2h_hwdata [24]);  // src/AHB.v(63)
  or \U_AHB/u40  (\U_AHB/n37 [1], gpio_out[1], \U_AHB/h2h_hwdata [1]);  // src/AHB.v(63)
  and \U_AHB/u41  (\U_AHB/n30 , \U_AHB/n1 , \U_AHB/h2h_haddr [2]);  // src/AHB.v(60)
  not \U_AHB/u42  (\U_AHB/n39 [31], \U_AHB/h2h_hwdata [31]);  // src/AHB.v(64)
  not \U_AHB/u43  (\U_AHB/n39 [30], \U_AHB/h2h_hwdata [30]);  // src/AHB.v(64)
  and \U_AHB/u44  (\U_AHB/n32 , \U_AHB/n1 , \U_AHB/h2h_haddr [3]);  // src/AHB.v(61)
  not \U_AHB/u45  (\U_AHB/n39 [29], \U_AHB/h2h_hwdata [29]);  // src/AHB.v(64)
  not \U_AHB/u46  (\U_AHB/n39 [28], \U_AHB/h2h_hwdata [28]);  // src/AHB.v(64)
  and \U_AHB/u47  (\U_AHB/n34 , \U_AHB/n1 , \U_AHB/h2h_haddr [4]);  // src/AHB.v(62)
  not \U_AHB/u48  (\U_AHB/n39 [27], \U_AHB/h2h_hwdata [27]);  // src/AHB.v(64)
  not \U_AHB/u49  (\U_AHB/n39 [26], \U_AHB/h2h_hwdata [26]);  // src/AHB.v(64)
  or \U_AHB/u5  (\U_AHB/n37 [23], gpio_out[23], \U_AHB/h2h_hwdata [23]);  // src/AHB.v(63)
  and \U_AHB/u50  (\U_AHB/n36 , \U_AHB/n1 , \U_AHB/h2h_haddr [7]);  // src/AHB.v(63)
  not \U_AHB/u51  (\U_AHB/n39 [25], \U_AHB/h2h_hwdata [25]);  // src/AHB.v(64)
  not \U_AHB/u52  (\U_AHB/n39 [24], \U_AHB/h2h_hwdata [24]);  // src/AHB.v(64)
  and \U_AHB/u53  (\U_AHB/n38 , \U_AHB/n1 , \U_AHB/h2h_haddr [8]);  // src/AHB.v(64)
  or \U_AHB/u54  (\U_AHB/n37 [0], gpio_out[0], \U_AHB/h2h_hwdata [0]);  // src/AHB.v(63)
  not \U_AHB/u55  (\U_AHB/n39 [0], \U_AHB/h2h_hwdata [0]);  // src/AHB.v(64)
  and \U_AHB/u56  (\U_AHB/n44 , \U_AHB/h2h_hwrite , \U_AHB/n43 );  // src/AHB.v(67)
  and \U_AHB/u57  (\U_AHB/n45 , \U_AHB/n44 , \U_AHB/h2h_haddr [5]);  // src/AHB.v(67)
  not \U_AHB/u58  (\U_AHB/n39 [23], \U_AHB/h2h_hwdata [23]);  // src/AHB.v(64)
  not \U_AHB/u59  (\U_AHB/n39 [22], \U_AHB/h2h_hwdata [22]);  // src/AHB.v(64)
  and \U_AHB/u6  (\U_AHB/n4 , \U_AHB/n1 , \U_AHB/h2h_haddr [6]);  // src/AHB.v(47)
  and \U_AHB/u60  (\U_AHB/n47 , \U_AHB/n44 , \U_AHB/h2h_haddr [6]);  // src/AHB.v(68)
  and \U_AHB/u61  (\U_AHB/n50 , \U_AHB/h2h_hwrite , \U_AHB/n49 );  // src/AHB.v(69)
  and \U_AHB/u62  (\U_AHB/n51 , \U_AHB/n50 , \U_AHB/h2h_haddr [2]);  // src/AHB.v(69)
  not \U_AHB/u63  (\U_AHB/n39 [21], \U_AHB/h2h_hwdata [21]);  // src/AHB.v(64)
  not \U_AHB/u64  (\U_AHB/n39 [20], \U_AHB/h2h_hwdata [20]);  // src/AHB.v(64)
  and \U_AHB/u65  (\U_AHB/n53 , \U_AHB/n50 , \U_AHB/h2h_haddr [3]);  // src/AHB.v(70)
  not \U_AHB/u66  (\U_AHB/n39 [19], \U_AHB/h2h_hwdata [19]);  // src/AHB.v(64)
  not \U_AHB/u67  (\U_AHB/n39 [18], \U_AHB/h2h_hwdata [18]);  // src/AHB.v(64)
  and \U_AHB/u68  (\U_AHB/n55 , \U_AHB/n50 , \U_AHB/h2h_haddr [4]);  // src/AHB.v(71)
  not \U_AHB/u69  (\U_AHB/n39 [17], \U_AHB/h2h_hwdata [17]);  // src/AHB.v(64)
  and \U_AHB/u7  (\U_AHB/n7 , \U_AHB/h2h_hwrite , \U_AHB/n6 );  // src/AHB.v(48)
  not \U_AHB/u70  (\U_AHB/n39 [16], \U_AHB/h2h_hwdata [16]);  // src/AHB.v(64)
  and \U_AHB/u71  (\U_AHB/n57 , \U_AHB/n50 , \U_AHB/h2h_haddr [5]);  // src/AHB.v(72)
  not \U_AHB/u72  (\U_AHB/n39 [15], \U_AHB/h2h_hwdata [15]);  // src/AHB.v(64)
  not \U_AHB/u73  (\U_AHB/n39 [14], \U_AHB/h2h_hwdata [14]);  // src/AHB.v(64)
  and \U_AHB/u74  (\U_AHB/n59 , \U_AHB/n50 , \U_AHB/h2h_haddr [6]);  // src/AHB.v(73)
  not \U_AHB/u75  (\U_AHB/n39 [13], \U_AHB/h2h_hwdata [13]);  // src/AHB.v(64)
  not \U_AHB/u76  (\U_AHB/n39 [12], \U_AHB/h2h_hwdata [12]);  // src/AHB.v(64)
  and \U_AHB/u77  (\U_AHB/n61 , \U_AHB/n50 , \U_AHB/h2h_haddr [7]);  // src/AHB.v(74)
  not \U_AHB/u78  (\U_AHB/n39 [11], \U_AHB/h2h_hwdata [11]);  // src/AHB.v(64)
  not \U_AHB/u79  (\U_AHB/n39 [10], \U_AHB/h2h_hwdata [10]);  // src/AHB.v(64)
  and \U_AHB/u8  (\U_AHB/n8 , \U_AHB/n7 , \U_AHB/h2h_haddr [2]);  // src/AHB.v(48)
  and \U_AHB/u80  (\U_AHB/n63 , \U_AHB/n50 , \U_AHB/h2h_haddr [8]);  // src/AHB.v(75)
  not \U_AHB/u81  (\U_AHB/n39 [9], \U_AHB/h2h_hwdata [9]);  // src/AHB.v(64)
  not \U_AHB/u82  (\U_AHB/n39 [8], \U_AHB/h2h_hwdata [8]);  // src/AHB.v(64)
  and \U_AHB/u83  (\U_AHB/n65 , \U_AHB/n50 , \U_AHB/h2h_haddr [9]);  // src/AHB.v(76)
  not \U_AHB/u84  (\U_AHB/n39 [7], \U_AHB/h2h_hwdata [7]);  // src/AHB.v(64)
  not \U_AHB/u85  (\U_AHB/n39 [6], \U_AHB/h2h_hwdata [6]);  // src/AHB.v(64)
  and \U_AHB/u86  (\U_AHB/n67 , \U_AHB/n50 , \U_AHB/h2h_haddr [10]);  // src/AHB.v(77)
  not \U_AHB/u87  (\U_AHB/n39 [5], \U_AHB/h2h_hwdata [5]);  // src/AHB.v(64)
  not \U_AHB/u88  (\U_AHB/n39 [4], \U_AHB/h2h_hwdata [4]);  // src/AHB.v(64)
  and \U_AHB/u89  (\U_AHB/n69 , \U_AHB/n50 , \U_AHB/h2h_haddr [11]);  // src/AHB.v(78)
  or \U_AHB/u9  (\U_AHB/n37 [22], gpio_out[22], \U_AHB/h2h_hwdata [22]);  // src/AHB.v(63)
  not \U_AHB/u90  (\U_AHB/n39 [3], \U_AHB/h2h_hwdata [3]);  // src/AHB.v(64)
  not \U_AHB/u91  (\U_AHB/n39 [2], \U_AHB/h2h_hwdata [2]);  // src/AHB.v(64)
  and \U_AHB/u92  (\U_AHB/n71 , \U_AHB/n50 , \U_AHB/h2h_haddr [12]);  // src/AHB.v(79)
  not \U_AHB/u93  (\U_AHB/n39 [1], \U_AHB/h2h_hwdata [1]);  // src/AHB.v(64)
  and \U_AHB/u94  (\U_AHB/n40 [31], gpio_out[31], \U_AHB/n39 [31]);  // src/AHB.v(64)
  and \U_AHB/u95  (\U_AHB/n73 , \U_AHB/n44 , \U_AHB/h2h_haddr [2]);  // src/AHB.v(80)
  and \U_AHB/u96  (\U_AHB/n40 [30], gpio_out[30], \U_AHB/n39 [30]);  // src/AHB.v(64)
  and \U_AHB/u97  (\U_AHB/n40 [29], gpio_out[29], \U_AHB/n39 [29]);  // src/AHB.v(64)
  and \U_AHB/u98  (\U_AHB/n75 , \U_AHB/n44 , \U_AHB/h2h_haddr [3]);  // src/AHB.v(81)
  and \U_AHB/u99  (\U_AHB/n40 [28], gpio_out[28], \U_AHB/n39 [28]);  // src/AHB.v(64)
  EF2_PHY_PLL #(
    .CLKC0_CPHASE(4),
    .CLKC0_DIV(5),
    .CLKC0_DIV2_ENABLE("DISABLE"),
    .CLKC0_DUTY(0.500000),
    .CLKC0_DUTY50("ENABLE"),
    .CLKC0_DUTY_INT(3),
    .CLKC0_ENABLE("ENABLE"),
    .CLKC0_FPHASE(0),
    .CLKC1_CPHASE(9),
    .CLKC1_DIV(10),
    .CLKC1_DIV2_ENABLE("DISABLE"),
    .CLKC1_DUTY(0.500000),
    .CLKC1_DUTY50("ENABLE"),
    .CLKC1_DUTY_INT(5),
    .CLKC1_ENABLE("ENABLE"),
    .CLKC1_FPHASE(0),
    .CLKC2_CPHASE(39),
    .CLKC2_DIV(40),
    .CLKC2_DIV2_ENABLE("DISABLE"),
    .CLKC2_ENABLE("ENABLE"),
    .CLKC2_FPHASE(0),
    .CLKC3_CPHASE(124),
    .CLKC3_DIV(125),
    .CLKC3_DIV2_ENABLE("DISABLE"),
    .CLKC3_ENABLE("ENABLE"),
    .CLKC3_FPHASE(0),
    .CLKC4_CPHASE(1),
    .CLKC4_DIV(1),
    .CLKC4_DIV2_ENABLE("DISABLE"),
    .CLKC4_ENABLE("DISABLE"),
    .CLKC4_FPHASE(0),
    .CLKC5_CPHASE(1),
    .CLKC5_DIV(1),
    .CLKC5_DIV2_ENABLE("DISABLE"),
    .CLKC5_ENABLE("DISABLE"),
    .CLKC6_CPHASE(1),
    .CLKC6_DIV(1),
    .CLKC6_DIV2_ENABLE("DISABLE"),
    .CLKC6_ENABLE("DISABLE"),
    .DERIVE_PLL_CLOCKS("DISABLE"),
    .DPHASE_SOURCE("DISABLE"),
    .DYNCFG("DISABLE"),
    .FBCLK_DIV(40),
    .FEEDBK_MODE("NOCOMP"),
    .FEEDBK_PATH("VCO_PHASE_0"),
    .FIN("25.000"),
    .FREQ_LOCK_ACCURACY(2),
    .FREQ_OFFSET("0.000000"),
    .FREQ_OFFSET_INT("0"),
    .GEN_BASIC_CLOCK("DISABLE"),
    .GMC_GAIN(6),
    .GMC_TEST(14),
    .HIGH_SPEED_EN("ENABLE"),
    .ICP_CURRENT(3),
    .IF_ESCLKSTSW("DISABLE"),
    .INTFB_WAKE("DISABLE"),
    .INTPI(3),
    .KVCO(6),
    .LPF_CAPACITOR(3),
    .LPF_RESISTOR(2),
    .NORESET("DISABLE"),
    .ODIV_MUXC0("DIV"),
    .ODIV_MUXC1("DIV"),
    .ODIV_MUXC2("DIV"),
    .ODIV_MUXC3("DIV"),
    .ODIV_MUXC4("DIV"),
    .OFFSET_MODE("EXT"),
    .PLLC2RST_ENA("DISABLE"),
    .PLLC34RST_ENA("DISABLE"),
    .PLLMRST_ENA("DISABLE"),
    .PLLRST_ENA("ENABLE"),
    .PLL_LOCK_MODE(0),
    .PREDIV_MUXC0("VCO"),
    .PREDIV_MUXC1("VCO"),
    .PREDIV_MUXC2("VCO"),
    .PREDIV_MUXC3("VCO"),
    .PREDIV_MUXC4("VCO"),
    .PREDIV_MUXC5("VCO"),
    .PREDIV_MUXC6("VCO"),
    .PU_INTP("DISABLE"),
    .REFCLK_DIV(1),
    .REFCLK_SEL("INTERNAL"),
    .SSC_AMP("0.000000"),
    .SSC_ENABLE("DISABLE"),
    .SSC_FREQ_DIV(0),
    .SSC_MODE("Down"),
    .SSC_RNGE(0),
    .STDBY_ENABLE("DISABLE"),
    .STDBY_VCO_ENA("DISABLE"),
    .SYNC_ENABLE("DISABLE"),
    .VCO_NORESET("DISABLE"))
    \U_PLL/pll_inst  (
    .daddr(6'b000000),
    .dclk(1'b0),
    .dcs(1'b0),
    .di(8'b00000000),
    .dsm_refclk(1'b0),
    .dsm_rst(1'b0),
    .dwe(1'b0),
    .fbclk(1'b0),
    .frac_offset_valid(1'b0),
    .psclk(1'b0),
    .psclksel(3'b000),
    .psdown(1'b0),
    .psstep(1'b0),
    .refclk(clkin),
    .reset(1'b0),
    .ssc_en(1'b0),
    .stdby(1'b0),
    .clkc({open_n101,open_n102,open_n103,open_n104,clk25m,clk100m,open_n105}),
    .extlock(rstn));  // al_ip/PLL.v(92)
  add_pu32_pu32_o32 add0 (
    .i0(timer),
    .i1(32'b00000000000000000000000000000001),
    .o(n2));  // CPLD_SOC_AHB_TOP.v(35)
  eq_w32 eq0 (
    .i0(timer),
    .i1(32'b00001011111010111100000111111111),
    .o(n1));  // CPLD_SOC_AHB_TOP.v(32)
  eq_w32 eq1 (
    .i0(timer),
    .i1(32'b00000010111110101111000001111111),
    .o(n4));  // CPLD_SOC_AHB_TOP.v(42)
  eq_w32 eq2 (
    .i0(timer),
    .i1(32'b00000101111101011110000011111111),
    .o(n5));  // CPLD_SOC_AHB_TOP.v(44)
  eq_w32 eq3 (
    .i0(timer),
    .i1(32'b00001000111100001101000101111111),
    .o(n6));  // CPLD_SOC_AHB_TOP.v(46)
  binary_mux_s1_w1 mux0_b0 (
    .i0(n2[0]),
    .i1(1'b0),
    .sel(n1),
    .o(n3[0]));  // CPLD_SOC_AHB_TOP.v(35)
  binary_mux_s1_w1 mux0_b1 (
    .i0(n2[1]),
    .i1(1'b0),
    .sel(n1),
    .o(n3[1]));  // CPLD_SOC_AHB_TOP.v(35)
  binary_mux_s1_w1 mux0_b10 (
    .i0(n2[10]),
    .i1(1'b0),
    .sel(n1),
    .o(n3[10]));  // CPLD_SOC_AHB_TOP.v(35)
  binary_mux_s1_w1 mux0_b11 (
    .i0(n2[11]),
    .i1(1'b0),
    .sel(n1),
    .o(n3[11]));  // CPLD_SOC_AHB_TOP.v(35)
  binary_mux_s1_w1 mux0_b12 (
    .i0(n2[12]),
    .i1(1'b0),
    .sel(n1),
    .o(n3[12]));  // CPLD_SOC_AHB_TOP.v(35)
  binary_mux_s1_w1 mux0_b13 (
    .i0(n2[13]),
    .i1(1'b0),
    .sel(n1),
    .o(n3[13]));  // CPLD_SOC_AHB_TOP.v(35)
  binary_mux_s1_w1 mux0_b14 (
    .i0(n2[14]),
    .i1(1'b0),
    .sel(n1),
    .o(n3[14]));  // CPLD_SOC_AHB_TOP.v(35)
  binary_mux_s1_w1 mux0_b15 (
    .i0(n2[15]),
    .i1(1'b0),
    .sel(n1),
    .o(n3[15]));  // CPLD_SOC_AHB_TOP.v(35)
  binary_mux_s1_w1 mux0_b16 (
    .i0(n2[16]),
    .i1(1'b0),
    .sel(n1),
    .o(n3[16]));  // CPLD_SOC_AHB_TOP.v(35)
  binary_mux_s1_w1 mux0_b17 (
    .i0(n2[17]),
    .i1(1'b0),
    .sel(n1),
    .o(n3[17]));  // CPLD_SOC_AHB_TOP.v(35)
  binary_mux_s1_w1 mux0_b18 (
    .i0(n2[18]),
    .i1(1'b0),
    .sel(n1),
    .o(n3[18]));  // CPLD_SOC_AHB_TOP.v(35)
  binary_mux_s1_w1 mux0_b19 (
    .i0(n2[19]),
    .i1(1'b0),
    .sel(n1),
    .o(n3[19]));  // CPLD_SOC_AHB_TOP.v(35)
  binary_mux_s1_w1 mux0_b2 (
    .i0(n2[2]),
    .i1(1'b0),
    .sel(n1),
    .o(n3[2]));  // CPLD_SOC_AHB_TOP.v(35)
  binary_mux_s1_w1 mux0_b20 (
    .i0(n2[20]),
    .i1(1'b0),
    .sel(n1),
    .o(n3[20]));  // CPLD_SOC_AHB_TOP.v(35)
  binary_mux_s1_w1 mux0_b21 (
    .i0(n2[21]),
    .i1(1'b0),
    .sel(n1),
    .o(n3[21]));  // CPLD_SOC_AHB_TOP.v(35)
  binary_mux_s1_w1 mux0_b22 (
    .i0(n2[22]),
    .i1(1'b0),
    .sel(n1),
    .o(n3[22]));  // CPLD_SOC_AHB_TOP.v(35)
  binary_mux_s1_w1 mux0_b23 (
    .i0(n2[23]),
    .i1(1'b0),
    .sel(n1),
    .o(n3[23]));  // CPLD_SOC_AHB_TOP.v(35)
  binary_mux_s1_w1 mux0_b24 (
    .i0(n2[24]),
    .i1(1'b0),
    .sel(n1),
    .o(n3[24]));  // CPLD_SOC_AHB_TOP.v(35)
  binary_mux_s1_w1 mux0_b25 (
    .i0(n2[25]),
    .i1(1'b0),
    .sel(n1),
    .o(n3[25]));  // CPLD_SOC_AHB_TOP.v(35)
  binary_mux_s1_w1 mux0_b26 (
    .i0(n2[26]),
    .i1(1'b0),
    .sel(n1),
    .o(n3[26]));  // CPLD_SOC_AHB_TOP.v(35)
  binary_mux_s1_w1 mux0_b27 (
    .i0(n2[27]),
    .i1(1'b0),
    .sel(n1),
    .o(n3[27]));  // CPLD_SOC_AHB_TOP.v(35)
  binary_mux_s1_w1 mux0_b28 (
    .i0(n2[28]),
    .i1(1'b0),
    .sel(n1),
    .o(n3[28]));  // CPLD_SOC_AHB_TOP.v(35)
  binary_mux_s1_w1 mux0_b29 (
    .i0(n2[29]),
    .i1(1'b0),
    .sel(n1),
    .o(n3[29]));  // CPLD_SOC_AHB_TOP.v(35)
  binary_mux_s1_w1 mux0_b3 (
    .i0(n2[3]),
    .i1(1'b0),
    .sel(n1),
    .o(n3[3]));  // CPLD_SOC_AHB_TOP.v(35)
  binary_mux_s1_w1 mux0_b30 (
    .i0(n2[30]),
    .i1(1'b0),
    .sel(n1),
    .o(n3[30]));  // CPLD_SOC_AHB_TOP.v(35)
  binary_mux_s1_w1 mux0_b31 (
    .i0(n2[31]),
    .i1(1'b0),
    .sel(n1),
    .o(n3[31]));  // CPLD_SOC_AHB_TOP.v(35)
  binary_mux_s1_w1 mux0_b4 (
    .i0(n2[4]),
    .i1(1'b0),
    .sel(n1),
    .o(n3[4]));  // CPLD_SOC_AHB_TOP.v(35)
  binary_mux_s1_w1 mux0_b5 (
    .i0(n2[5]),
    .i1(1'b0),
    .sel(n1),
    .o(n3[5]));  // CPLD_SOC_AHB_TOP.v(35)
  binary_mux_s1_w1 mux0_b6 (
    .i0(n2[6]),
    .i1(1'b0),
    .sel(n1),
    .o(n3[6]));  // CPLD_SOC_AHB_TOP.v(35)
  binary_mux_s1_w1 mux0_b7 (
    .i0(n2[7]),
    .i1(1'b0),
    .sel(n1),
    .o(n3[7]));  // CPLD_SOC_AHB_TOP.v(35)
  binary_mux_s1_w1 mux0_b8 (
    .i0(n2[8]),
    .i1(1'b0),
    .sel(n1),
    .o(n3[8]));  // CPLD_SOC_AHB_TOP.v(35)
  binary_mux_s1_w1 mux0_b9 (
    .i0(n2[9]),
    .i1(1'b0),
    .sel(n1),
    .o(n3[9]));  // CPLD_SOC_AHB_TOP.v(35)
  binary_mux_s1_w1 mux1_b2 (
    .i0(ledout[2]),
    .i1(1'b1),
    .sel(n1),
    .o(n7[2]));  // CPLD_SOC_AHB_TOP.v(49)
  binary_mux_s1_w1 mux1_b3 (
    .i0(ledout[3]),
    .i1(1'b0),
    .sel(n1),
    .o(n7[3]));  // CPLD_SOC_AHB_TOP.v(49)
  and mux2_b0_sel_is_0 (mux2_b0_sel_is_0_o, n6_neg, n1_neg);
  AL_MUX mux2_b1 (
    .i0(1'b1),
    .i1(ledout[1]),
    .sel(mux2_b0_sel_is_0_o),
    .o(n8[1]));
  binary_mux_s1_w1 mux2_b2 (
    .i0(n7[2]),
    .i1(1'b0),
    .sel(n6),
    .o(n8[2]));  // CPLD_SOC_AHB_TOP.v(49)
  and mux3_b0_sel_is_2 (mux3_b0_sel_is_2_o, n5_neg, mux2_b0_sel_is_0_o);
  binary_mux_s1_w1 mux3_b1 (
    .i0(n8[1]),
    .i1(1'b0),
    .sel(n5),
    .o(n9[1]));  // CPLD_SOC_AHB_TOP.v(49)
  and mux3_b3_sel_is_0 (mux3_b3_sel_is_0_o, n5_neg, n6_neg);
  binary_mux_s1_w1 mux4_b1 (
    .i0(n9[1]),
    .i1(1'b1),
    .sel(n4),
    .o(n10[1]));  // CPLD_SOC_AHB_TOP.v(49)
  AL_MUX mux4_b2 (
    .i0(1'b1),
    .i1(n8[2]),
    .sel(mux4_b2_sel_is_0_o),
    .o(n10[2]));
  and mux4_b2_sel_is_0 (mux4_b2_sel_is_0_o, n4_neg, n5_neg);
  AL_MUX mux4_b3 (
    .i0(1'b1),
    .i1(n7[3]),
    .sel(mux4_b3_sel_is_2_o),
    .o(n10[3]));
  and mux4_b3_sel_is_2 (mux4_b3_sel_is_2_o, n4_neg, mux3_b3_sel_is_0_o);
  not n1_inv (n1_neg, n1);
  not n4_inv (n4_neg, n4);
  not n5_inv (n5_neg, n5);
  not n6_inv (n6_neg, n6);
  not \pwm_start_stop[16]_inv  (\pwm_start_stop[16]_neg , pwm_start_stop[16]);
  not \pwm_start_stop[17]_inv  (\pwm_start_stop[17]_neg , pwm_start_stop[17]);
  not \pwm_start_stop[18]_inv  (\pwm_start_stop[18]_neg , pwm_start_stop[18]);
  not \pwm_start_stop[19]_inv  (\pwm_start_stop[19]_neg , pwm_start_stop[19]);
  not \pwm_start_stop[20]_inv  (\pwm_start_stop[20]_neg , pwm_start_stop[20]);
  not \pwm_start_stop[21]_inv  (\pwm_start_stop[21]_neg , pwm_start_stop[21]);
  not \pwm_start_stop[22]_inv  (\pwm_start_stop[22]_neg , pwm_start_stop[22]);
  not \pwm_start_stop[23]_inv  (\pwm_start_stop[23]_neg , pwm_start_stop[23]);
  not \pwm_start_stop[24]_inv  (\pwm_start_stop[24]_neg , pwm_start_stop[24]);
  not \pwm_start_stop[25]_inv  (\pwm_start_stop[25]_neg , pwm_start_stop[25]);
  not \pwm_start_stop[26]_inv  (\pwm_start_stop[26]_neg , pwm_start_stop[26]);
  not \pwm_start_stop[27]_inv  (\pwm_start_stop[27]_neg , pwm_start_stop[27]);
  not \pwm_start_stop[28]_inv  (\pwm_start_stop[28]_neg , pwm_start_stop[28]);
  not \pwm_start_stop[29]_inv  (\pwm_start_stop[29]_neg , pwm_start_stop[29]);
  not \pwm_start_stop[30]_inv  (\pwm_start_stop[30]_neg , pwm_start_stop[30]);
  not \pwm_start_stop[31]_inv  (\pwm_start_stop[31]_neg , pwm_start_stop[31]);
  reg_ar_as_w1 reg0_b0 (
    .clk(clk25m),
    .d(n3[0]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(timer[0]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b1 (
    .clk(clk25m),
    .d(n3[1]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(timer[1]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b10 (
    .clk(clk25m),
    .d(n3[10]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(timer[10]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b11 (
    .clk(clk25m),
    .d(n3[11]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(timer[11]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b12 (
    .clk(clk25m),
    .d(n3[12]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(timer[12]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b13 (
    .clk(clk25m),
    .d(n3[13]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(timer[13]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b14 (
    .clk(clk25m),
    .d(n3[14]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(timer[14]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b15 (
    .clk(clk25m),
    .d(n3[15]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(timer[15]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b16 (
    .clk(clk25m),
    .d(n3[16]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(timer[16]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b17 (
    .clk(clk25m),
    .d(n3[17]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(timer[17]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b18 (
    .clk(clk25m),
    .d(n3[18]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(timer[18]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b19 (
    .clk(clk25m),
    .d(n3[19]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(timer[19]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b2 (
    .clk(clk25m),
    .d(n3[2]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(timer[2]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b20 (
    .clk(clk25m),
    .d(n3[20]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(timer[20]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b21 (
    .clk(clk25m),
    .d(n3[21]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(timer[21]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b22 (
    .clk(clk25m),
    .d(n3[22]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(timer[22]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b23 (
    .clk(clk25m),
    .d(n3[23]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(timer[23]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b24 (
    .clk(clk25m),
    .d(n3[24]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(timer[24]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b25 (
    .clk(clk25m),
    .d(n3[25]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(timer[25]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b26 (
    .clk(clk25m),
    .d(n3[26]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(timer[26]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b27 (
    .clk(clk25m),
    .d(n3[27]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(timer[27]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b28 (
    .clk(clk25m),
    .d(n3[28]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(timer[28]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b29 (
    .clk(clk25m),
    .d(n3[29]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(timer[29]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b3 (
    .clk(clk25m),
    .d(n3[3]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(timer[3]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b30 (
    .clk(clk25m),
    .d(n3[30]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(timer[30]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b31 (
    .clk(clk25m),
    .d(n3[31]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(timer[31]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b4 (
    .clk(clk25m),
    .d(n3[4]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(timer[4]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b5 (
    .clk(clk25m),
    .d(n3[5]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(timer[5]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b6 (
    .clk(clk25m),
    .d(n3[6]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(timer[6]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b7 (
    .clk(clk25m),
    .d(n3[7]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(timer[7]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b8 (
    .clk(clk25m),
    .d(n3[8]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(timer[8]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_ar_as_w1 reg0_b9 (
    .clk(clk25m),
    .d(n3[9]),
    .en(1'b1),
    .reset(~rst_n),
    .set(1'b0),
    .q(timer[9]));  // CPLD_SOC_AHB_TOP.v(35)
  reg_sr_as_w1 reg1_b0 (
    .clk(clk25m),
    .d(1'b1),
    .en(~mux3_b0_sel_is_2_o),
    .reset(n4),
    .set(~rst_n),
    .q(ledout[0]));  // CPLD_SOC_AHB_TOP.v(49)
  reg_ar_as_w1 reg1_b1 (
    .clk(clk25m),
    .d(n10[1]),
    .en(1'b1),
    .reset(1'b0),
    .set(~rst_n),
    .q(ledout[1]));  // CPLD_SOC_AHB_TOP.v(49)
  reg_ar_as_w1 reg1_b2 (
    .clk(clk25m),
    .d(n10[2]),
    .en(1'b1),
    .reset(1'b0),
    .set(~rst_n),
    .q(ledout[2]));  // CPLD_SOC_AHB_TOP.v(49)
  reg_ar_as_w1 reg1_b3 (
    .clk(clk25m),
    .d(n10[3]),
    .en(1'b1),
    .reset(1'b0),
    .set(~rst_n),
    .q(ledout[3]));  // CPLD_SOC_AHB_TOP.v(49)
  and u10 (n18, limit_l[7], limit_r[7]);  // CPLD_SOC_AHB_TOP.v(127)
  and u11 (n19, limit_l[8], limit_r[8]);  // CPLD_SOC_AHB_TOP.v(128)
  and u12 (n20, limit_l[9], limit_r[9]);  // CPLD_SOC_AHB_TOP.v(129)
  and u13 (n21, limit_l[10], limit_r[10]);  // CPLD_SOC_AHB_TOP.v(130)
  and u14 (n22, limit_l[11], limit_r[11]);  // CPLD_SOC_AHB_TOP.v(131)
  and u15 (n23, limit_l[12], limit_r[12]);  // CPLD_SOC_AHB_TOP.v(132)
  and u16 (n24, limit_l[13], limit_r[13]);  // CPLD_SOC_AHB_TOP.v(133)
  and u17 (n25, limit_l[14], limit_r[14]);  // CPLD_SOC_AHB_TOP.v(134)
  and u18 (n26, limit_l[15], limit_r[15]);  // CPLD_SOC_AHB_TOP.v(135)
  and u3 (n11, limit_l[0], limit_r[0]);  // CPLD_SOC_AHB_TOP.v(120)
  and u4 (n12, limit_l[1], limit_r[1]);  // CPLD_SOC_AHB_TOP.v(121)
  and u5 (n13, limit_l[2], limit_r[2]);  // CPLD_SOC_AHB_TOP.v(122)
  and u6 (n14, limit_l[3], limit_r[3]);  // CPLD_SOC_AHB_TOP.v(123)
  and u7 (n15, limit_l[4], limit_r[4]);  // CPLD_SOC_AHB_TOP.v(124)
  and u8 (n16, limit_l[5], limit_r[5]);  // CPLD_SOC_AHB_TOP.v(125)
  and u9 (n17, limit_l[6], limit_r[6]);  // CPLD_SOC_AHB_TOP.v(126)

endmodule 

module reg_ar_as_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  parameter REGSET = "RESET";
  wire enout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_DFF #(
    .INI((REGSET == "SET") ? 1'b1 : 1'b0))
    u_seq0 (
    .clk(clk),
    .d(enout),
    .reset(reset),
    .set(set),
    .q(q));

endmodule 

module AL_BUFKEEP
  (
  i,
  o
  );

  input i;
  output o;

  parameter KEEP = "OUT";

  buf u1 (o, i);

endmodule 

module eq_w27
  (
  i0,
  i1,
  o
  );

  input [26:0] i0;
  input [26:0] i1;
  output o;

  wire \or_or_or_or_xor_i0[0_o ;
  wire \or_or_or_xor_i0[0]_i_o ;
  wire \or_or_or_xor_i0[13]__o ;
  wire \or_or_xor_i0[0]_i1[0_o ;
  wire \or_or_xor_i0[13]_i1[_o ;
  wire \or_or_xor_i0[16]_i1[_o ;
  wire \or_or_xor_i0[20]_i1[_o ;
  wire \or_or_xor_i0[23]_i1[_o ;
  wire \or_or_xor_i0[6]_i1[6_o ;
  wire \or_or_xor_i0[9]_i1[9_o ;
  wire \or_xor_i0[0]_i1[0]_o_o ;
  wire \or_xor_i0[11]_i1[11]_o ;
  wire \or_xor_i0[13]_i1[13]_o ;
  wire \or_xor_i0[14]_i1[14]_o ;
  wire \or_xor_i0[16]_i1[16]_o ;
  wire \or_xor_i0[18]_i1[18]_o ;
  wire \or_xor_i0[1]_i1[1]_o_o ;
  wire \or_xor_i0[20]_i1[20]_o ;
  wire \or_xor_i0[21]_i1[21]_o ;
  wire \or_xor_i0[23]_i1[23]_o ;
  wire \or_xor_i0[25]_i1[25]_o ;
  wire \or_xor_i0[3]_i1[3]_o_o ;
  wire \or_xor_i0[4]_i1[4]_o_o ;
  wire \or_xor_i0[6]_i1[6]_o_o ;
  wire \or_xor_i0[7]_i1[7]_o_o ;
  wire \or_xor_i0[9]_i1[9]_o_o ;
  wire \xor_i0[0]_i1[0]_o ;
  wire \xor_i0[10]_i1[10]_o ;
  wire \xor_i0[11]_i1[11]_o ;
  wire \xor_i0[12]_i1[12]_o ;
  wire \xor_i0[13]_i1[13]_o ;
  wire \xor_i0[14]_i1[14]_o ;
  wire \xor_i0[15]_i1[15]_o ;
  wire \xor_i0[16]_i1[16]_o ;
  wire \xor_i0[17]_i1[17]_o ;
  wire \xor_i0[18]_i1[18]_o ;
  wire \xor_i0[19]_i1[19]_o ;
  wire \xor_i0[1]_i1[1]_o ;
  wire \xor_i0[20]_i1[20]_o ;
  wire \xor_i0[21]_i1[21]_o ;
  wire \xor_i0[22]_i1[22]_o ;
  wire \xor_i0[23]_i1[23]_o ;
  wire \xor_i0[24]_i1[24]_o ;
  wire \xor_i0[25]_i1[25]_o ;
  wire \xor_i0[26]_i1[26]_o ;
  wire \xor_i0[2]_i1[2]_o ;
  wire \xor_i0[3]_i1[3]_o ;
  wire \xor_i0[4]_i1[4]_o ;
  wire \xor_i0[5]_i1[5]_o ;
  wire \xor_i0[6]_i1[6]_o ;
  wire \xor_i0[7]_i1[7]_o ;
  wire \xor_i0[8]_i1[8]_o ;
  wire \xor_i0[9]_i1[9]_o ;

  not none_diff (o, \or_or_or_or_xor_i0[0_o );
  or \or_or_or_or_xor_i0[0  (\or_or_or_or_xor_i0[0_o , \or_or_or_xor_i0[0]_i_o , \or_or_or_xor_i0[13]__o );
  or \or_or_or_xor_i0[0]_i  (\or_or_or_xor_i0[0]_i_o , \or_or_xor_i0[0]_i1[0_o , \or_or_xor_i0[6]_i1[6_o );
  or \or_or_or_xor_i0[13]_  (\or_or_or_xor_i0[13]__o , \or_or_xor_i0[13]_i1[_o , \or_or_xor_i0[20]_i1[_o );
  or \or_or_xor_i0[0]_i1[0  (\or_or_xor_i0[0]_i1[0_o , \or_xor_i0[0]_i1[0]_o_o , \or_xor_i0[3]_i1[3]_o_o );
  or \or_or_xor_i0[13]_i1[  (\or_or_xor_i0[13]_i1[_o , \or_xor_i0[13]_i1[13]_o , \or_or_xor_i0[16]_i1[_o );
  or \or_or_xor_i0[16]_i1[  (\or_or_xor_i0[16]_i1[_o , \or_xor_i0[16]_i1[16]_o , \or_xor_i0[18]_i1[18]_o );
  or \or_or_xor_i0[20]_i1[  (\or_or_xor_i0[20]_i1[_o , \or_xor_i0[20]_i1[20]_o , \or_or_xor_i0[23]_i1[_o );
  or \or_or_xor_i0[23]_i1[  (\or_or_xor_i0[23]_i1[_o , \or_xor_i0[23]_i1[23]_o , \or_xor_i0[25]_i1[25]_o );
  or \or_or_xor_i0[6]_i1[6  (\or_or_xor_i0[6]_i1[6_o , \or_xor_i0[6]_i1[6]_o_o , \or_or_xor_i0[9]_i1[9_o );
  or \or_or_xor_i0[9]_i1[9  (\or_or_xor_i0[9]_i1[9_o , \or_xor_i0[9]_i1[9]_o_o , \or_xor_i0[11]_i1[11]_o );
  or \or_xor_i0[0]_i1[0]_o  (\or_xor_i0[0]_i1[0]_o_o , \xor_i0[0]_i1[0]_o , \or_xor_i0[1]_i1[1]_o_o );
  or \or_xor_i0[11]_i1[11]  (\or_xor_i0[11]_i1[11]_o , \xor_i0[11]_i1[11]_o , \xor_i0[12]_i1[12]_o );
  or \or_xor_i0[13]_i1[13]  (\or_xor_i0[13]_i1[13]_o , \xor_i0[13]_i1[13]_o , \or_xor_i0[14]_i1[14]_o );
  or \or_xor_i0[14]_i1[14]  (\or_xor_i0[14]_i1[14]_o , \xor_i0[14]_i1[14]_o , \xor_i0[15]_i1[15]_o );
  or \or_xor_i0[16]_i1[16]  (\or_xor_i0[16]_i1[16]_o , \xor_i0[16]_i1[16]_o , \xor_i0[17]_i1[17]_o );
  or \or_xor_i0[18]_i1[18]  (\or_xor_i0[18]_i1[18]_o , \xor_i0[18]_i1[18]_o , \xor_i0[19]_i1[19]_o );
  or \or_xor_i0[1]_i1[1]_o  (\or_xor_i0[1]_i1[1]_o_o , \xor_i0[1]_i1[1]_o , \xor_i0[2]_i1[2]_o );
  or \or_xor_i0[20]_i1[20]  (\or_xor_i0[20]_i1[20]_o , \xor_i0[20]_i1[20]_o , \or_xor_i0[21]_i1[21]_o );
  or \or_xor_i0[21]_i1[21]  (\or_xor_i0[21]_i1[21]_o , \xor_i0[21]_i1[21]_o , \xor_i0[22]_i1[22]_o );
  or \or_xor_i0[23]_i1[23]  (\or_xor_i0[23]_i1[23]_o , \xor_i0[23]_i1[23]_o , \xor_i0[24]_i1[24]_o );
  or \or_xor_i0[25]_i1[25]  (\or_xor_i0[25]_i1[25]_o , \xor_i0[25]_i1[25]_o , \xor_i0[26]_i1[26]_o );
  or \or_xor_i0[3]_i1[3]_o  (\or_xor_i0[3]_i1[3]_o_o , \xor_i0[3]_i1[3]_o , \or_xor_i0[4]_i1[4]_o_o );
  or \or_xor_i0[4]_i1[4]_o  (\or_xor_i0[4]_i1[4]_o_o , \xor_i0[4]_i1[4]_o , \xor_i0[5]_i1[5]_o );
  or \or_xor_i0[6]_i1[6]_o  (\or_xor_i0[6]_i1[6]_o_o , \xor_i0[6]_i1[6]_o , \or_xor_i0[7]_i1[7]_o_o );
  or \or_xor_i0[7]_i1[7]_o  (\or_xor_i0[7]_i1[7]_o_o , \xor_i0[7]_i1[7]_o , \xor_i0[8]_i1[8]_o );
  or \or_xor_i0[9]_i1[9]_o  (\or_xor_i0[9]_i1[9]_o_o , \xor_i0[9]_i1[9]_o , \xor_i0[10]_i1[10]_o );
  xor \xor_i0[0]_i1[0]  (\xor_i0[0]_i1[0]_o , i0[0], i1[0]);
  xor \xor_i0[10]_i1[10]  (\xor_i0[10]_i1[10]_o , i0[10], i1[10]);
  xor \xor_i0[11]_i1[11]  (\xor_i0[11]_i1[11]_o , i0[11], i1[11]);
  xor \xor_i0[12]_i1[12]  (\xor_i0[12]_i1[12]_o , i0[12], i1[12]);
  xor \xor_i0[13]_i1[13]  (\xor_i0[13]_i1[13]_o , i0[13], i1[13]);
  xor \xor_i0[14]_i1[14]  (\xor_i0[14]_i1[14]_o , i0[14], i1[14]);
  xor \xor_i0[15]_i1[15]  (\xor_i0[15]_i1[15]_o , i0[15], i1[15]);
  xor \xor_i0[16]_i1[16]  (\xor_i0[16]_i1[16]_o , i0[16], i1[16]);
  xor \xor_i0[17]_i1[17]  (\xor_i0[17]_i1[17]_o , i0[17], i1[17]);
  xor \xor_i0[18]_i1[18]  (\xor_i0[18]_i1[18]_o , i0[18], i1[18]);
  xor \xor_i0[19]_i1[19]  (\xor_i0[19]_i1[19]_o , i0[19], i1[19]);
  xor \xor_i0[1]_i1[1]  (\xor_i0[1]_i1[1]_o , i0[1], i1[1]);
  xor \xor_i0[20]_i1[20]  (\xor_i0[20]_i1[20]_o , i0[20], i1[20]);
  xor \xor_i0[21]_i1[21]  (\xor_i0[21]_i1[21]_o , i0[21], i1[21]);
  xor \xor_i0[22]_i1[22]  (\xor_i0[22]_i1[22]_o , i0[22], i1[22]);
  xor \xor_i0[23]_i1[23]  (\xor_i0[23]_i1[23]_o , i0[23], i1[23]);
  xor \xor_i0[24]_i1[24]  (\xor_i0[24]_i1[24]_o , i0[24], i1[24]);
  xor \xor_i0[25]_i1[25]  (\xor_i0[25]_i1[25]_o , i0[25], i1[25]);
  xor \xor_i0[26]_i1[26]  (\xor_i0[26]_i1[26]_o , i0[26], i1[26]);
  xor \xor_i0[2]_i1[2]  (\xor_i0[2]_i1[2]_o , i0[2], i1[2]);
  xor \xor_i0[3]_i1[3]  (\xor_i0[3]_i1[3]_o , i0[3], i1[3]);
  xor \xor_i0[4]_i1[4]  (\xor_i0[4]_i1[4]_o , i0[4], i1[4]);
  xor \xor_i0[5]_i1[5]  (\xor_i0[5]_i1[5]_o , i0[5], i1[5]);
  xor \xor_i0[6]_i1[6]  (\xor_i0[6]_i1[6]_o , i0[6], i1[6]);
  xor \xor_i0[7]_i1[7]  (\xor_i0[7]_i1[7]_o , i0[7], i1[7]);
  xor \xor_i0[8]_i1[8]  (\xor_i0[8]_i1[8]_o , i0[8], i1[8]);
  xor \xor_i0[9]_i1[9]  (\xor_i0[9]_i1[9]_o , i0[9], i1[9]);

endmodule 

module eq_w24
  (
  i0,
  i1,
  o
  );

  input [23:0] i0;
  input [23:0] i1;
  output o;

  wire \or_or_or_or_xor_i0[0_o ;
  wire \or_or_or_xor_i0[0]_i_o ;
  wire \or_or_or_xor_i0[12]__o ;
  wire \or_or_xor_i0[0]_i1[0_o ;
  wire \or_or_xor_i0[12]_i1[_o ;
  wire \or_or_xor_i0[18]_i1[_o ;
  wire \or_or_xor_i0[6]_i1[6_o ;
  wire \or_xor_i0[0]_i1[0]_o_o ;
  wire \or_xor_i0[10]_i1[10]_o ;
  wire \or_xor_i0[12]_i1[12]_o ;
  wire \or_xor_i0[13]_i1[13]_o ;
  wire \or_xor_i0[15]_i1[15]_o ;
  wire \or_xor_i0[16]_i1[16]_o ;
  wire \or_xor_i0[18]_i1[18]_o ;
  wire \or_xor_i0[19]_i1[19]_o ;
  wire \or_xor_i0[1]_i1[1]_o_o ;
  wire \or_xor_i0[21]_i1[21]_o ;
  wire \or_xor_i0[22]_i1[22]_o ;
  wire \or_xor_i0[3]_i1[3]_o_o ;
  wire \or_xor_i0[4]_i1[4]_o_o ;
  wire \or_xor_i0[6]_i1[6]_o_o ;
  wire \or_xor_i0[7]_i1[7]_o_o ;
  wire \or_xor_i0[9]_i1[9]_o_o ;
  wire \xor_i0[0]_i1[0]_o ;
  wire \xor_i0[10]_i1[10]_o ;
  wire \xor_i0[11]_i1[11]_o ;
  wire \xor_i0[12]_i1[12]_o ;
  wire \xor_i0[13]_i1[13]_o ;
  wire \xor_i0[14]_i1[14]_o ;
  wire \xor_i0[15]_i1[15]_o ;
  wire \xor_i0[16]_i1[16]_o ;
  wire \xor_i0[17]_i1[17]_o ;
  wire \xor_i0[18]_i1[18]_o ;
  wire \xor_i0[19]_i1[19]_o ;
  wire \xor_i0[1]_i1[1]_o ;
  wire \xor_i0[20]_i1[20]_o ;
  wire \xor_i0[21]_i1[21]_o ;
  wire \xor_i0[22]_i1[22]_o ;
  wire \xor_i0[23]_i1[23]_o ;
  wire \xor_i0[2]_i1[2]_o ;
  wire \xor_i0[3]_i1[3]_o ;
  wire \xor_i0[4]_i1[4]_o ;
  wire \xor_i0[5]_i1[5]_o ;
  wire \xor_i0[6]_i1[6]_o ;
  wire \xor_i0[7]_i1[7]_o ;
  wire \xor_i0[8]_i1[8]_o ;
  wire \xor_i0[9]_i1[9]_o ;

  not none_diff (o, \or_or_or_or_xor_i0[0_o );
  or \or_or_or_or_xor_i0[0  (\or_or_or_or_xor_i0[0_o , \or_or_or_xor_i0[0]_i_o , \or_or_or_xor_i0[12]__o );
  or \or_or_or_xor_i0[0]_i  (\or_or_or_xor_i0[0]_i_o , \or_or_xor_i0[0]_i1[0_o , \or_or_xor_i0[6]_i1[6_o );
  or \or_or_or_xor_i0[12]_  (\or_or_or_xor_i0[12]__o , \or_or_xor_i0[12]_i1[_o , \or_or_xor_i0[18]_i1[_o );
  or \or_or_xor_i0[0]_i1[0  (\or_or_xor_i0[0]_i1[0_o , \or_xor_i0[0]_i1[0]_o_o , \or_xor_i0[3]_i1[3]_o_o );
  or \or_or_xor_i0[12]_i1[  (\or_or_xor_i0[12]_i1[_o , \or_xor_i0[12]_i1[12]_o , \or_xor_i0[15]_i1[15]_o );
  or \or_or_xor_i0[18]_i1[  (\or_or_xor_i0[18]_i1[_o , \or_xor_i0[18]_i1[18]_o , \or_xor_i0[21]_i1[21]_o );
  or \or_or_xor_i0[6]_i1[6  (\or_or_xor_i0[6]_i1[6_o , \or_xor_i0[6]_i1[6]_o_o , \or_xor_i0[9]_i1[9]_o_o );
  or \or_xor_i0[0]_i1[0]_o  (\or_xor_i0[0]_i1[0]_o_o , \xor_i0[0]_i1[0]_o , \or_xor_i0[1]_i1[1]_o_o );
  or \or_xor_i0[10]_i1[10]  (\or_xor_i0[10]_i1[10]_o , \xor_i0[10]_i1[10]_o , \xor_i0[11]_i1[11]_o );
  or \or_xor_i0[12]_i1[12]  (\or_xor_i0[12]_i1[12]_o , \xor_i0[12]_i1[12]_o , \or_xor_i0[13]_i1[13]_o );
  or \or_xor_i0[13]_i1[13]  (\or_xor_i0[13]_i1[13]_o , \xor_i0[13]_i1[13]_o , \xor_i0[14]_i1[14]_o );
  or \or_xor_i0[15]_i1[15]  (\or_xor_i0[15]_i1[15]_o , \xor_i0[15]_i1[15]_o , \or_xor_i0[16]_i1[16]_o );
  or \or_xor_i0[16]_i1[16]  (\or_xor_i0[16]_i1[16]_o , \xor_i0[16]_i1[16]_o , \xor_i0[17]_i1[17]_o );
  or \or_xor_i0[18]_i1[18]  (\or_xor_i0[18]_i1[18]_o , \xor_i0[18]_i1[18]_o , \or_xor_i0[19]_i1[19]_o );
  or \or_xor_i0[19]_i1[19]  (\or_xor_i0[19]_i1[19]_o , \xor_i0[19]_i1[19]_o , \xor_i0[20]_i1[20]_o );
  or \or_xor_i0[1]_i1[1]_o  (\or_xor_i0[1]_i1[1]_o_o , \xor_i0[1]_i1[1]_o , \xor_i0[2]_i1[2]_o );
  or \or_xor_i0[21]_i1[21]  (\or_xor_i0[21]_i1[21]_o , \xor_i0[21]_i1[21]_o , \or_xor_i0[22]_i1[22]_o );
  or \or_xor_i0[22]_i1[22]  (\or_xor_i0[22]_i1[22]_o , \xor_i0[22]_i1[22]_o , \xor_i0[23]_i1[23]_o );
  or \or_xor_i0[3]_i1[3]_o  (\or_xor_i0[3]_i1[3]_o_o , \xor_i0[3]_i1[3]_o , \or_xor_i0[4]_i1[4]_o_o );
  or \or_xor_i0[4]_i1[4]_o  (\or_xor_i0[4]_i1[4]_o_o , \xor_i0[4]_i1[4]_o , \xor_i0[5]_i1[5]_o );
  or \or_xor_i0[6]_i1[6]_o  (\or_xor_i0[6]_i1[6]_o_o , \xor_i0[6]_i1[6]_o , \or_xor_i0[7]_i1[7]_o_o );
  or \or_xor_i0[7]_i1[7]_o  (\or_xor_i0[7]_i1[7]_o_o , \xor_i0[7]_i1[7]_o , \xor_i0[8]_i1[8]_o );
  or \or_xor_i0[9]_i1[9]_o  (\or_xor_i0[9]_i1[9]_o_o , \xor_i0[9]_i1[9]_o , \or_xor_i0[10]_i1[10]_o );
  xor \xor_i0[0]_i1[0]  (\xor_i0[0]_i1[0]_o , i0[0], i1[0]);
  xor \xor_i0[10]_i1[10]  (\xor_i0[10]_i1[10]_o , i0[10], i1[10]);
  xor \xor_i0[11]_i1[11]  (\xor_i0[11]_i1[11]_o , i0[11], i1[11]);
  xor \xor_i0[12]_i1[12]  (\xor_i0[12]_i1[12]_o , i0[12], i1[12]);
  xor \xor_i0[13]_i1[13]  (\xor_i0[13]_i1[13]_o , i0[13], i1[13]);
  xor \xor_i0[14]_i1[14]  (\xor_i0[14]_i1[14]_o , i0[14], i1[14]);
  xor \xor_i0[15]_i1[15]  (\xor_i0[15]_i1[15]_o , i0[15], i1[15]);
  xor \xor_i0[16]_i1[16]  (\xor_i0[16]_i1[16]_o , i0[16], i1[16]);
  xor \xor_i0[17]_i1[17]  (\xor_i0[17]_i1[17]_o , i0[17], i1[17]);
  xor \xor_i0[18]_i1[18]  (\xor_i0[18]_i1[18]_o , i0[18], i1[18]);
  xor \xor_i0[19]_i1[19]  (\xor_i0[19]_i1[19]_o , i0[19], i1[19]);
  xor \xor_i0[1]_i1[1]  (\xor_i0[1]_i1[1]_o , i0[1], i1[1]);
  xor \xor_i0[20]_i1[20]  (\xor_i0[20]_i1[20]_o , i0[20], i1[20]);
  xor \xor_i0[21]_i1[21]  (\xor_i0[21]_i1[21]_o , i0[21], i1[21]);
  xor \xor_i0[22]_i1[22]  (\xor_i0[22]_i1[22]_o , i0[22], i1[22]);
  xor \xor_i0[23]_i1[23]  (\xor_i0[23]_i1[23]_o , i0[23], i1[23]);
  xor \xor_i0[2]_i1[2]  (\xor_i0[2]_i1[2]_o , i0[2], i1[2]);
  xor \xor_i0[3]_i1[3]  (\xor_i0[3]_i1[3]_o , i0[3], i1[3]);
  xor \xor_i0[4]_i1[4]  (\xor_i0[4]_i1[4]_o , i0[4], i1[4]);
  xor \xor_i0[5]_i1[5]  (\xor_i0[5]_i1[5]_o , i0[5], i1[5]);
  xor \xor_i0[6]_i1[6]  (\xor_i0[6]_i1[6]_o , i0[6], i1[6]);
  xor \xor_i0[7]_i1[7]  (\xor_i0[7]_i1[7]_o , i0[7], i1[7]);
  xor \xor_i0[8]_i1[8]  (\xor_i0[8]_i1[8]_o , i0[8], i1[8]);
  xor \xor_i0[9]_i1[9]  (\xor_i0[9]_i1[9]_o , i0[9], i1[9]);

endmodule 

module binary_mux_s1_w1
  (
  i0,
  i1,
  sel,
  o
  );

  input i0;
  input i1;
  input sel;
  output o;


  AL_MUX al_mux_b0_0_0 (
    .i0(i0),
    .i1(i1),
    .sel(sel),
    .o(o));

endmodule 

module ne_w24
  (
  i0,
  i1,
  o
  );

  input [23:0] i0;
  input [23:0] i1;
  output o;

  wire [23:0] diff;

  or any_diff (o, diff[0], diff[1], diff[2], diff[3], diff[4], diff[5], diff[6], diff[7], diff[8], diff[9], diff[10], diff[11], diff[12], diff[13], diff[14], diff[15], diff[16], diff[17], diff[18], diff[19], diff[20], diff[21], diff[22], diff[23]);
  xor diff_0 (diff[0], i0[0], i1[0]);
  xor diff_1 (diff[1], i0[1], i1[1]);
  xor diff_10 (diff[10], i0[10], i1[10]);
  xor diff_11 (diff[11], i0[11], i1[11]);
  xor diff_12 (diff[12], i0[12], i1[12]);
  xor diff_13 (diff[13], i0[13], i1[13]);
  xor diff_14 (diff[14], i0[14], i1[14]);
  xor diff_15 (diff[15], i0[15], i1[15]);
  xor diff_16 (diff[16], i0[16], i1[16]);
  xor diff_17 (diff[17], i0[17], i1[17]);
  xor diff_18 (diff[18], i0[18], i1[18]);
  xor diff_19 (diff[19], i0[19], i1[19]);
  xor diff_2 (diff[2], i0[2], i1[2]);
  xor diff_20 (diff[20], i0[20], i1[20]);
  xor diff_21 (diff[21], i0[21], i1[21]);
  xor diff_22 (diff[22], i0[22], i1[22]);
  xor diff_23 (diff[23], i0[23], i1[23]);
  xor diff_3 (diff[3], i0[3], i1[3]);
  xor diff_4 (diff[4], i0[4], i1[4]);
  xor diff_5 (diff[5], i0[5], i1[5]);
  xor diff_6 (diff[6], i0[6], i1[6]);
  xor diff_7 (diff[7], i0[7], i1[7]);
  xor diff_8 (diff[8], i0[8], i1[8]);
  xor diff_9 (diff[9], i0[9], i1[9]);

endmodule 

module reg_sr_ss_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  parameter REGSET = "RESET";
  wire enout;
  wire resetout;
  wire setout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_MUX u_reset0 (
    .i0(setout),
    .i1(1'b0),
    .sel(reset),
    .o(resetout));
  AL_DFF #(
    .INI((REGSET == "SET") ? 1'b1 : 1'b0))
    u_seq0 (
    .clk(clk),
    .d(resetout),
    .reset(1'b0),
    .set(1'b0),
    .q(q));
  AL_MUX u_set0 (
    .i0(enout),
    .i1(1'b1),
    .sel(set),
    .o(setout));

endmodule 

module reg_sr_as_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  parameter REGSET = "RESET";
  wire enout;
  wire resetout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_MUX u_reset0 (
    .i0(enout),
    .i1(1'b0),
    .sel(reset),
    .o(resetout));
  AL_DFF #(
    .INI((REGSET == "SET") ? 1'b1 : 1'b0))
    u_seq0 (
    .clk(clk),
    .d(resetout),
    .reset(1'b0),
    .set(set),
    .q(q));

endmodule 

module reg_ar_ss_w1
  (
  clk,
  d,
  en,
  reset,
  set,
  q
  );

  input clk;
  input d;
  input en;
  input reset;
  input set;
  output q;

  parameter REGSET = "RESET";
  wire enout;
  wire setout;

  AL_MUX u_en0 (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_DFF #(
    .INI((REGSET == "SET") ? 1'b1 : 1'b0))
    u_seq0 (
    .clk(clk),
    .d(setout),
    .reset(reset),
    .set(1'b0),
    .q(q));
  AL_MUX u_set0 (
    .i0(enout),
    .i1(1'b1),
    .sel(set),
    .o(setout));

endmodule 

module add_pu27_mu27_o27
  (
  i0,
  i1,
  o
  );

  input [26:0] i0;
  input [26:0] i1;
  output [26:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a10;
  wire net_a11;
  wire net_a12;
  wire net_a13;
  wire net_a14;
  wire net_a15;
  wire net_a16;
  wire net_a17;
  wire net_a18;
  wire net_a19;
  wire net_a2;
  wire net_a20;
  wire net_a21;
  wire net_a22;
  wire net_a23;
  wire net_a24;
  wire net_a25;
  wire net_a26;
  wire net_a3;
  wire net_a4;
  wire net_a5;
  wire net_a6;
  wire net_a7;
  wire net_a8;
  wire net_a9;
  wire net_b0;
  wire net_b1;
  wire net_b10;
  wire net_b11;
  wire net_b12;
  wire net_b13;
  wire net_b14;
  wire net_b15;
  wire net_b16;
  wire net_b17;
  wire net_b18;
  wire net_b19;
  wire net_b2;
  wire net_b20;
  wire net_b21;
  wire net_b22;
  wire net_b23;
  wire net_b24;
  wire net_b25;
  wire net_b26;
  wire net_b3;
  wire net_b4;
  wire net_b5;
  wire net_b6;
  wire net_b7;
  wire net_b8;
  wire net_b9;
  wire net_cout0;
  wire net_cout1;
  wire net_cout10;
  wire net_cout11;
  wire net_cout12;
  wire net_cout13;
  wire net_cout14;
  wire net_cout15;
  wire net_cout16;
  wire net_cout17;
  wire net_cout18;
  wire net_cout19;
  wire net_cout2;
  wire net_cout20;
  wire net_cout21;
  wire net_cout22;
  wire net_cout23;
  wire net_cout24;
  wire net_cout25;
  wire net_cout26;
  wire net_cout3;
  wire net_cout4;
  wire net_cout5;
  wire net_cout6;
  wire net_cout7;
  wire net_cout8;
  wire net_cout9;
  wire net_nb0;
  wire net_nb1;
  wire net_nb10;
  wire net_nb11;
  wire net_nb12;
  wire net_nb13;
  wire net_nb14;
  wire net_nb15;
  wire net_nb16;
  wire net_nb17;
  wire net_nb18;
  wire net_nb19;
  wire net_nb2;
  wire net_nb20;
  wire net_nb21;
  wire net_nb22;
  wire net_nb23;
  wire net_nb24;
  wire net_nb25;
  wire net_nb26;
  wire net_nb3;
  wire net_nb4;
  wire net_nb5;
  wire net_nb6;
  wire net_nb7;
  wire net_nb8;
  wire net_nb9;
  wire net_sum0;
  wire net_sum1;
  wire net_sum10;
  wire net_sum11;
  wire net_sum12;
  wire net_sum13;
  wire net_sum14;
  wire net_sum15;
  wire net_sum16;
  wire net_sum17;
  wire net_sum18;
  wire net_sum19;
  wire net_sum2;
  wire net_sum20;
  wire net_sum21;
  wire net_sum22;
  wire net_sum23;
  wire net_sum24;
  wire net_sum25;
  wire net_sum26;
  wire net_sum3;
  wire net_sum4;
  wire net_sum5;
  wire net_sum6;
  wire net_sum7;
  wire net_sum8;
  wire net_sum9;

  assign net_a26 = i0[26];
  assign net_a25 = i0[25];
  assign net_a24 = i0[24];
  assign net_a23 = i0[23];
  assign net_a22 = i0[22];
  assign net_a21 = i0[21];
  assign net_a20 = i0[20];
  assign net_a19 = i0[19];
  assign net_a18 = i0[18];
  assign net_a17 = i0[17];
  assign net_a16 = i0[16];
  assign net_a15 = i0[15];
  assign net_a14 = i0[14];
  assign net_a13 = i0[13];
  assign net_a12 = i0[12];
  assign net_a11 = i0[11];
  assign net_a10 = i0[10];
  assign net_a9 = i0[9];
  assign net_a8 = i0[8];
  assign net_a7 = i0[7];
  assign net_a6 = i0[6];
  assign net_a5 = i0[5];
  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b26 = i1[26];
  assign net_b25 = i1[25];
  assign net_b24 = i1[24];
  assign net_b23 = i1[23];
  assign net_b22 = i1[22];
  assign net_b21 = i1[21];
  assign net_b20 = i1[20];
  assign net_b19 = i1[19];
  assign net_b18 = i1[18];
  assign net_b17 = i1[17];
  assign net_b16 = i1[16];
  assign net_b15 = i1[15];
  assign net_b14 = i1[14];
  assign net_b13 = i1[13];
  assign net_b12 = i1[12];
  assign net_b11 = i1[11];
  assign net_b10 = i1[10];
  assign net_b9 = i1[9];
  assign net_b8 = i1[8];
  assign net_b7 = i1[7];
  assign net_b6 = i1[6];
  assign net_b5 = i1[5];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[26] = net_sum26;
  assign o[25] = net_sum25;
  assign o[24] = net_sum24;
  assign o[23] = net_sum23;
  assign o[22] = net_sum22;
  assign o[21] = net_sum21;
  assign o[20] = net_sum20;
  assign o[19] = net_sum19;
  assign o[18] = net_sum18;
  assign o[17] = net_sum17;
  assign o[16] = net_sum16;
  assign o[15] = net_sum15;
  assign o[14] = net_sum14;
  assign o[13] = net_sum13;
  assign o[12] = net_sum12;
  assign o[11] = net_sum11;
  assign o[10] = net_sum10;
  assign o[9] = net_sum9;
  assign o[8] = net_sum8;
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_nb0),
    .c(1'b1),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_nb1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_10 (
    .a(net_a10),
    .b(net_nb10),
    .c(net_cout9),
    .cout(net_cout10),
    .sum(net_sum10));
  AL_FADD comp_11 (
    .a(net_a11),
    .b(net_nb11),
    .c(net_cout10),
    .cout(net_cout11),
    .sum(net_sum11));
  AL_FADD comp_12 (
    .a(net_a12),
    .b(net_nb12),
    .c(net_cout11),
    .cout(net_cout12),
    .sum(net_sum12));
  AL_FADD comp_13 (
    .a(net_a13),
    .b(net_nb13),
    .c(net_cout12),
    .cout(net_cout13),
    .sum(net_sum13));
  AL_FADD comp_14 (
    .a(net_a14),
    .b(net_nb14),
    .c(net_cout13),
    .cout(net_cout14),
    .sum(net_sum14));
  AL_FADD comp_15 (
    .a(net_a15),
    .b(net_nb15),
    .c(net_cout14),
    .cout(net_cout15),
    .sum(net_sum15));
  AL_FADD comp_16 (
    .a(net_a16),
    .b(net_nb16),
    .c(net_cout15),
    .cout(net_cout16),
    .sum(net_sum16));
  AL_FADD comp_17 (
    .a(net_a17),
    .b(net_nb17),
    .c(net_cout16),
    .cout(net_cout17),
    .sum(net_sum17));
  AL_FADD comp_18 (
    .a(net_a18),
    .b(net_nb18),
    .c(net_cout17),
    .cout(net_cout18),
    .sum(net_sum18));
  AL_FADD comp_19 (
    .a(net_a19),
    .b(net_nb19),
    .c(net_cout18),
    .cout(net_cout19),
    .sum(net_sum19));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_nb2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_20 (
    .a(net_a20),
    .b(net_nb20),
    .c(net_cout19),
    .cout(net_cout20),
    .sum(net_sum20));
  AL_FADD comp_21 (
    .a(net_a21),
    .b(net_nb21),
    .c(net_cout20),
    .cout(net_cout21),
    .sum(net_sum21));
  AL_FADD comp_22 (
    .a(net_a22),
    .b(net_nb22),
    .c(net_cout21),
    .cout(net_cout22),
    .sum(net_sum22));
  AL_FADD comp_23 (
    .a(net_a23),
    .b(net_nb23),
    .c(net_cout22),
    .cout(net_cout23),
    .sum(net_sum23));
  AL_FADD comp_24 (
    .a(net_a24),
    .b(net_nb24),
    .c(net_cout23),
    .cout(net_cout24),
    .sum(net_sum24));
  AL_FADD comp_25 (
    .a(net_a25),
    .b(net_nb25),
    .c(net_cout24),
    .cout(net_cout25),
    .sum(net_sum25));
  AL_FADD comp_26 (
    .a(net_a26),
    .b(net_nb26),
    .c(net_cout25),
    .cout(net_cout26),
    .sum(net_sum26));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_nb3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_nb4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_5 (
    .a(net_a5),
    .b(net_nb5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_6 (
    .a(net_a6),
    .b(net_nb6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_7 (
    .a(net_a7),
    .b(net_nb7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));
  AL_FADD comp_8 (
    .a(net_a8),
    .b(net_nb8),
    .c(net_cout7),
    .cout(net_cout8),
    .sum(net_sum8));
  AL_FADD comp_9 (
    .a(net_a9),
    .b(net_nb9),
    .c(net_cout8),
    .cout(net_cout9),
    .sum(net_sum9));
  not inv_b0 (net_nb0, net_b0);
  not inv_b1 (net_nb1, net_b1);
  not inv_b10 (net_nb10, net_b10);
  not inv_b11 (net_nb11, net_b11);
  not inv_b12 (net_nb12, net_b12);
  not inv_b13 (net_nb13, net_b13);
  not inv_b14 (net_nb14, net_b14);
  not inv_b15 (net_nb15, net_b15);
  not inv_b16 (net_nb16, net_b16);
  not inv_b17 (net_nb17, net_b17);
  not inv_b18 (net_nb18, net_b18);
  not inv_b19 (net_nb19, net_b19);
  not inv_b2 (net_nb2, net_b2);
  not inv_b20 (net_nb20, net_b20);
  not inv_b21 (net_nb21, net_b21);
  not inv_b22 (net_nb22, net_b22);
  not inv_b23 (net_nb23, net_b23);
  not inv_b24 (net_nb24, net_b24);
  not inv_b25 (net_nb25, net_b25);
  not inv_b26 (net_nb26, net_b26);
  not inv_b3 (net_nb3, net_b3);
  not inv_b4 (net_nb4, net_b4);
  not inv_b5 (net_nb5, net_b5);
  not inv_b6 (net_nb6, net_b6);
  not inv_b7 (net_nb7, net_b7);
  not inv_b8 (net_nb8, net_b8);
  not inv_b9 (net_nb9, net_b9);

endmodule 

module add_pu24_mu24_o24
  (
  i0,
  i1,
  o
  );

  input [23:0] i0;
  input [23:0] i1;
  output [23:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a10;
  wire net_a11;
  wire net_a12;
  wire net_a13;
  wire net_a14;
  wire net_a15;
  wire net_a16;
  wire net_a17;
  wire net_a18;
  wire net_a19;
  wire net_a2;
  wire net_a20;
  wire net_a21;
  wire net_a22;
  wire net_a23;
  wire net_a3;
  wire net_a4;
  wire net_a5;
  wire net_a6;
  wire net_a7;
  wire net_a8;
  wire net_a9;
  wire net_b0;
  wire net_b1;
  wire net_b10;
  wire net_b11;
  wire net_b12;
  wire net_b13;
  wire net_b14;
  wire net_b15;
  wire net_b16;
  wire net_b17;
  wire net_b18;
  wire net_b19;
  wire net_b2;
  wire net_b20;
  wire net_b21;
  wire net_b22;
  wire net_b23;
  wire net_b3;
  wire net_b4;
  wire net_b5;
  wire net_b6;
  wire net_b7;
  wire net_b8;
  wire net_b9;
  wire net_cout0;
  wire net_cout1;
  wire net_cout10;
  wire net_cout11;
  wire net_cout12;
  wire net_cout13;
  wire net_cout14;
  wire net_cout15;
  wire net_cout16;
  wire net_cout17;
  wire net_cout18;
  wire net_cout19;
  wire net_cout2;
  wire net_cout20;
  wire net_cout21;
  wire net_cout22;
  wire net_cout23;
  wire net_cout3;
  wire net_cout4;
  wire net_cout5;
  wire net_cout6;
  wire net_cout7;
  wire net_cout8;
  wire net_cout9;
  wire net_nb0;
  wire net_nb1;
  wire net_nb10;
  wire net_nb11;
  wire net_nb12;
  wire net_nb13;
  wire net_nb14;
  wire net_nb15;
  wire net_nb16;
  wire net_nb17;
  wire net_nb18;
  wire net_nb19;
  wire net_nb2;
  wire net_nb20;
  wire net_nb21;
  wire net_nb22;
  wire net_nb23;
  wire net_nb3;
  wire net_nb4;
  wire net_nb5;
  wire net_nb6;
  wire net_nb7;
  wire net_nb8;
  wire net_nb9;
  wire net_sum0;
  wire net_sum1;
  wire net_sum10;
  wire net_sum11;
  wire net_sum12;
  wire net_sum13;
  wire net_sum14;
  wire net_sum15;
  wire net_sum16;
  wire net_sum17;
  wire net_sum18;
  wire net_sum19;
  wire net_sum2;
  wire net_sum20;
  wire net_sum21;
  wire net_sum22;
  wire net_sum23;
  wire net_sum3;
  wire net_sum4;
  wire net_sum5;
  wire net_sum6;
  wire net_sum7;
  wire net_sum8;
  wire net_sum9;

  assign net_a23 = i0[23];
  assign net_a22 = i0[22];
  assign net_a21 = i0[21];
  assign net_a20 = i0[20];
  assign net_a19 = i0[19];
  assign net_a18 = i0[18];
  assign net_a17 = i0[17];
  assign net_a16 = i0[16];
  assign net_a15 = i0[15];
  assign net_a14 = i0[14];
  assign net_a13 = i0[13];
  assign net_a12 = i0[12];
  assign net_a11 = i0[11];
  assign net_a10 = i0[10];
  assign net_a9 = i0[9];
  assign net_a8 = i0[8];
  assign net_a7 = i0[7];
  assign net_a6 = i0[6];
  assign net_a5 = i0[5];
  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b23 = i1[23];
  assign net_b22 = i1[22];
  assign net_b21 = i1[21];
  assign net_b20 = i1[20];
  assign net_b19 = i1[19];
  assign net_b18 = i1[18];
  assign net_b17 = i1[17];
  assign net_b16 = i1[16];
  assign net_b15 = i1[15];
  assign net_b14 = i1[14];
  assign net_b13 = i1[13];
  assign net_b12 = i1[12];
  assign net_b11 = i1[11];
  assign net_b10 = i1[10];
  assign net_b9 = i1[9];
  assign net_b8 = i1[8];
  assign net_b7 = i1[7];
  assign net_b6 = i1[6];
  assign net_b5 = i1[5];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[23] = net_sum23;
  assign o[22] = net_sum22;
  assign o[21] = net_sum21;
  assign o[20] = net_sum20;
  assign o[19] = net_sum19;
  assign o[18] = net_sum18;
  assign o[17] = net_sum17;
  assign o[16] = net_sum16;
  assign o[15] = net_sum15;
  assign o[14] = net_sum14;
  assign o[13] = net_sum13;
  assign o[12] = net_sum12;
  assign o[11] = net_sum11;
  assign o[10] = net_sum10;
  assign o[9] = net_sum9;
  assign o[8] = net_sum8;
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_nb0),
    .c(1'b1),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_nb1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_10 (
    .a(net_a10),
    .b(net_nb10),
    .c(net_cout9),
    .cout(net_cout10),
    .sum(net_sum10));
  AL_FADD comp_11 (
    .a(net_a11),
    .b(net_nb11),
    .c(net_cout10),
    .cout(net_cout11),
    .sum(net_sum11));
  AL_FADD comp_12 (
    .a(net_a12),
    .b(net_nb12),
    .c(net_cout11),
    .cout(net_cout12),
    .sum(net_sum12));
  AL_FADD comp_13 (
    .a(net_a13),
    .b(net_nb13),
    .c(net_cout12),
    .cout(net_cout13),
    .sum(net_sum13));
  AL_FADD comp_14 (
    .a(net_a14),
    .b(net_nb14),
    .c(net_cout13),
    .cout(net_cout14),
    .sum(net_sum14));
  AL_FADD comp_15 (
    .a(net_a15),
    .b(net_nb15),
    .c(net_cout14),
    .cout(net_cout15),
    .sum(net_sum15));
  AL_FADD comp_16 (
    .a(net_a16),
    .b(net_nb16),
    .c(net_cout15),
    .cout(net_cout16),
    .sum(net_sum16));
  AL_FADD comp_17 (
    .a(net_a17),
    .b(net_nb17),
    .c(net_cout16),
    .cout(net_cout17),
    .sum(net_sum17));
  AL_FADD comp_18 (
    .a(net_a18),
    .b(net_nb18),
    .c(net_cout17),
    .cout(net_cout18),
    .sum(net_sum18));
  AL_FADD comp_19 (
    .a(net_a19),
    .b(net_nb19),
    .c(net_cout18),
    .cout(net_cout19),
    .sum(net_sum19));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_nb2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_20 (
    .a(net_a20),
    .b(net_nb20),
    .c(net_cout19),
    .cout(net_cout20),
    .sum(net_sum20));
  AL_FADD comp_21 (
    .a(net_a21),
    .b(net_nb21),
    .c(net_cout20),
    .cout(net_cout21),
    .sum(net_sum21));
  AL_FADD comp_22 (
    .a(net_a22),
    .b(net_nb22),
    .c(net_cout21),
    .cout(net_cout22),
    .sum(net_sum22));
  AL_FADD comp_23 (
    .a(net_a23),
    .b(net_nb23),
    .c(net_cout22),
    .cout(net_cout23),
    .sum(net_sum23));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_nb3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_nb4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_5 (
    .a(net_a5),
    .b(net_nb5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_6 (
    .a(net_a6),
    .b(net_nb6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_7 (
    .a(net_a7),
    .b(net_nb7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));
  AL_FADD comp_8 (
    .a(net_a8),
    .b(net_nb8),
    .c(net_cout7),
    .cout(net_cout8),
    .sum(net_sum8));
  AL_FADD comp_9 (
    .a(net_a9),
    .b(net_nb9),
    .c(net_cout8),
    .cout(net_cout9),
    .sum(net_sum9));
  not inv_b0 (net_nb0, net_b0);
  not inv_b1 (net_nb1, net_b1);
  not inv_b10 (net_nb10, net_b10);
  not inv_b11 (net_nb11, net_b11);
  not inv_b12 (net_nb12, net_b12);
  not inv_b13 (net_nb13, net_b13);
  not inv_b14 (net_nb14, net_b14);
  not inv_b15 (net_nb15, net_b15);
  not inv_b16 (net_nb16, net_b16);
  not inv_b17 (net_nb17, net_b17);
  not inv_b18 (net_nb18, net_b18);
  not inv_b19 (net_nb19, net_b19);
  not inv_b2 (net_nb2, net_b2);
  not inv_b20 (net_nb20, net_b20);
  not inv_b21 (net_nb21, net_b21);
  not inv_b22 (net_nb22, net_b22);
  not inv_b23 (net_nb23, net_b23);
  not inv_b3 (net_nb3, net_b3);
  not inv_b4 (net_nb4, net_b4);
  not inv_b5 (net_nb5, net_b5);
  not inv_b6 (net_nb6, net_b6);
  not inv_b7 (net_nb7, net_b7);
  not inv_b8 (net_nb8, net_b8);
  not inv_b9 (net_nb9, net_b9);

endmodule 

module eq_w2
  (
  i0,
  i1,
  o
  );

  input [1:0] i0;
  input [1:0] i1;
  output o;

  wire \or_xor_i0[0]_i1[0]_o_o ;
  wire \xor_i0[0]_i1[0]_o ;
  wire \xor_i0[1]_i1[1]_o ;

  not none_diff (o, \or_xor_i0[0]_i1[0]_o_o );
  or \or_xor_i0[0]_i1[0]_o  (\or_xor_i0[0]_i1[0]_o_o , \xor_i0[0]_i1[0]_o , \xor_i0[1]_i1[1]_o );
  xor \xor_i0[0]_i1[0]  (\xor_i0[0]_i1[0]_o , i0[0], i1[0]);
  xor \xor_i0[1]_i1[1]  (\xor_i0[1]_i1[1]_o , i0[1], i1[1]);

endmodule 

module add_pu32_pu32_o32
  (
  i0,
  i1,
  o
  );

  input [31:0] i0;
  input [31:0] i1;
  output [31:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a10;
  wire net_a11;
  wire net_a12;
  wire net_a13;
  wire net_a14;
  wire net_a15;
  wire net_a16;
  wire net_a17;
  wire net_a18;
  wire net_a19;
  wire net_a2;
  wire net_a20;
  wire net_a21;
  wire net_a22;
  wire net_a23;
  wire net_a24;
  wire net_a25;
  wire net_a26;
  wire net_a27;
  wire net_a28;
  wire net_a29;
  wire net_a3;
  wire net_a30;
  wire net_a31;
  wire net_a4;
  wire net_a5;
  wire net_a6;
  wire net_a7;
  wire net_a8;
  wire net_a9;
  wire net_b0;
  wire net_b1;
  wire net_b10;
  wire net_b11;
  wire net_b12;
  wire net_b13;
  wire net_b14;
  wire net_b15;
  wire net_b16;
  wire net_b17;
  wire net_b18;
  wire net_b19;
  wire net_b2;
  wire net_b20;
  wire net_b21;
  wire net_b22;
  wire net_b23;
  wire net_b24;
  wire net_b25;
  wire net_b26;
  wire net_b27;
  wire net_b28;
  wire net_b29;
  wire net_b3;
  wire net_b30;
  wire net_b31;
  wire net_b4;
  wire net_b5;
  wire net_b6;
  wire net_b7;
  wire net_b8;
  wire net_b9;
  wire net_cout0;
  wire net_cout1;
  wire net_cout10;
  wire net_cout11;
  wire net_cout12;
  wire net_cout13;
  wire net_cout14;
  wire net_cout15;
  wire net_cout16;
  wire net_cout17;
  wire net_cout18;
  wire net_cout19;
  wire net_cout2;
  wire net_cout20;
  wire net_cout21;
  wire net_cout22;
  wire net_cout23;
  wire net_cout24;
  wire net_cout25;
  wire net_cout26;
  wire net_cout27;
  wire net_cout28;
  wire net_cout29;
  wire net_cout3;
  wire net_cout30;
  wire net_cout31;
  wire net_cout4;
  wire net_cout5;
  wire net_cout6;
  wire net_cout7;
  wire net_cout8;
  wire net_cout9;
  wire net_sum0;
  wire net_sum1;
  wire net_sum10;
  wire net_sum11;
  wire net_sum12;
  wire net_sum13;
  wire net_sum14;
  wire net_sum15;
  wire net_sum16;
  wire net_sum17;
  wire net_sum18;
  wire net_sum19;
  wire net_sum2;
  wire net_sum20;
  wire net_sum21;
  wire net_sum22;
  wire net_sum23;
  wire net_sum24;
  wire net_sum25;
  wire net_sum26;
  wire net_sum27;
  wire net_sum28;
  wire net_sum29;
  wire net_sum3;
  wire net_sum30;
  wire net_sum31;
  wire net_sum4;
  wire net_sum5;
  wire net_sum6;
  wire net_sum7;
  wire net_sum8;
  wire net_sum9;

  assign net_a31 = i0[31];
  assign net_a30 = i0[30];
  assign net_a29 = i0[29];
  assign net_a28 = i0[28];
  assign net_a27 = i0[27];
  assign net_a26 = i0[26];
  assign net_a25 = i0[25];
  assign net_a24 = i0[24];
  assign net_a23 = i0[23];
  assign net_a22 = i0[22];
  assign net_a21 = i0[21];
  assign net_a20 = i0[20];
  assign net_a19 = i0[19];
  assign net_a18 = i0[18];
  assign net_a17 = i0[17];
  assign net_a16 = i0[16];
  assign net_a15 = i0[15];
  assign net_a14 = i0[14];
  assign net_a13 = i0[13];
  assign net_a12 = i0[12];
  assign net_a11 = i0[11];
  assign net_a10 = i0[10];
  assign net_a9 = i0[9];
  assign net_a8 = i0[8];
  assign net_a7 = i0[7];
  assign net_a6 = i0[6];
  assign net_a5 = i0[5];
  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b31 = i1[31];
  assign net_b30 = i1[30];
  assign net_b29 = i1[29];
  assign net_b28 = i1[28];
  assign net_b27 = i1[27];
  assign net_b26 = i1[26];
  assign net_b25 = i1[25];
  assign net_b24 = i1[24];
  assign net_b23 = i1[23];
  assign net_b22 = i1[22];
  assign net_b21 = i1[21];
  assign net_b20 = i1[20];
  assign net_b19 = i1[19];
  assign net_b18 = i1[18];
  assign net_b17 = i1[17];
  assign net_b16 = i1[16];
  assign net_b15 = i1[15];
  assign net_b14 = i1[14];
  assign net_b13 = i1[13];
  assign net_b12 = i1[12];
  assign net_b11 = i1[11];
  assign net_b10 = i1[10];
  assign net_b9 = i1[9];
  assign net_b8 = i1[8];
  assign net_b7 = i1[7];
  assign net_b6 = i1[6];
  assign net_b5 = i1[5];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[31] = net_sum31;
  assign o[30] = net_sum30;
  assign o[29] = net_sum29;
  assign o[28] = net_sum28;
  assign o[27] = net_sum27;
  assign o[26] = net_sum26;
  assign o[25] = net_sum25;
  assign o[24] = net_sum24;
  assign o[23] = net_sum23;
  assign o[22] = net_sum22;
  assign o[21] = net_sum21;
  assign o[20] = net_sum20;
  assign o[19] = net_sum19;
  assign o[18] = net_sum18;
  assign o[17] = net_sum17;
  assign o[16] = net_sum16;
  assign o[15] = net_sum15;
  assign o[14] = net_sum14;
  assign o[13] = net_sum13;
  assign o[12] = net_sum12;
  assign o[11] = net_sum11;
  assign o[10] = net_sum10;
  assign o[9] = net_sum9;
  assign o[8] = net_sum8;
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_b0),
    .c(1'b0),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_b1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_10 (
    .a(net_a10),
    .b(net_b10),
    .c(net_cout9),
    .cout(net_cout10),
    .sum(net_sum10));
  AL_FADD comp_11 (
    .a(net_a11),
    .b(net_b11),
    .c(net_cout10),
    .cout(net_cout11),
    .sum(net_sum11));
  AL_FADD comp_12 (
    .a(net_a12),
    .b(net_b12),
    .c(net_cout11),
    .cout(net_cout12),
    .sum(net_sum12));
  AL_FADD comp_13 (
    .a(net_a13),
    .b(net_b13),
    .c(net_cout12),
    .cout(net_cout13),
    .sum(net_sum13));
  AL_FADD comp_14 (
    .a(net_a14),
    .b(net_b14),
    .c(net_cout13),
    .cout(net_cout14),
    .sum(net_sum14));
  AL_FADD comp_15 (
    .a(net_a15),
    .b(net_b15),
    .c(net_cout14),
    .cout(net_cout15),
    .sum(net_sum15));
  AL_FADD comp_16 (
    .a(net_a16),
    .b(net_b16),
    .c(net_cout15),
    .cout(net_cout16),
    .sum(net_sum16));
  AL_FADD comp_17 (
    .a(net_a17),
    .b(net_b17),
    .c(net_cout16),
    .cout(net_cout17),
    .sum(net_sum17));
  AL_FADD comp_18 (
    .a(net_a18),
    .b(net_b18),
    .c(net_cout17),
    .cout(net_cout18),
    .sum(net_sum18));
  AL_FADD comp_19 (
    .a(net_a19),
    .b(net_b19),
    .c(net_cout18),
    .cout(net_cout19),
    .sum(net_sum19));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_b2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_20 (
    .a(net_a20),
    .b(net_b20),
    .c(net_cout19),
    .cout(net_cout20),
    .sum(net_sum20));
  AL_FADD comp_21 (
    .a(net_a21),
    .b(net_b21),
    .c(net_cout20),
    .cout(net_cout21),
    .sum(net_sum21));
  AL_FADD comp_22 (
    .a(net_a22),
    .b(net_b22),
    .c(net_cout21),
    .cout(net_cout22),
    .sum(net_sum22));
  AL_FADD comp_23 (
    .a(net_a23),
    .b(net_b23),
    .c(net_cout22),
    .cout(net_cout23),
    .sum(net_sum23));
  AL_FADD comp_24 (
    .a(net_a24),
    .b(net_b24),
    .c(net_cout23),
    .cout(net_cout24),
    .sum(net_sum24));
  AL_FADD comp_25 (
    .a(net_a25),
    .b(net_b25),
    .c(net_cout24),
    .cout(net_cout25),
    .sum(net_sum25));
  AL_FADD comp_26 (
    .a(net_a26),
    .b(net_b26),
    .c(net_cout25),
    .cout(net_cout26),
    .sum(net_sum26));
  AL_FADD comp_27 (
    .a(net_a27),
    .b(net_b27),
    .c(net_cout26),
    .cout(net_cout27),
    .sum(net_sum27));
  AL_FADD comp_28 (
    .a(net_a28),
    .b(net_b28),
    .c(net_cout27),
    .cout(net_cout28),
    .sum(net_sum28));
  AL_FADD comp_29 (
    .a(net_a29),
    .b(net_b29),
    .c(net_cout28),
    .cout(net_cout29),
    .sum(net_sum29));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_b3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_30 (
    .a(net_a30),
    .b(net_b30),
    .c(net_cout29),
    .cout(net_cout30),
    .sum(net_sum30));
  AL_FADD comp_31 (
    .a(net_a31),
    .b(net_b31),
    .c(net_cout30),
    .cout(net_cout31),
    .sum(net_sum31));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_b4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_5 (
    .a(net_a5),
    .b(net_b5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_6 (
    .a(net_a6),
    .b(net_b6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_7 (
    .a(net_a7),
    .b(net_b7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));
  AL_FADD comp_8 (
    .a(net_a8),
    .b(net_b8),
    .c(net_cout7),
    .cout(net_cout8),
    .sum(net_sum8));
  AL_FADD comp_9 (
    .a(net_a9),
    .b(net_b9),
    .c(net_cout8),
    .cout(net_cout9),
    .sum(net_sum9));

endmodule 

module eq_w32
  (
  i0,
  i1,
  o
  );

  input [31:0] i0;
  input [31:0] i1;
  output o;

  wire or_or_or_or_or_xor_i_o;
  wire \or_or_or_or_xor_i0[0_o ;
  wire \or_or_or_or_xor_i0[1_o ;
  wire \or_or_or_xor_i0[0]_i_o ;
  wire \or_or_or_xor_i0[16]__o ;
  wire \or_or_or_xor_i0[24]__o ;
  wire \or_or_or_xor_i0[8]_i_o ;
  wire \or_or_xor_i0[0]_i1[0_o ;
  wire \or_or_xor_i0[12]_i1[_o ;
  wire \or_or_xor_i0[16]_i1[_o ;
  wire \or_or_xor_i0[20]_i1[_o ;
  wire \or_or_xor_i0[24]_i1[_o ;
  wire \or_or_xor_i0[28]_i1[_o ;
  wire \or_or_xor_i0[4]_i1[4_o ;
  wire \or_or_xor_i0[8]_i1[8_o ;
  wire \or_xor_i0[0]_i1[0]_o_o ;
  wire \or_xor_i0[10]_i1[10]_o ;
  wire \or_xor_i0[12]_i1[12]_o ;
  wire \or_xor_i0[14]_i1[14]_o ;
  wire \or_xor_i0[16]_i1[16]_o ;
  wire \or_xor_i0[18]_i1[18]_o ;
  wire \or_xor_i0[20]_i1[20]_o ;
  wire \or_xor_i0[22]_i1[22]_o ;
  wire \or_xor_i0[24]_i1[24]_o ;
  wire \or_xor_i0[26]_i1[26]_o ;
  wire \or_xor_i0[28]_i1[28]_o ;
  wire \or_xor_i0[2]_i1[2]_o_o ;
  wire \or_xor_i0[30]_i1[30]_o ;
  wire \or_xor_i0[4]_i1[4]_o_o ;
  wire \or_xor_i0[6]_i1[6]_o_o ;
  wire \or_xor_i0[8]_i1[8]_o_o ;
  wire \xor_i0[0]_i1[0]_o ;
  wire \xor_i0[10]_i1[10]_o ;
  wire \xor_i0[11]_i1[11]_o ;
  wire \xor_i0[12]_i1[12]_o ;
  wire \xor_i0[13]_i1[13]_o ;
  wire \xor_i0[14]_i1[14]_o ;
  wire \xor_i0[15]_i1[15]_o ;
  wire \xor_i0[16]_i1[16]_o ;
  wire \xor_i0[17]_i1[17]_o ;
  wire \xor_i0[18]_i1[18]_o ;
  wire \xor_i0[19]_i1[19]_o ;
  wire \xor_i0[1]_i1[1]_o ;
  wire \xor_i0[20]_i1[20]_o ;
  wire \xor_i0[21]_i1[21]_o ;
  wire \xor_i0[22]_i1[22]_o ;
  wire \xor_i0[23]_i1[23]_o ;
  wire \xor_i0[24]_i1[24]_o ;
  wire \xor_i0[25]_i1[25]_o ;
  wire \xor_i0[26]_i1[26]_o ;
  wire \xor_i0[27]_i1[27]_o ;
  wire \xor_i0[28]_i1[28]_o ;
  wire \xor_i0[29]_i1[29]_o ;
  wire \xor_i0[2]_i1[2]_o ;
  wire \xor_i0[30]_i1[30]_o ;
  wire \xor_i0[31]_i1[31]_o ;
  wire \xor_i0[3]_i1[3]_o ;
  wire \xor_i0[4]_i1[4]_o ;
  wire \xor_i0[5]_i1[5]_o ;
  wire \xor_i0[6]_i1[6]_o ;
  wire \xor_i0[7]_i1[7]_o ;
  wire \xor_i0[8]_i1[8]_o ;
  wire \xor_i0[9]_i1[9]_o ;

  not none_diff (o, or_or_or_or_or_xor_i_o);
  or or_or_or_or_or_xor_i (or_or_or_or_or_xor_i_o, \or_or_or_or_xor_i0[0_o , \or_or_or_or_xor_i0[1_o );
  or \or_or_or_or_xor_i0[0  (\or_or_or_or_xor_i0[0_o , \or_or_or_xor_i0[0]_i_o , \or_or_or_xor_i0[8]_i_o );
  or \or_or_or_or_xor_i0[1  (\or_or_or_or_xor_i0[1_o , \or_or_or_xor_i0[16]__o , \or_or_or_xor_i0[24]__o );
  or \or_or_or_xor_i0[0]_i  (\or_or_or_xor_i0[0]_i_o , \or_or_xor_i0[0]_i1[0_o , \or_or_xor_i0[4]_i1[4_o );
  or \or_or_or_xor_i0[16]_  (\or_or_or_xor_i0[16]__o , \or_or_xor_i0[16]_i1[_o , \or_or_xor_i0[20]_i1[_o );
  or \or_or_or_xor_i0[24]_  (\or_or_or_xor_i0[24]__o , \or_or_xor_i0[24]_i1[_o , \or_or_xor_i0[28]_i1[_o );
  or \or_or_or_xor_i0[8]_i  (\or_or_or_xor_i0[8]_i_o , \or_or_xor_i0[8]_i1[8_o , \or_or_xor_i0[12]_i1[_o );
  or \or_or_xor_i0[0]_i1[0  (\or_or_xor_i0[0]_i1[0_o , \or_xor_i0[0]_i1[0]_o_o , \or_xor_i0[2]_i1[2]_o_o );
  or \or_or_xor_i0[12]_i1[  (\or_or_xor_i0[12]_i1[_o , \or_xor_i0[12]_i1[12]_o , \or_xor_i0[14]_i1[14]_o );
  or \or_or_xor_i0[16]_i1[  (\or_or_xor_i0[16]_i1[_o , \or_xor_i0[16]_i1[16]_o , \or_xor_i0[18]_i1[18]_o );
  or \or_or_xor_i0[20]_i1[  (\or_or_xor_i0[20]_i1[_o , \or_xor_i0[20]_i1[20]_o , \or_xor_i0[22]_i1[22]_o );
  or \or_or_xor_i0[24]_i1[  (\or_or_xor_i0[24]_i1[_o , \or_xor_i0[24]_i1[24]_o , \or_xor_i0[26]_i1[26]_o );
  or \or_or_xor_i0[28]_i1[  (\or_or_xor_i0[28]_i1[_o , \or_xor_i0[28]_i1[28]_o , \or_xor_i0[30]_i1[30]_o );
  or \or_or_xor_i0[4]_i1[4  (\or_or_xor_i0[4]_i1[4_o , \or_xor_i0[4]_i1[4]_o_o , \or_xor_i0[6]_i1[6]_o_o );
  or \or_or_xor_i0[8]_i1[8  (\or_or_xor_i0[8]_i1[8_o , \or_xor_i0[8]_i1[8]_o_o , \or_xor_i0[10]_i1[10]_o );
  or \or_xor_i0[0]_i1[0]_o  (\or_xor_i0[0]_i1[0]_o_o , \xor_i0[0]_i1[0]_o , \xor_i0[1]_i1[1]_o );
  or \or_xor_i0[10]_i1[10]  (\or_xor_i0[10]_i1[10]_o , \xor_i0[10]_i1[10]_o , \xor_i0[11]_i1[11]_o );
  or \or_xor_i0[12]_i1[12]  (\or_xor_i0[12]_i1[12]_o , \xor_i0[12]_i1[12]_o , \xor_i0[13]_i1[13]_o );
  or \or_xor_i0[14]_i1[14]  (\or_xor_i0[14]_i1[14]_o , \xor_i0[14]_i1[14]_o , \xor_i0[15]_i1[15]_o );
  or \or_xor_i0[16]_i1[16]  (\or_xor_i0[16]_i1[16]_o , \xor_i0[16]_i1[16]_o , \xor_i0[17]_i1[17]_o );
  or \or_xor_i0[18]_i1[18]  (\or_xor_i0[18]_i1[18]_o , \xor_i0[18]_i1[18]_o , \xor_i0[19]_i1[19]_o );
  or \or_xor_i0[20]_i1[20]  (\or_xor_i0[20]_i1[20]_o , \xor_i0[20]_i1[20]_o , \xor_i0[21]_i1[21]_o );
  or \or_xor_i0[22]_i1[22]  (\or_xor_i0[22]_i1[22]_o , \xor_i0[22]_i1[22]_o , \xor_i0[23]_i1[23]_o );
  or \or_xor_i0[24]_i1[24]  (\or_xor_i0[24]_i1[24]_o , \xor_i0[24]_i1[24]_o , \xor_i0[25]_i1[25]_o );
  or \or_xor_i0[26]_i1[26]  (\or_xor_i0[26]_i1[26]_o , \xor_i0[26]_i1[26]_o , \xor_i0[27]_i1[27]_o );
  or \or_xor_i0[28]_i1[28]  (\or_xor_i0[28]_i1[28]_o , \xor_i0[28]_i1[28]_o , \xor_i0[29]_i1[29]_o );
  or \or_xor_i0[2]_i1[2]_o  (\or_xor_i0[2]_i1[2]_o_o , \xor_i0[2]_i1[2]_o , \xor_i0[3]_i1[3]_o );
  or \or_xor_i0[30]_i1[30]  (\or_xor_i0[30]_i1[30]_o , \xor_i0[30]_i1[30]_o , \xor_i0[31]_i1[31]_o );
  or \or_xor_i0[4]_i1[4]_o  (\or_xor_i0[4]_i1[4]_o_o , \xor_i0[4]_i1[4]_o , \xor_i0[5]_i1[5]_o );
  or \or_xor_i0[6]_i1[6]_o  (\or_xor_i0[6]_i1[6]_o_o , \xor_i0[6]_i1[6]_o , \xor_i0[7]_i1[7]_o );
  or \or_xor_i0[8]_i1[8]_o  (\or_xor_i0[8]_i1[8]_o_o , \xor_i0[8]_i1[8]_o , \xor_i0[9]_i1[9]_o );
  xor \xor_i0[0]_i1[0]  (\xor_i0[0]_i1[0]_o , i0[0], i1[0]);
  xor \xor_i0[10]_i1[10]  (\xor_i0[10]_i1[10]_o , i0[10], i1[10]);
  xor \xor_i0[11]_i1[11]  (\xor_i0[11]_i1[11]_o , i0[11], i1[11]);
  xor \xor_i0[12]_i1[12]  (\xor_i0[12]_i1[12]_o , i0[12], i1[12]);
  xor \xor_i0[13]_i1[13]  (\xor_i0[13]_i1[13]_o , i0[13], i1[13]);
  xor \xor_i0[14]_i1[14]  (\xor_i0[14]_i1[14]_o , i0[14], i1[14]);
  xor \xor_i0[15]_i1[15]  (\xor_i0[15]_i1[15]_o , i0[15], i1[15]);
  xor \xor_i0[16]_i1[16]  (\xor_i0[16]_i1[16]_o , i0[16], i1[16]);
  xor \xor_i0[17]_i1[17]  (\xor_i0[17]_i1[17]_o , i0[17], i1[17]);
  xor \xor_i0[18]_i1[18]  (\xor_i0[18]_i1[18]_o , i0[18], i1[18]);
  xor \xor_i0[19]_i1[19]  (\xor_i0[19]_i1[19]_o , i0[19], i1[19]);
  xor \xor_i0[1]_i1[1]  (\xor_i0[1]_i1[1]_o , i0[1], i1[1]);
  xor \xor_i0[20]_i1[20]  (\xor_i0[20]_i1[20]_o , i0[20], i1[20]);
  xor \xor_i0[21]_i1[21]  (\xor_i0[21]_i1[21]_o , i0[21], i1[21]);
  xor \xor_i0[22]_i1[22]  (\xor_i0[22]_i1[22]_o , i0[22], i1[22]);
  xor \xor_i0[23]_i1[23]  (\xor_i0[23]_i1[23]_o , i0[23], i1[23]);
  xor \xor_i0[24]_i1[24]  (\xor_i0[24]_i1[24]_o , i0[24], i1[24]);
  xor \xor_i0[25]_i1[25]  (\xor_i0[25]_i1[25]_o , i0[25], i1[25]);
  xor \xor_i0[26]_i1[26]  (\xor_i0[26]_i1[26]_o , i0[26], i1[26]);
  xor \xor_i0[27]_i1[27]  (\xor_i0[27]_i1[27]_o , i0[27], i1[27]);
  xor \xor_i0[28]_i1[28]  (\xor_i0[28]_i1[28]_o , i0[28], i1[28]);
  xor \xor_i0[29]_i1[29]  (\xor_i0[29]_i1[29]_o , i0[29], i1[29]);
  xor \xor_i0[2]_i1[2]  (\xor_i0[2]_i1[2]_o , i0[2], i1[2]);
  xor \xor_i0[30]_i1[30]  (\xor_i0[30]_i1[30]_o , i0[30], i1[30]);
  xor \xor_i0[31]_i1[31]  (\xor_i0[31]_i1[31]_o , i0[31], i1[31]);
  xor \xor_i0[3]_i1[3]  (\xor_i0[3]_i1[3]_o , i0[3], i1[3]);
  xor \xor_i0[4]_i1[4]  (\xor_i0[4]_i1[4]_o , i0[4], i1[4]);
  xor \xor_i0[5]_i1[5]  (\xor_i0[5]_i1[5]_o , i0[5], i1[5]);
  xor \xor_i0[6]_i1[6]  (\xor_i0[6]_i1[6]_o , i0[6], i1[6]);
  xor \xor_i0[7]_i1[7]  (\xor_i0[7]_i1[7]_o , i0[7], i1[7]);
  xor \xor_i0[8]_i1[8]  (\xor_i0[8]_i1[8]_o , i0[8], i1[8]);
  xor \xor_i0[9]_i1[9]  (\xor_i0[9]_i1[9]_o , i0[9], i1[9]);

endmodule 

module AL_MUX
  (
  input i0,
  input i1,
  input sel,
  output o
  );

  wire not_sel, sel_i0, sel_i1;
  not u0 (not_sel, sel);
  and u1 (sel_i1, sel, i1);
  and u2 (sel_i0, not_sel, i0);
  or u3 (o, sel_i1, sel_i0);

endmodule

module AL_DFF
  (
  input reset,
  input set,
  input clk,
  input d,
  output reg q
  );

  parameter INI = 1'b0;

  always @(posedge reset or posedge set or posedge clk)
  begin
    if (reset)
      q <= 1'b0;
    else if (set)
      q <= 1'b1;
    else
      q <= d;
  end

endmodule

module AL_FADD
  (
  input a,
  input b,
  input c,
  output sum,
  output cout
  );

  wire prop;
  wire not_prop;
  wire sel_i0;
  wire sel_i1;

  xor u0 (prop, a, b);
  xor u1 (sum, prop, c);
  not u2 (not_prop, prop);
  and u3 (sel_i1, prop, c);
  and u4 (sel_i0, not_prop, a);
  or  u5 (cout, sel_i0, sel_i1);

endmodule

